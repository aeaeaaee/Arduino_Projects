PK
     B"BY.u��� �    cirkitFile.json{"raven_core_version":15,"hardware_version":0,"pin_to_graph":{"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg"],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg":["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2"],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1":["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg"],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos":["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2"],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg"],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg"],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos":["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg":["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2"],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29_polarity-pos":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29_polarity-neg":[],"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29":[],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4"],"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_0":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_1":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_2":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_3":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_6":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_7":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_8":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_9":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_10":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_11":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_12":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_13":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14":["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15":["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_16":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_17":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_19":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_22":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_23":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_24":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_25":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5"],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_27":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_28":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_29":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_30":[],"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_31":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos"],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_1":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg"],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14"],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15"],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_5":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_6":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_7":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_8":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_9":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_10":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_11":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_12":[],"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_13":[],"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos"],"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5"],"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg"],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3"],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg"],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg"],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3":["pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7"],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15"],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16":["pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos":["pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos":["pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg":["pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1"],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28":["pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0"],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28_polarity-neg":[],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg":["pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1"],"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29_polarity-pos":[],"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29_polarity-neg":[],"pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28"],"pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg"],"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28"],"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg"],"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos"],"pin-type-component_5102790f-a871-47d9-83fd-2bf45f8f7bb8_0":[],"pin-type-component_5102790f-a871-47d9-83fd-2bf45f8f7bb8_1":[],"pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16"],"pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos"],"pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_0":[],"pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_1":[],"pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_2":[],"pin-type-component_27363330-fd4d-4d48-8fe5-7e75a0bb5506_0":[],"pin-type-component_27363330-fd4d-4d48-8fe5-7e75a0bb5506_1":[],"pin-type-component_9cd4866e-171b-4689-8c74-d7df80f41d58_0":[],"pin-type-component_9cd4866e-171b-4689-8c74-d7df80f41d58_1":[],"pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_0":[],"pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_1":[],"pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_2":[],"pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_0":[],"pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_1":[],"pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_2":[],"pin-type-component_ad1269e6-5014-4c59-af62-685c40e02898_0":[],"pin-type-component_ad1269e6-5014-4c59-af62-685c40e02898_1":[],"pin-type-component_f533a25e-c11a-427c-a4aa-e80fef74288c_0":[],"pin-type-component_f533a25e-c11a-427c-a4aa-e80fef74288c_1":[],"pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8"],"pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3"],"pin-type-component_6e804c70-7bd6-41c1-bf62-acd23076114e_0":[],"pin-type-component_6e804c70-7bd6-41c1-bf62-acd23076114e_1":[],"pin-type-component_dd2abdd4-ed36-4c43-9689-d56c6cb3bd68_0":[],"pin-type-component_dd2abdd4-ed36-4c43-9689-d56c6cb3bd68_1":[],"pin-type-component_66bf0903-9a55-463b-bc47-49eeb06f5fc3_0":[],"pin-type-component_66bf0903-9a55-463b-bc47-49eeb06f5fc3_1":[],"pin-type-component_3845c3bd-f40d-4978-9482-daa8afda013f_0":[],"pin-type-component_3845c3bd-f40d-4978-9482-daa8afda013f_1":[],"pin-type-component_d0b06877-9f19-4217-938d-d5d876016b19_0":[],"pin-type-component_d0b06877-9f19-4217-938d-d5d876016b19_1":[],"pin-type-component_0db723b4-8ee7-4aa5-8efd-d1c37793e604_0":[],"pin-type-component_0db723b4-8ee7-4aa5-8efd-d1c37793e604_1":[],"pin-type-component_d2a8b258-269a-4d63-87df-4ce160f1790a_0":[],"pin-type-component_d2a8b258-269a-4d63-87df-4ce160f1790a_1":[],"pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1"],"pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6"],"pin-type-component_f4f47a18-edf3-46de-9608-c6b22e0dc54e_0":[],"pin-type-component_f4f47a18-edf3-46de-9608-c6b22e0dc54e_1":[]},"pin_to_color":{"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg":"#189AB4","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg":"#189AB4","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1":"#683D3B","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg":"#189AB4","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos":"#FF0000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2":"#189AB4","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg":"#189AB4","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg":"#189AB4","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg":"#189AB4","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5":"#e2e600","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6":"#e70404","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8":"#e70404","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9":"#FF0000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17":"#1ddd03","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos":"#FF0000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg":"#189AB4","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29_polarity-pos":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29_polarity-neg":"#000000","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29":"#000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos":"#FF0000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg":"#189AB4","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_0":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_1":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_2":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_3":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4":"#FF0000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5":"#189AB4","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_6":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_7":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_8":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_9":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_10":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_11":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_12":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_13":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14":"#0E4CA1","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15":"#FFE502","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_16":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_17":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18":"#5ecd13","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_19":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20":"#14db25","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21":"#1ddd03","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_22":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_23":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_24":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_25":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26":"#e2e600","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_27":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_28":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_29":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_30":"#000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_31":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0":"#FF0000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_1":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2":"#189AB4","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3":"#0E4CA1","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4":"#FFE502","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_5":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_6":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_7":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_8":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_9":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_10":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_11":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_12":"#000000","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_13":"#000000","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0":"#FF0000","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1":"#e2e600","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2":"#189AB4","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg":"#189AB4","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg":"#189AB4","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg":"#189AB4","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3":"#189AB4","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg":"#189AB4","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7":"#189AB4","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8":"#e75a0d","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos":"#FF0000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10":"#e75a0d","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11":"#e75a0d","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos":"#FF0000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12":"#FF0000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg":"#189AB4","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15":"#189AB4","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16":"#083a36","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos":"#FF0000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19":"#14db25","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos":"#FF0000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23":"#5ecd13","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg":"#189AB4","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28":"#f20202","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28_polarity-neg":"#000000","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg":"#189AB4","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29_polarity-pos":"#000000","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29_polarity-neg":"#000000","pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0":"#f20202","pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1":"#189AB4","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0":"#f20202","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1":"#189AB4","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2":"#FF0000","pin-type-component_5102790f-a871-47d9-83fd-2bf45f8f7bb8_0":"#000000","pin-type-component_5102790f-a871-47d9-83fd-2bf45f8f7bb8_1":"#000000","pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0":"#083a36","pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1":"#FF0000","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_0":"#000000","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_1":"#000000","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_2":"#000000","pin-type-component_27363330-fd4d-4d48-8fe5-7e75a0bb5506_0":"#000000","pin-type-component_27363330-fd4d-4d48-8fe5-7e75a0bb5506_1":"#000000","pin-type-component_9cd4866e-171b-4689-8c74-d7df80f41d58_0":"#000000","pin-type-component_9cd4866e-171b-4689-8c74-d7df80f41d58_1":"#000000","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_0":"#000000","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_1":"#000000","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_2":"#000000","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_0":"#000000","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_1":"#000000","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_2":"#000000","pin-type-component_ad1269e6-5014-4c59-af62-685c40e02898_0":"#000000","pin-type-component_ad1269e6-5014-4c59-af62-685c40e02898_1":"#000000","pin-type-component_f533a25e-c11a-427c-a4aa-e80fef74288c_0":"#000000","pin-type-component_f533a25e-c11a-427c-a4aa-e80fef74288c_1":"#000000","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0":"#e75a0d","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1":"#189AB4","pin-type-component_6e804c70-7bd6-41c1-bf62-acd23076114e_0":"#000000","pin-type-component_6e804c70-7bd6-41c1-bf62-acd23076114e_1":"#000000","pin-type-component_dd2abdd4-ed36-4c43-9689-d56c6cb3bd68_0":"#000000","pin-type-component_dd2abdd4-ed36-4c43-9689-d56c6cb3bd68_1":"#000000","pin-type-component_66bf0903-9a55-463b-bc47-49eeb06f5fc3_0":"#000000","pin-type-component_66bf0903-9a55-463b-bc47-49eeb06f5fc3_1":"#000000","pin-type-component_3845c3bd-f40d-4978-9482-daa8afda013f_0":"#000000","pin-type-component_3845c3bd-f40d-4978-9482-daa8afda013f_1":"#000000","pin-type-component_d0b06877-9f19-4217-938d-d5d876016b19_0":"#000000","pin-type-component_d0b06877-9f19-4217-938d-d5d876016b19_1":"#000000","pin-type-component_0db723b4-8ee7-4aa5-8efd-d1c37793e604_0":"#000000","pin-type-component_0db723b4-8ee7-4aa5-8efd-d1c37793e604_1":"#000000","pin-type-component_d2a8b258-269a-4d63-87df-4ce160f1790a_0":"#000000","pin-type-component_d2a8b258-269a-4d63-87df-4ce160f1790a_1":"#000000","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0":"#683D3B","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1":"#e70404","pin-type-component_f4f47a18-edf3-46de-9608-c6b22e0dc54e_0":"#000000","pin-type-component_f4f47a18-edf3-46de-9608-c6b22e0dc54e_1":"#000000"},"pin_to_state":{"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29_polarity-neg":"neutral","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos":"neutral","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_0":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_1":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_2":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_3":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_6":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_7":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_8":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_9":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_10":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_11":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_12":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_13":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_16":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_17":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_19":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_22":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_23":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_24":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_25":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_27":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_28":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_29":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_30":"neutral","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_31":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_1":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_5":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_6":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_7":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_8":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_9":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_10":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_11":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_12":"neutral","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_13":"neutral","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0":"neutral","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1":"neutral","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg":"neutral","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29_polarity-pos":"neutral","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29_polarity-neg":"neutral","pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0":"neutral","pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1":"neutral","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0":"neutral","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1":"neutral","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2":"neutral","pin-type-component_5102790f-a871-47d9-83fd-2bf45f8f7bb8_0":"neutral","pin-type-component_5102790f-a871-47d9-83fd-2bf45f8f7bb8_1":"neutral","pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0":"neutral","pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1":"neutral","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_0":"neutral","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_1":"neutral","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_2":"neutral","pin-type-component_27363330-fd4d-4d48-8fe5-7e75a0bb5506_0":"neutral","pin-type-component_27363330-fd4d-4d48-8fe5-7e75a0bb5506_1":"neutral","pin-type-component_9cd4866e-171b-4689-8c74-d7df80f41d58_0":"neutral","pin-type-component_9cd4866e-171b-4689-8c74-d7df80f41d58_1":"neutral","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_0":"neutral","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_1":"neutral","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_2":"neutral","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_0":"neutral","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_1":"neutral","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_2":"neutral","pin-type-component_ad1269e6-5014-4c59-af62-685c40e02898_0":"neutral","pin-type-component_ad1269e6-5014-4c59-af62-685c40e02898_1":"neutral","pin-type-component_f533a25e-c11a-427c-a4aa-e80fef74288c_0":"neutral","pin-type-component_f533a25e-c11a-427c-a4aa-e80fef74288c_1":"neutral","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0":"neutral","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1":"neutral","pin-type-component_6e804c70-7bd6-41c1-bf62-acd23076114e_0":"neutral","pin-type-component_6e804c70-7bd6-41c1-bf62-acd23076114e_1":"neutral","pin-type-component_dd2abdd4-ed36-4c43-9689-d56c6cb3bd68_0":"neutral","pin-type-component_dd2abdd4-ed36-4c43-9689-d56c6cb3bd68_1":"neutral","pin-type-component_66bf0903-9a55-463b-bc47-49eeb06f5fc3_0":"neutral","pin-type-component_66bf0903-9a55-463b-bc47-49eeb06f5fc3_1":"neutral","pin-type-component_3845c3bd-f40d-4978-9482-daa8afda013f_0":"neutral","pin-type-component_3845c3bd-f40d-4978-9482-daa8afda013f_1":"neutral","pin-type-component_d0b06877-9f19-4217-938d-d5d876016b19_0":"neutral","pin-type-component_d0b06877-9f19-4217-938d-d5d876016b19_1":"neutral","pin-type-component_0db723b4-8ee7-4aa5-8efd-d1c37793e604_0":"neutral","pin-type-component_0db723b4-8ee7-4aa5-8efd-d1c37793e604_1":"neutral","pin-type-component_d2a8b258-269a-4d63-87df-4ce160f1790a_0":"neutral","pin-type-component_d2a8b258-269a-4d63-87df-4ce160f1790a_1":"neutral","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0":"neutral","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1":"neutral","pin-type-component_f4f47a18-edf3-46de-9608-c6b22e0dc54e_0":"neutral","pin-type-component_f4f47a18-edf3-46de-9608-c6b22e0dc54e_1":"neutral"},"next_color_idx":17,"wires_placed_in_order":[["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos"],["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg"],["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28"],["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27"],["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos"],["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-neg"],["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14"],["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15"],["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8"],["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9"],["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5"],["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1"],["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg"],["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos"],["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg"],["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos"],["pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos"],["pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg"],["pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg"],["pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28"],["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0"],["pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos"],["pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16"],["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg"],["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23"],["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg"],["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19"],["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12"],["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11"],["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0"],["pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3"],["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg"],["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17"],["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9"],["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10"],["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg"],["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8"],["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5"],["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg"],["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-neg"],["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1"],["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg"],["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1"],["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg"],["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg"]],"wires_removed_and_placed_in_order":[[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos"]]],[[],[["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg"]]],[[],[["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28"]]],[[],[["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27"]]],[[],[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos"]]],[[],[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-neg"]]],[[],[["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14"]]],[[],[["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15"]]],[[],[["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8"]]],[[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0"]],[]],[[],[["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9"]]],[[],[["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5"]]],[[],[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1"]]],[[],[["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg"]]],[[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos"]],[]],[[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-neg"]],[]],[[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2"]],[]],[[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0"]],[]],[[],[["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos"]]],[[],[["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg"]]],[[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0"]],[]],[[],[["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos"]]],[[],[["pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg"]]],[[],[["pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg"]]],[[],[["pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28"]]],[[],[["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos"]]],[[],[["pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19"]]],[[],[["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12"]]],[[],[["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0"]]],[[],[["pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg"]]],[[],[["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17"]]],[[],[["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9"]]],[[],[["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[],[["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg"]]],[[],[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8"]]],[[],[["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5"]]],[[],[["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg"]]],[[],[["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-neg"]]],[[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1"]],[]],[[],[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1"]]],[[],[]],[[],[]],[[],[]],[[],[]],[[["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg"]],[]],[[],[["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg"]]],[[["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-neg"]],[]],[[],[["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1"]]],[[],[["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg"]]],[[],[["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg"]]]],"arduino_state":"arduino_off","pin_to_uid":{"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg":"0000000000000027","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg":"0000000000000008","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1":"0000000000000026","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg":"0000000000000029","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos":"0000000000000006","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2":"0000000000000028","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg":"0000000000000028","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg":"0000000000000017","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_3_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg":"0000000000000029","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_4_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_4_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_5_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5":"0000000000000007","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6":"0000000000000025","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_6_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_7_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_7_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8":"0000000000000025","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_8_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9":"0000000000000023","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_9_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_10_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_10_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_11_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_11_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_12_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_12_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_13_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_13_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_14_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_14_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_15_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_15_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_16_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_16_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17":"0000000000000022","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_17_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_18_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_18_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_19_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_19_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_20_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_20_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_21_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_21_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_22_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_22_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_23_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_23_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_24_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_24_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_25_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_25_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_26_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_26_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_27_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_27_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_28_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos":"0000000000000002","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg":"0000000000000003","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29_polarity-pos":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_29_polarity-neg":"_","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29":"_","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos":"0000000000000000","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg":"0000000000000001","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_0":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_1":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_2":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_3":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4":"0000000000000000","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5":"0000000000000001","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_6":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_7":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_8":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_9":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_10":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_11":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_12":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_13":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14":"0000000000000004","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15":"0000000000000005","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_16":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_17":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18":"0000000000000016","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_19":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20":"0000000000000018","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21":"0000000000000022","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_22":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_23":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_24":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_25":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26":"0000000000000007","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_27":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_28":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_29":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_30":"_","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_31":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0":"0000000000000002","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_1":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2":"0000000000000003","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3":"0000000000000004","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4":"0000000000000005","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_5":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_6":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_7":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_8":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_9":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_10":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_11":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_12":"_","pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_13":"_","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0":"0000000000000006","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1":"0000000000000007","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2":"0000000000000008","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_0_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_0_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg":"0000000000000021","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_1_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg":"0000000000000027","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_2_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg":"0000000000000017","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3":"0000000000000021","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg":"0000000000000024","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_4_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_5_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_5_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_6_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_6_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7":"0000000000000024","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_7_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_8_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8":"0000000000000020","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos":"0000000000000023","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_9_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10":"0000000000000020","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_10_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_11_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11":"0000000000000020","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos":"0000000000000019","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12":"0000000000000019","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg":"0000000000000015","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_13_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_14_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_14_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15":"0000000000000015","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_15_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16":"0000000000000014","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_16_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_17_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_17_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_18_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_18_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos":"0000000000000013","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19":"0000000000000018","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos":"0000000000000009","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_20_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_21_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_21_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_22_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_22_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23":"0000000000000016","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg":"0000000000000010","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_23_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_24_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_24_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_25_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_25_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_26_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_26_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_27_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_27_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28":"0000000000000012","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_28_polarity-neg":"_","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg":"0000000000000011","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29_polarity-pos":"_","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_1_29_polarity-neg":"_","pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0":"0000000000000012","pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1":"0000000000000011","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0":"0000000000000012","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1":"0000000000000010","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2":"0000000000000009","pin-type-component_5102790f-a871-47d9-83fd-2bf45f8f7bb8_0":"_","pin-type-component_5102790f-a871-47d9-83fd-2bf45f8f7bb8_1":"_","pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0":"0000000000000014","pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1":"0000000000000013","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_0":"_","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_1":"_","pin-type-component_66f8bc17-eb1f-4e67-8117-33c0336c94e1_2":"_","pin-type-component_27363330-fd4d-4d48-8fe5-7e75a0bb5506_0":"_","pin-type-component_27363330-fd4d-4d48-8fe5-7e75a0bb5506_1":"_","pin-type-component_9cd4866e-171b-4689-8c74-d7df80f41d58_0":"_","pin-type-component_9cd4866e-171b-4689-8c74-d7df80f41d58_1":"_","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_0":"_","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_1":"_","pin-type-component_f975c783-09a0-4388-b00b-397fe1665b1b_2":"_","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_0":"_","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_1":"_","pin-type-component_626de387-bf3e-496c-ace3-9cc07bcbcca7_2":"_","pin-type-component_ad1269e6-5014-4c59-af62-685c40e02898_0":"_","pin-type-component_ad1269e6-5014-4c59-af62-685c40e02898_1":"_","pin-type-component_f533a25e-c11a-427c-a4aa-e80fef74288c_0":"_","pin-type-component_f533a25e-c11a-427c-a4aa-e80fef74288c_1":"_","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0":"0000000000000020","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1":"0000000000000021","pin-type-component_6e804c70-7bd6-41c1-bf62-acd23076114e_0":"_","pin-type-component_6e804c70-7bd6-41c1-bf62-acd23076114e_1":"_","pin-type-component_dd2abdd4-ed36-4c43-9689-d56c6cb3bd68_0":"_","pin-type-component_dd2abdd4-ed36-4c43-9689-d56c6cb3bd68_1":"_","pin-type-component_66bf0903-9a55-463b-bc47-49eeb06f5fc3_0":"_","pin-type-component_66bf0903-9a55-463b-bc47-49eeb06f5fc3_1":"_","pin-type-component_3845c3bd-f40d-4978-9482-daa8afda013f_0":"_","pin-type-component_3845c3bd-f40d-4978-9482-daa8afda013f_1":"_","pin-type-component_d0b06877-9f19-4217-938d-d5d876016b19_0":"_","pin-type-component_d0b06877-9f19-4217-938d-d5d876016b19_1":"_","pin-type-component_0db723b4-8ee7-4aa5-8efd-d1c37793e604_0":"_","pin-type-component_0db723b4-8ee7-4aa5-8efd-d1c37793e604_1":"_","pin-type-component_d2a8b258-269a-4d63-87df-4ce160f1790a_0":"_","pin-type-component_d2a8b258-269a-4d63-87df-4ce160f1790a_1":"_","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0":"0000000000000026","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1":"0000000000000025","pin-type-component_f4f47a18-edf3-46de-9608-c6b22e0dc54e_0":"_","pin-type-component_f4f47a18-edf3-46de-9608-c6b22e0dc54e_1":"_"},"component_id_to_pins":{"29e3d5cd-3224-413d-a062-740822a04b1a":["0","1","2","3","4","5","6","7","8","9","10","11","12","13","14","15","16","17","18","19","20","21","22","23","24","25","26","27","28","29","30","31"],"7c6bc105-c394-4a64-9521-bc44ceff98b5":["0","1","2","3","4","5","6","7","8","9","10","11","12","13"],"55a7ce7b-e804-4a1d-a1f9-171e9b277f34":["0","1","2"],"f6061ec8-9e0f-477d-a581-f856789f23b7":["0","1"],"c8450809-2f14-4f14-a78c-76b5cd3da1ad":["0","1","2"],"5102790f-a871-47d9-83fd-2bf45f8f7bb8":["0","1"],"7396e91b-5bcd-46e1-a8f1-738735f2592c":["0","1"],"66f8bc17-eb1f-4e67-8117-33c0336c94e1":["0","1","2"],"27363330-fd4d-4d48-8fe5-7e75a0bb5506":["0","1"],"9cd4866e-171b-4689-8c74-d7df80f41d58":["0","1"],"f975c783-09a0-4388-b00b-397fe1665b1b":["0","1","2"],"626de387-bf3e-496c-ace3-9cc07bcbcca7":["0","1","2"],"ad1269e6-5014-4c59-af62-685c40e02898":["0","1"],"f533a25e-c11a-427c-a4aa-e80fef74288c":["0","1"],"57050f69-0988-4a51-890c-d90af2acaf50":["0","1"],"6e804c70-7bd6-41c1-bf62-acd23076114e":["0","1"],"dd2abdd4-ed36-4c43-9689-d56c6cb3bd68":["0","1"],"66bf0903-9a55-463b-bc47-49eeb06f5fc3":["0","1"],"3845c3bd-f40d-4978-9482-daa8afda013f":["0","1"],"d0b06877-9f19-4217-938d-d5d876016b19":["0","1"],"0db723b4-8ee7-4aa5-8efd-d1c37793e604":["0","1"],"d2a8b258-269a-4d63-87df-4ce160f1790a":["0","1"],"52600675-74b1-4d29-91eb-2baa5606d76d":["0","1"],"f4f47a18-edf3-46de-9608-c6b22e0dc54e":["0","1"]},"uid_to_net":{"_":[],"0000000000000000":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos"],"0000000000000001":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg"],"0000000000000004":["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14"],"0000000000000005":["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15"],"0000000000000007":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5","pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26","pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1"],"0000000000000008":["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg"],"0000000000000002":["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos"],"0000000000000003":["pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg"],"0000000000000006":["pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos"],"0000000000000009":["pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos"],"0000000000000010":["pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg"],"0000000000000011":["pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg"],"0000000000000012":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28","pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0","pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0"],"0000000000000013":["pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos"],"0000000000000014":["pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16"],"0000000000000015":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg"],"0000000000000016":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23"],"0000000000000018":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19"],"0000000000000019":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12"],"0000000000000020":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0","pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10"],"0000000000000021":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3","pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg"],"0000000000000022":["pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17"],"0000000000000023":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9"],"0000000000000024":["pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7","pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg"],"0000000000000025":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8","pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1"],"0000000000000027":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg"],"0000000000000017":["pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg"],"0000000000000026":["pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0","pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1"],"0000000000000028":["pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg"],"0000000000000029":["pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg","pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg"]},"uid_to_text_label":{"0000000000000000":"Net 0","0000000000000001":"Net 1","0000000000000004":"Net 4","0000000000000005":"Net 5","0000000000000007":"Net 7","0000000000000008":"Net 8","0000000000000002":"Net 2","0000000000000003":"Net 3","0000000000000006":"Net 6","0000000000000009":"Net 9","0000000000000010":"Net 10","0000000000000011":"Net 11","0000000000000012":"Net 12","0000000000000013":"Net 13","0000000000000014":"Net 14","0000000000000015":"Net 15","0000000000000016":"Net 16","0000000000000018":"Net 18","0000000000000019":"Net 19","0000000000000020":"Net 20","0000000000000021":"Net 21","0000000000000022":"Net 22","0000000000000023":"Net 23","0000000000000024":"Net 24","0000000000000025":"Net 25","0000000000000027":"Net 27","0000000000000017":"Net 17","0000000000000026":"Net 26","0000000000000028":"Net 28","0000000000000029":"Net 29"},"all_breadboard_info_list":["0daba328-b819-4a1a-a3d8-5e73b2ecc506_30_2_True_685.5_115.5_right","039b408b-a8df-42ed-a12c-4cde63707cd1_30_2_True_685.5_-214.49999999999994_right"],"breadboard_info_list":["0daba328-b819-4a1a-a3d8-5e73b2ecc506_30_2_True_685.5_115.5_right","039b408b-a8df-42ed-a12c-4cde63707cd1_30_2_True_685.5_-214.49999999999994_right"],"componentsData":[{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[666.25,687.5],"typeId":"23db5403-7550-740c-a02b-8b3755757442","componentVersion":1,"instanceId":"29e3d5cd-3224-413d-a062-740822a04b1a","orientation":"up","circleData":[[647.5,830],[662.5,830],[677.5,830],[692.5,830],[707.5,830],[722.5,830],[737.5,830],[752.5,830],[782.5,830],[797.5,830],[812.5,830],[827.5,830],[842.5,830],[857.5,830],[593.5,545],[608.5,545],[623.5,545],[638.5,545],[653.5,545],[668.5,545],[683.5,545],[698.5,545],[713.5,545],[728.5,545],[752.5,545],[767.5,545],[782.5,545],[797.5,545],[812.5,545],[827.5,545],[842.5,545],[857.5,545]],"code":"511,folder,{\"name\":\"sketch\",\"id\":\"150270f7-b12d-4166-be2e-509828e22d68\",\"explorerHtmlId\":\"0569ae18-232c-49e3-be3b-646b8247db87\",\"nameHtmlId\":\"ee0fcf06-ad7d-47bf-9c3d-b2a5b83bcfa2\",\"nameInputHtmlId\":\"ddea2923-1aaf-40e4-98f6-de5db4c57f60\",\"explorerChildHtmlId\":\"53ec99de-33e8-427c-bbde-613cbdc2b11c\",\"explorerCarrotOpenHtmlId\":\"7e532488-8e85-4f3d-a880-e710ae014762\",\"explorerCarrotClosedHtmlId\":\"5e197ce9-fa18-4fc3-8b86-f6cae3f26a51\",\"arduinoBoardFqbn\":\"arduino:avr:uno\",\"arduinoBoardName\":\"\",\"arduinoPortAddress\":\"\"},2,381,file,{\"name\":\"sketch.ino\",\"id\":\"8a5c93f8-f3d8-4e26-8f3e-115506dfd38b\",\"explorerHtmlId\":\"cc5ddb5a-0805-409d-aa3f-eeb5617ebf47\",\"nameHtmlId\":\"147e2f34-bee7-4f33-a4b7-90102166d760\",\"nameInputHtmlId\":\"6346fa8a-6941-4d16-affb-e53e34292ee0\",\"code\":\"void setup() {\\n  // put your setup code here, to run once:\\n\\n}\\n\\nvoid loop() {\\n  // put your main code here, to run repeatedly:\\n\\n}\"},0,252,file,{\"name\":\"documentation.txt\",\"id\":\"72133dff-1840-42c0-9291-56e8010612df\",\"explorerHtmlId\":\"5ad05b0a-e556-4bbb-a5c8-fd446c8b9c2b\",\"nameHtmlId\":\"c6580758-d35c-4bbb-bae4-1304bcad8f38\",\"nameInputHtmlId\":\"3083c783-86a7-4b1e-b0a5-832fa79ccef6\",\"code\":\"\"},0,","codeLabelPosition":[666.25,530],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"1980","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[354.942634,282.5],"typeId":"c2a735ad-a15e-2230-31cf-c702f9ea7cb5","componentVersion":1,"instanceId":"7c6bc105-c394-4a64-9521-bc44ceff98b5","orientation":"up","circleData":[[317.5,320],[332.500012,320],[347.500024,320],[362.500036,320],[377.500048,320],[392.5000585,320],[431.00025999999997,296.21438750000004],[431.0004685,286.76545250000004],[431.00025999999997,277.316726],[431.00025999999997,267.86779250000006],[278.999632,268.55597750000004],[278.9994235,278.004752],[278.999632,287.4535265],[278.999632,296.9022995]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1021.6797835,246.77594000000005],"typeId":"5eb4ee00-1bfb-4094-b0b7-76a195dc2829","componentVersion":7,"instanceId":"55a7ce7b-e804-4a1d-a1f9-171e9b277f34","orientation":"up","circleData":[[1007.5,320],[1021.3190215,320.454302],[1036.1842344999998,320.9489255]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[242.2312435,-24.50060499999995],"typeId":"75a91b20-33fe-4043-8d25-b0ca953a6307","componentVersion":3,"instanceId":"f6061ec8-9e0f-477d-a581-f856789f23b7","orientation":"right","circleData":[[392.5,-70],[392.50000000000006,-54.3574795]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[588.4745245,-281.92794549999996],"typeId":"1e489b6c-0e9c-4f1b-98f8-b8590afb7732","componentVersion":1,"instanceId":"c8450809-2f14-4f14-a78c-76b5cd3da1ad","orientation":"up","circleData":[[557.5,-189.99999999999997],[587.5,-189.99999999999997],[617.5,-189.99999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Capacitance":{"type":"double","name":"Capacitance","value":"2.2e-7","unit":"F","showOnComp":true,"required":true}},"position":[588.3404767320466,-52.59148187187603],"typeId":"2c229afa-5375-44c6-9069-3781267c16db","componentVersion":1,"instanceId":"5102790f-a871-47d9-83fd-2bf45f8f7bb8","orientation":"up","circleData":[[542.5,-39.99999999999995],[617.5000000000002,-39.99999999999995]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[784.616947,-266.63191149999994],"typeId":"a0726024-2717-468d-bcb0-1ef57233b392","componentVersion":3,"instanceId":"7396e91b-5bcd-46e1-a8f1-738735f2592c","orientation":"up","circleData":[[707.5,-174.99999999999994],[670,-174.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"976","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[706.747,-99.01224999999985],"typeId":"bf357ed6-dccd-a67c-b3c8-1a96cf58f9a4","componentVersion":1,"instanceId":"66f8bc17-eb1f-4e67-8117-33c0336c94e1","orientation":"up","circleData":[[692.5,-54.99999999999994],[707.497003,-54.99999999999994],[722.4940015,-54.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"type":"double","name":"Resistance","value":"220","unit":"Ω","showOnComp":true,"required":true,"validRange":[0,9007199254740991]},"Tolerance":{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},"Number Of Bands":{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}},"position":[648.4322648810503,-24.999999999999947],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"27363330-fd4d-4d48-8fe5-7e75a0bb5506","orientation":"up","circleData":[[602.5,-24.999999999999947],[677.5,-24.999999999999947]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[684.16975,-121.70724999999999],"typeId":"82d731d1-c75f-e131-c68f-ff0e81dc6210","componentVersion":1,"instanceId":"9cd4866e-171b-4689-8c74-d7df80f41d58","orientation":"up","circleData":[[677.5,-39.99999999999994],[692.5045,-39.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"976","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[766.7470000000001,-9.012249999999952],"typeId":"bf357ed6-dccd-a67c-b3c8-1a96cf58f9a4","componentVersion":1,"instanceId":"f975c783-09a0-4388-b00b-397fe1665b1b","orientation":"up","circleData":[[752.5,35.000000000000036],[767.4970030000002,35.000000000000036],[782.4940015,35.000000000000036]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"976","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[811.7470000000001,215.98774999999995],"typeId":"bf357ed6-dccd-a67c-b3c8-1a96cf58f9a4","componentVersion":1,"instanceId":"626de387-bf3e-496c-ace3-9cc07bcbcca7","orientation":"up","circleData":[[797.5,259.9999999999999],[812.4970030000002,259.9999999999999],[827.4940015,259.9999999999999]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[744.16975,-31.707250000000037],"typeId":"82d731d1-c75f-e131-c68f-ff0e81dc6210","componentVersion":1,"instanceId":"ad1269e6-5014-4c59-af62-685c40e02898","orientation":"up","circleData":[[737.5,50.00000000000001],[752.5045,50.00000000000001]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"type":"double","name":"Resistance","value":"220","unit":"Ω","showOnComp":true,"required":true,"validRange":[0,9007199254740991]},"Tolerance":{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},"Number Of Bands":{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}},"position":[708.4322648810503,65],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"f533a25e-c11a-427c-a4aa-e80fef74288c","orientation":"up","circleData":[[662.5,65],[737.5,65]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"711","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[1312.6375,54.765546500000006],"typeId":"bd390fed-95a0-8dd4-98ea-cc81efdfc30b","componentVersion":1,"instanceId":"57050f69-0988-4a51-890c-d90af2acaf50","orientation":"up","circleData":[[1187.5,50.00000000000002],[1187.5,65.59140950000003]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Capacitance":{"type":"double","name":"Capacitance","value":"2.2e-7","unit":"F","showOnComp":true,"required":true}},"position":[873.3404767320467,22.40851812812395],"typeId":"2c229afa-5375-44c6-9069-3781267c16db","componentVersion":1,"instanceId":"6e804c70-7bd6-41c1-bf62-acd23076114e","orientation":"up","circleData":[[827.5,35.000000000000036],[902.5000000000002,35.000000000000036]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[854.2614504999999,94.93749950000006],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"dd2abdd4-ed36-4c43-9689-d56c6cb3bd68","orientation":"up","circleData":[[827.5,95],[902.5,95]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[789.16975,193.2927499999998],"typeId":"82d731d1-c75f-e131-c68f-ff0e81dc6210","componentVersion":1,"instanceId":"66bf0903-9a55-463b-bc47-49eeb06f5fc3","orientation":"up","circleData":[[782.5,275],[797.5045,275]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"Resistance":{"type":"double","name":"Resistance","value":"220","unit":"Ω","showOnComp":true,"required":true,"validRange":[0,9007199254740991]},"Tolerance":{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},"Number Of Bands":{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}},"position":[738.4322648810503,290],"typeId":"72c75556-baa3-04e7-55a5-e13f447c8c5a","componentVersion":1,"instanceId":"3845c3bd-f40d-4978-9482-daa8afda013f","orientation":"up","circleData":[[692.5,290],[767.5,290]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[804.16975,-151.70725],"typeId":"82d731d1-c75f-e131-c68f-ff0e81dc6210","componentVersion":1,"instanceId":"d0b06877-9f19-4217-938d-d5d876016b19","orientation":"up","circleData":[[797.5,-69.99999999999997],[812.5045,-69.99999999999997]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[819.16975,-136.70724999999993],"typeId":"82d731d1-c75f-e131-c68f-ff0e81dc6210","componentVersion":1,"instanceId":"0db723b4-8ee7-4aa5-8efd-d1c37793e604","orientation":"up","circleData":[[812.5,-54.99999999999994],[827.5045,-54.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[834.16975,-121.70724999999993],"typeId":"82d731d1-c75f-e131-c68f-ff0e81dc6210","componentVersion":1,"instanceId":"d2a8b258-269a-4d63-87df-4ce160f1790a","orientation":"up","circleData":[[827.5,-39.99999999999994],[842.5045,-39.99999999999994]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{},"position":[1353.337777,282.3988715000001],"typeId":"6635379e-9371-f184-7e48-a00d3644b40e","componentVersion":1,"instanceId":"52600675-74b1-4d29-91eb-2baa5606d76d","orientation":"up","circleData":[[1202.5,395],[1202.552413,381.733166]],"cirkitStudioVersion":"1.3.3"},{"compProperties":{"mpn":{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},"manufacturer":{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}},"position":[884.2614504999999,289.93749950000006],"typeId":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","componentVersion":1,"instanceId":"f4f47a18-edf3-46de-9608-c6b22e0dc54e","orientation":"up","circleData":[[857.5,290],[932.5,290]],"cirkitStudioVersion":"1.3.3"}],"bounds":{"top":"-389.54555","left":"75.87034","width":"1464.63281","height":"1244.54555","x":"75.87034","y":"-389.54555"},"cachedBreadboardPrettyViewWires":["{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos\",\"rawStartPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_4\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"707.5000000000_830.0000000000\\\",\\\"707.5000000000_875.0000000000\\\",\\\"400.0000000000_875.0000000000\\\",\\\"400.0000000000_470.0000000000\\\",\\\"512.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg\",\"rawStartPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_5\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_29_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"722.5000000000_830.0000000000\\\",\\\"722.5000000000_860.0000000000\\\",\\\"422.5000000000_860.0000000000\\\",\\\"422.5000000000_485.0000000000\\\",\\\"512.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#0E4CA1\",\"startPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14\",\"endPinId\":\"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3\",\"rawStartPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_14\",\"rawEndPinId\":\"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_3\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"593.5000000000_545.0000000000\\\",\\\"593.5000000000_425.0000000000\\\",\\\"362.5000360000_425.0000000000\\\",\\\"362.5000360000_320.0000000000\\\"]}\"}","{\"color\":\"#FFE502\",\"startPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15\",\"endPinId\":\"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4\",\"rawStartPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_15\",\"rawEndPinId\":\"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_4\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"608.5000000000_545.0000000000\\\",\\\"608.5000000000_417.5000000000\\\",\\\"377.5000480000_417.5000000000\\\",\\\"377.5000480000_320.0000000000\\\"]}\"}","{\"color\":\"#e2e600\",\"startPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5\",\"endPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_4\",\"rawEndPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_26\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_425.0000000000\\\",\\\"872.5000000000_515.0000000000\\\",\\\"782.5000000000_515.0000000000\\\",\\\"782.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#e2e600\",\"startPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5\",\"endPinId\":\"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_5_0\",\"rawEndPinId\":\"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"872.5000000000_365.0000000000\\\",\\\"872.5000000000_342.5000000000\\\",\\\"1021.3190215000_342.5000000000\\\",\\\"1021.3190215000_320.4543020000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg\",\"rawStartPinId\":\"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_2\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_0_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1036.1842345000_320.9489255000\\\",\\\"1036.1842345000_335.0000000000\\\",\\\"1037.5000000000_335.0000000000\\\",\\\"1037.5000000000_485.0000000000\\\",\\\"947.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos\",\"rawStartPinId\":\"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_0\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"317.5000000000_320.0000000000\\\",\\\"317.5000000000_440.0000000000\\\",\\\"527.5000000000_440.0000000000\\\",\\\"527.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg\",\"rawStartPinId\":\"pin-type-component_7c6bc105-c394-4a64-9521-bc44ceff98b5_2\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_28_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"347.5000240000_320.0000000000\\\",\\\"347.5000240000_455.0000000000\\\",\\\"527.5000000000_455.0000000000\\\",\\\"527.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos\",\"rawStartPinId\":\"pin-type-component_55a7ce7b-e804-4a1d-a1f9-171e9b277f34_0\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_1_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"1007.5000000000_320.0000000000\\\",\\\"1007.5000000000_432.5000000000\\\",\\\"932.5000000000_432.5000000000\\\",\\\"932.5000000000_470.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos\",\"rawStartPinId\":\"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_2\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_20_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"617.5000000000_-190.0000000000\\\",\\\"617.5000000000_-160.0000000000\\\",\\\"647.5000000000_-160.0000000000\\\",\\\"647.5000000000_-130.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg\",\"rawStartPinId\":\"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_1\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"587.5000000000_-190.0000000000\\\",\\\"587.5000000000_-160.0000000000\\\",\\\"602.5000000000_-160.0000000000\\\",\\\"602.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg\",\"rawStartPinId\":\"pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_1\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_29_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"392.5000000000_-54.3574795000\\\",\\\"422.5000000000_-54.3574795000\\\",\\\"422.5000000000_-115.0000000000\\\",\\\"512.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#f20202\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28\",\"endPinId\":\"pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_0\",\"rawEndPinId\":\"pin-type-component_f6061ec8-9e0f-477d-a581-f856789f23b7_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"527.5000000000_-70.0000000000\\\",\\\"392.5000000000_-70.0000000000\\\"]}\"}","{\"color\":\"#f20202\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28\",\"endPinId\":\"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_0_28_1\",\"rawEndPinId\":\"pin-type-component_c8450809-2f14-4f14-a78c-76b5cd3da1ad_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"527.5000000000_-55.0000000000\\\",\\\"557.5000000000_-55.0000000000\\\",\\\"557.5000000000_-190.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos\",\"rawStartPinId\":\"pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_1\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_19_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"670.0000000000_-175.0000000000\\\",\\\"662.5000000000_-175.0000000000\\\",\\\"662.5000000000_-130.0000000000\\\"]}\"}","{\"color\":\"#083a36\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16\",\"endPinId\":\"pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_0_16_0\",\"rawEndPinId\":\"pin-type-component_7396e91b-5bcd-46e1-a8f1-738735f2592c_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"707.5000000000_-70.0000000000\\\",\\\"700.0000000000_-70.0000000000\\\",\\\"700.0000000000_-175.0000000000\\\",\\\"707.5000000000_-175.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_0_15_2\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_13_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"722.5000000000_-40.0000000000\\\",\\\"752.5000000000_-40.0000000000\\\",\\\"752.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#5ecd13\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23\",\"endPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_0_23_4\",\"rawEndPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_18\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"602.5000000000_-10.0000000000\\\",\\\"602.5000000000_515.0000000000\\\",\\\"653.5000000000_515.0000000000\\\",\\\"653.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#14db25\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19\",\"endPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_1_19_3\",\"rawEndPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_20\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"662.5000000000_80.0000000000\\\",\\\"662.5000000000_515.0000000000\\\",\\\"683.5000000000_515.0000000000\\\",\\\"683.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_1_12_1\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_12_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"767.5000000000_50.0000000000\\\",\\\"767.5000000000_-130.0000000000\\\"]}\"}","{\"color\":\"#e75a0d\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8\",\"endPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_1\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_50.0000000000\\\",\\\"782.5000000000_50.0000000000\\\"]}\"}","{\"color\":\"#e75a0d\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8\",\"endPinId\":\"pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_1_8_2\",\"rawEndPinId\":\"pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"827.5000000000_65.0000000000\\\",\\\"827.5000000000_80.0000000000\\\",\\\"1172.5000000000_80.0000000000\\\",\\\"1172.5000000000_50.0000000000\\\",\\\"1187.5000000000_50.0000000000\\\"]}\"}","{\"color\":\"#e75a0d\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10\",\"endPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_0_10_1\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_1_11_2\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"797.5000000000_-55.0000000000\\\",\\\"797.5000000000_65.0000000000\\\",\\\"782.5000000000_65.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3\",\"endPinId\":\"pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_2\",\"rawEndPinId\":\"pin-type-component_57050f69-0988-4a51-890c-d90af2acaf50_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_65.0000000000\\\",\\\"1172.5000000000_65.0000000000\\\",\\\"1172.5000000000_65.5914095000\\\",\\\"1187.5000000000_65.5914095000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_1_3_1\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_1_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_50.0000000000\\\",\\\"932.5000000000_50.0000000000\\\",\\\"932.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#1ddd03\",\"startPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17\",\"endPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_17_3\",\"rawEndPinId\":\"pin-type-component_29e3d5cd-3224-413d-a062-740822a04b1a_21\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"692.5000000000_305.0000000000\\\",\\\"692.5000000000_515.0000000000\\\",\\\"698.5000000000_515.0000000000\\\",\\\"698.5000000000_545.0000000000\\\"]}\"}","{\"color\":\"#FF0000\",\"startPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_9_1\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_9_polarity-pos\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"812.5000000000_275.0000000000\\\",\\\"812.5000000000_-130.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7\",\"endPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_039b408b-a8df-42ed-a12c-4cde63707cd1_0_7_3\",\"rawEndPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_4_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"842.5000000000_-25.0000000000\\\",\\\"887.5000000000_-25.0000000000\\\",\\\"887.5000000000_-115.0000000000\\\"]}\"}","{\"color\":\"#e70404\",\"startPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6\",\"endPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_1\",\"rawEndPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_8_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"857.5000000000_275.0000000000\\\",\\\"827.5000000000_275.0000000000\\\"]}\"}","{\"color\":\"#e70404\",\"startPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6\",\"endPinId\":\"pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_6_0\",\"rawEndPinId\":\"pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_1\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"857.5000000000_260.0000000000\\\",\\\"857.5000000000_177.5000000000\\\",\\\"1157.5000000000_177.5000000000\\\",\\\"1157.5000000000_381.7331660000\\\",\\\"1202.5524130000_381.7331660000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg\",\"rawStartPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_2_polarity-neg\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_0_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"917.5000000000_-115.0000000000\\\",\\\"1015.0000000000_-115.0000000000\\\",\\\"1015.0000000000_215.0000000000\\\",\\\"947.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg\",\"rawStartPinId\":\"pin-type-power-rail_039b408b-a8df-42ed-a12c-4cde63707cd1_0_3_polarity-neg\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_2_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"902.5000000000_-115.0000000000\\\",\\\"1097.5000000000_-115.0000000000\\\",\\\"1097.5000000000_485.0000000000\\\",\\\"917.5000000000_485.0000000000\\\"]}\"}","{\"color\":\"#683D3B\",\"startPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1\",\"endPinId\":\"pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_3\",\"rawEndPinId\":\"pin-type-component_52600675-74b1-4d29-91eb-2baa5606d76d_0\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"932.5000000000_305.0000000000\\\",\\\"1157.5000000000_305.0000000000\\\",\\\"1157.5000000000_395.0000000000\\\",\\\"1202.5000000000_395.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-breadboard_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg\",\"rawStartPinId\":\"pin-type-breadboard-sub-pin_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_1\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_2_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"917.5000000000_275.0000000000\\\",\\\"917.5000000000_215.0000000000\\\"]}\"}","{\"color\":\"#189AB4\",\"startPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg\",\"endPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg\",\"rawStartPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_0_1_polarity-neg\",\"rawEndPinId\":\"pin-type-power-rail_0daba328-b819-4a1a-a3d8-5e73b2ecc506_1_3_polarity-neg\",\"pointPath\":\"{\\\"listOfPointStrings\\\":[\\\"932.5000000000_215.0000000000\\\",\\\"932.5000000000_350.0000000000\\\",\\\"902.5000000000_350.0000000000\\\",\\\"902.5000000000_485.0000000000\\\"]}\"}"],"projectDescription":""}PK
     B"BY               jsons/PK
     B"BY�h���`  �`     jsons/user_defined.json{"type":"user_defined","version":"0.0.1","subtypes":[{"subtypeName":"Arduino UNO","category":["Microcontroller"],"userDefined":false,"id":"23db5403-7550-740c-a02b-8b3755757442","subtypeDescription":"","subtypePic":"0b351edc-7875-4477-b820-546ce15be531.png","fqbn":"arduino:avr:uno","pinInfo":{"numDisplayCols":"29.5","numDisplayRows":"21","pins":[{"uniquePinIdString":"0","positionMil":"1350,100","isAnchorPin":true,"label":"UNUSED"},{"uniquePinIdString":"1","positionMil":"1450,100","isAnchorPin":false,"label":"IOREF"},{"uniquePinIdString":"2","positionMil":"1550,100","isAnchorPin":false,"label":"Reset"},{"uniquePinIdString":"3","positionMil":"1650,100","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"4","positionMil":"1750,100","isAnchorPin":false,"label":"5V"},{"uniquePinIdString":"5","positionMil":"1850,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"6","positionMil":"1950,100","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"2050,100","isAnchorPin":false,"label":"Vin"},{"uniquePinIdString":"8","positionMil":"2250,100","isAnchorPin":false,"label":"A0"},{"uniquePinIdString":"9","positionMil":"2350,100","isAnchorPin":false,"label":"A1"},{"uniquePinIdString":"10","positionMil":"2450,100","isAnchorPin":false,"label":"A2"},{"uniquePinIdString":"11","positionMil":"2550,100","isAnchorPin":false,"label":"A3"},{"uniquePinIdString":"12","positionMil":"2650,100","isAnchorPin":false,"label":"A4"},{"uniquePinIdString":"13","positionMil":"2750,100","isAnchorPin":false,"label":"A5"},{"uniquePinIdString":"14","positionMil":"990,2000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"15","positionMil":"1090,2000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"16","positionMil":"1190,2000","isAnchorPin":false,"label":"AREF"},{"uniquePinIdString":"17","positionMil":"1290,2000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"18","positionMil":"1390,2000","isAnchorPin":false,"label":"D13"},{"uniquePinIdString":"19","positionMil":"1490,2000","isAnchorPin":false,"label":"D12"},{"uniquePinIdString":"20","positionMil":"1590,2000","isAnchorPin":false,"label":"D11"},{"uniquePinIdString":"21","positionMil":"1690,2000","isAnchorPin":false,"label":"D10"},{"uniquePinIdString":"22","positionMil":"1790,2000","isAnchorPin":false,"label":"D9"},{"uniquePinIdString":"23","positionMil":"1890,2000","isAnchorPin":false,"label":"D8"},{"uniquePinIdString":"24","positionMil":"2050,2000","isAnchorPin":false,"label":"D7"},{"uniquePinIdString":"25","positionMil":"2150,2000","isAnchorPin":false,"label":"D6"},{"uniquePinIdString":"26","positionMil":"2250,2000","isAnchorPin":false,"label":"D5"},{"uniquePinIdString":"27","positionMil":"2350,2000","isAnchorPin":false,"label":"D4"},{"uniquePinIdString":"28","positionMil":"2450,2000","isAnchorPin":false,"label":"D3"},{"uniquePinIdString":"29","positionMil":"2550,2000","isAnchorPin":false,"label":"D2"},{"uniquePinIdString":"30","positionMil":"2650,2000","isAnchorPin":false,"label":"D1"},{"uniquePinIdString":"31","positionMil":"2750,2000","isAnchorPin":false,"label":"D0"}],"pinType":"wired"},"iconPic":"e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png","properties":[{"type":"string","name":"mpn","value":"A000066","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Arduino","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Adafruit TSL2591 High Dynamic Range Digital Light Sensor","category":["Adafruit"],"userDefined":false,"id":"c2a735ad-a15e-2230-31cf-c702f9ea7cb5","subtypeDescription":"","subtypePic":"e28c3bbb-5472-4456-9ec9-e60c5bfdece2.png","pinInfo":{"numDisplayCols":"10.72630","numDisplayRows":"7.00000","pins":[{"uniquePinIdString":"0","positionMil":"286.69744,100.00000","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"386.69752,100.00000","isAnchorPin":false,"label":"3.3V"},{"uniquePinIdString":"2","positionMil":"486.69760,100.00000","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"3","positionMil":"586.69768,100.00000","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"4","positionMil":"686.69776,100.00000","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"5","positionMil":"786.69783,100.00000","isAnchorPin":false,"label":"INT"},{"uniquePinIdString":"6","positionMil":"1043.36584,258.57075","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"7","positionMil":"1043.36723,321.56365","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"8","positionMil":"1043.36584,384.55516","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"9","positionMil":"1043.36584,447.54805","isAnchorPin":false,"label":"SCL"},{"uniquePinIdString":"10","positionMil":"30.02832,442.96015","isAnchorPin":false,"label":"GND"},{"uniquePinIdString":"11","positionMil":"30.02693,379.96832","isAnchorPin":false,"label":"VCC"},{"uniquePinIdString":"12","positionMil":"30.02832,316.97649","isAnchorPin":false,"label":"SDA"},{"uniquePinIdString":"13","positionMil":"30.02832,253.98467","isAnchorPin":false,"label":"SCL"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"1980","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"9a88a734-d46c-4092-86bc-e9f7b966a1ec.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"KY-015 DHT11","category":["User Defined"],"id":"5eb4ee00-1bfb-4094-b0b7-76a195dc2829","componentVersion":7,"userDefined":true,"subtypeDescription":"","subtypePic":"05596fff-4f8f-4556-8b1d-73ff55b6eaa8.png","iconPic":"e4b09d94-725a-4fc8-8861-adc4f6b1a3b4.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"5.51599","numDisplayRows":"9.68775","pins":[{"uniquePinIdString":"0","positionMil":"181.26761,-3.77290","isAnchorPin":true,"label":"5V"},{"uniquePinIdString":"1","positionMil":"273.39442,-6.80158","isAnchorPin":false,"label":"S"},{"uniquePinIdString":"2","positionMil":"372.49584,-10.09907","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Battery AAx5 7.5V","category":["User Defined"],"id":"75a91b20-33fe-4043-8d25-b0ca953a6307","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"c49304c6-1828-42f7-9c78-6513b79a7c1a.png","iconPic":"86ae6a4b-562d-4e93-9595-3c4b0d09f42e.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"26.75693","numDisplayRows":"20.84812","pins":[{"uniquePinIdString":"0","positionMil":"1034.51720,2044.19771","isAnchorPin":true,"label":"VCC"},{"uniquePinIdString":"1","positionMil":"1138.80067,2044.19771","isAnchorPin":false,"label":"GND"}],"pinType":"wired"},"properties":[]},{"subtypeName":"7805","category":["User Defined"],"id":"1e489b6c-0e9c-4f1b-98f8-b8590afb7732","componentVersion":1,"userDefined":true,"subtypeDescription":"","subtypePic":"43e4be74-284e-4582-91bd-e4a77387caa5.png","iconPic":"a3b4885c-2487-4906-a080-ee9b44acb175.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"6.46327","numDisplayRows":"13.01568","pins":[{"uniquePinIdString":"0","positionMil":"116.66667,37.93103","isAnchorPin":true,"label":"Vin"},{"uniquePinIdString":"1","positionMil":"316.66667,37.93103","isAnchorPin":false,"label":"Gnd"},{"uniquePinIdString":"2","positionMil":"516.66667,37.93103","isAnchorPin":false,"label":"Vout"}],"pinType":"wired"},"properties":[]},{"subtypeName":"Ceramic Capacitor","subtypeDescription":"","id":"2c229afa-5375-44c6-9069-3781267c16db","subtypePic":"7c9bed20-c7d7-43dc-b689-820375f46db8.png","category":["Basic"],"userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"44.10000,0.00000","endPositionMil":"44.10000,-200.00000","isAnchorPin":true,"label":"pin0"},{"uniquePinIdString":"1","startPositionMil":"144.33000,0.00000","endPositionMil":"144.33000,-200.00000","isAnchorPin":false,"label":"pin1"}],"numDisplayCols":"1.88360","numDisplayRows":"2.48270","pinType":"movable"},"properties":[{"type":"double","name":"Capacitance","value":"0.0000001","unit":"F","showOnComp":true,"required":true}],"iconPic":"7ade412b-fa94-47ea-987a-d6c9baa14438.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Humidifier","category":["User Defined"],"id":"a0726024-2717-468d-bcb0-1ef57233b392","componentVersion":3,"userDefined":true,"subtypeDescription":"","subtypePic":"4d53c106-8e41-4afb-b8f1-56dd58def1e6.png","iconPic":"d004afae-d6a3-4a65-a5d4-4f8d37106046.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"16.13983","numDisplayRows":"13.88119","pins":[{"uniquePinIdString":"0","positionMil":"292.87852,83.18009","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"42.87852,83.18009","isAnchorPin":false,"label":"5V"}],"pinType":"wired"},"properties":[]},{"subtypeName":"TIP120 Hi-Current Darlington Transistor","category":["Adafruit"],"userDefined":false,"id":"bf357ed6-dccd-a67c-b3c8-1a96cf58f9a4","subtypeDescription":"","subtypePic":"19f08d4b-a68c-4e36-96dd-32682874608f.png","pinInfo":{"numDisplayCols":"3.69980","numDisplayRows":"6.23170","pins":[{"uniquePinIdString":"0","positionMil":"90.01000,18.17000","isAnchorPin":true,"label":"BASE"},{"uniquePinIdString":"1","positionMil":"189.99002,18.17000","isAnchorPin":false,"label":"COLLECTOR"},{"uniquePinIdString":"2","positionMil":"289.97001,18.17000","isAnchorPin":false,"label":"EMITTER"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"976","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"5779bcfa-264f-4061-b24b-5c8b50561781.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LED: Two Pin (red)","subtypeDescription":"","id":"82d731d1-c75f-e131-c68f-ff0e81dc6210","category":["Output"],"userDefined":false,"subtypePic":"da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"62.87000,0.00000","endPositionMil":"62.87000,-341.89000","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"162.90000,0.00000","endPositionMil":"162.90000,-341.89000","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"2.14670","numDisplayRows":"4.05650","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"b96c8ad8-7845-422d-b49f-326b2968fdb8.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"TIP120 Hi-Current Darlington Transistor","category":["Adafruit"],"userDefined":false,"id":"bf357ed6-dccd-a67c-b3c8-1a96cf58f9a4","subtypeDescription":"","subtypePic":"19f08d4b-a68c-4e36-96dd-32682874608f.png","pinInfo":{"numDisplayCols":"3.69980","numDisplayRows":"6.23170","pins":[{"uniquePinIdString":"0","positionMil":"90.01000,18.17000","isAnchorPin":true,"label":"BASE"},{"uniquePinIdString":"1","positionMil":"189.99002,18.17000","isAnchorPin":false,"label":"COLLECTOR"},{"uniquePinIdString":"2","positionMil":"289.97001,18.17000","isAnchorPin":false,"label":"EMITTER"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"976","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"5779bcfa-264f-4061-b24b-5c8b50561781.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"TIP120 Hi-Current Darlington Transistor","category":["Adafruit"],"userDefined":false,"id":"bf357ed6-dccd-a67c-b3c8-1a96cf58f9a4","subtypeDescription":"","subtypePic":"19f08d4b-a68c-4e36-96dd-32682874608f.png","pinInfo":{"numDisplayCols":"3.69980","numDisplayRows":"6.23170","pins":[{"uniquePinIdString":"0","positionMil":"90.01000,18.17000","isAnchorPin":true,"label":"BASE"},{"uniquePinIdString":"1","positionMil":"189.99002,18.17000","isAnchorPin":false,"label":"COLLECTOR"},{"uniquePinIdString":"2","positionMil":"289.97001,18.17000","isAnchorPin":false,"label":"EMITTER"}],"pinType":"wired"},"properties":[{"type":"string","name":"mpn","value":"976","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"5779bcfa-264f-4061-b24b-5c8b50561781.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LED: Two Pin (red)","subtypeDescription":"","id":"82d731d1-c75f-e131-c68f-ff0e81dc6210","category":["Output"],"userDefined":false,"subtypePic":"da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"62.87000,0.00000","endPositionMil":"62.87000,-341.89000","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"162.90000,0.00000","endPositionMil":"162.90000,-341.89000","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"2.14670","numDisplayRows":"4.05650","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"b96c8ad8-7845-422d-b49f-326b2968fdb8.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"DC Motor","category":["Output"],"userDefined":false,"id":"bd390fed-95a0-8dd4-98ea-cc81efdfc30b","subtypeDescription":"","subtypePic":"f1393e3f-31c1-44d6-9d33-bf195c230c11.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"27.77778,432.60397","endPositionMil":"0.00000,418.71531","isAnchorPin":true,"label":"pin 1"},{"uniquePinIdString":"1","startPositionMil":"27.77778,314.77258","endPositionMil":"0.00000,314.77258","isAnchorPin":false,"label":"pin 2"}],"numDisplayCols":"16.68500","numDisplayRows":"7.73890","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"711","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Adafruit Industries","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"1ff35573-e276-4514-8c59-6294c96ecf57.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Ceramic Capacitor","subtypeDescription":"","id":"2c229afa-5375-44c6-9069-3781267c16db","subtypePic":"7c9bed20-c7d7-43dc-b689-820375f46db8.png","category":["Basic"],"userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"44.10000,0.00000","endPositionMil":"44.10000,-200.00000","isAnchorPin":true,"label":"pin0"},{"uniquePinIdString":"1","startPositionMil":"144.33000,0.00000","endPositionMil":"144.33000,-200.00000","isAnchorPin":false,"label":"pin1"}],"numDisplayCols":"1.88360","numDisplayRows":"2.48270","pinType":"movable"},"properties":[{"type":"double","name":"Capacitance","value":"0.0000001","unit":"F","showOnComp":true,"required":true}],"iconPic":"7ade412b-fa94-47ea-987a-d6c9baa14438.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LED: Two Pin (red)","subtypeDescription":"","id":"82d731d1-c75f-e131-c68f-ff0e81dc6210","category":["Output"],"userDefined":false,"subtypePic":"da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"62.87000,0.00000","endPositionMil":"62.87000,-341.89000","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"162.90000,0.00000","endPositionMil":"162.90000,-341.89000","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"2.14670","numDisplayRows":"4.05650","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"b96c8ad8-7845-422d-b49f-326b2968fdb8.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Resistor","category":["Basic"],"id":"72c75556-baa3-04e7-55a5-e13f447c8c5a","subtypeDescription":"","subtypePic":"bbfae99c-8036-4c5e-89fd-a87441410720.png","userDefined":false,"pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"-120.00000,50.00000","endPositionMil":"-250.00000,50.00000","isAnchorPin":true,"label":"pin1"},{"uniquePinIdString":"1","startPositionMil":"120.00000,50.00000","endPositionMil":"250.00000,50.00000","isAnchorPin":false,"label":"pin2"}],"numDisplayCols":"0","numDisplayRows":"1","pinType":"movable"},"properties":[{"type":"double","name":"Resistance","value":200,"unit":"Ω","showOnComp":true,"required":true,"validRange":[0,70000]},{"type":"dropdown","name":"Tolerance","value":"5%","options":["0.25%","0.1%","0.5%","1%","2%","5%","10%"],"showOnComp":false,"required":true},{"type":"dropdown","name":"Number Of Bands","value":5,"options":[4,5,6],"showOnComp":false,"required":true}],"iconPic":"a262aa33-74c4-460b-b0ad-c746896f6744.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LED: Two Pin (red)","subtypeDescription":"","id":"82d731d1-c75f-e131-c68f-ff0e81dc6210","category":["Output"],"userDefined":false,"subtypePic":"da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"62.87000,0.00000","endPositionMil":"62.87000,-341.89000","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"162.90000,0.00000","endPositionMil":"162.90000,-341.89000","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"2.14670","numDisplayRows":"4.05650","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"b96c8ad8-7845-422d-b49f-326b2968fdb8.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LED: Two Pin (red)","subtypeDescription":"","id":"82d731d1-c75f-e131-c68f-ff0e81dc6210","category":["Output"],"userDefined":false,"subtypePic":"da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"62.87000,0.00000","endPositionMil":"62.87000,-341.89000","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"162.90000,0.00000","endPositionMil":"162.90000,-341.89000","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"2.14670","numDisplayRows":"4.05650","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"b96c8ad8-7845-422d-b49f-326b2968fdb8.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"LED: Two Pin (red)","subtypeDescription":"","id":"82d731d1-c75f-e131-c68f-ff0e81dc6210","category":["Output"],"userDefined":false,"subtypePic":"da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"62.87000,0.00000","endPositionMil":"62.87000,-341.89000","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"162.90000,0.00000","endPositionMil":"162.90000,-341.89000","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"2.14670","numDisplayRows":"4.05650","pinType":"movable"},"properties":[{"type":"string","name":"mpn","value":"HLMP-3762","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"Broadcom","unit":"","showOnComp":false,"userVisible":false,"required":true}],"iconPic":"b96c8ad8-7845-422d-b49f-326b2968fdb8.png","componentVersion":1,"imageLocation":"local_cache"},{"subtypeName":"Fan","category":["Output"],"userDefined":true,"id":"6635379e-9371-f184-7e48-a00d3644b40e","subtypeDescription":"","subtypePic":"146a6d58-0553-42c9-b8c7-03425202d69a.png","iconPic":"d1a57a69-e5a0-4805-bdaf-8d975fdf5bdb.png","imageLocation":"local_cache","pinInfo":{"numDisplayCols":"23.62205","numDisplayRows":"19.68504","pins":[{"uniquePinIdString":"0","positionMil":"175.51732,233.57781","isAnchorPin":true,"label":"GND"},{"uniquePinIdString":"1","positionMil":"175.86674,322.02337","isAnchorPin":false,"label":"5V"}],"pinType":"wired"},"properties":[],"componentVersion":1},{"subtypeName":"Diode","category":["Basic"],"userDefined":false,"id":"5a48a43f-03ea-4bbd-9afd-312205a4efd6","subtypeDescription":"","subtypePic":"a7e3301e-fb46-458d-916f-a05c0bde95f4.png","pinInfo":{"pins":[{"uniquePinIdString":"0","startPositionMil":"14.54166,49.58333","endPositionMil":"29.08333,49.58333","isAnchorPin":true,"label":"cathode"},{"uniquePinIdString":"1","startPositionMil":"385.90267,49.58333","endPositionMil":"400.44434,49.58333","isAnchorPin":false,"label":"anode"}],"numDisplayCols":"4.14986","numDisplayRows":"1.00000","pinType":"movable"},"iconPic":"4bf63cb1-3675-4452-8ab6-1403298522d5.png","properties":[{"type":"string","name":"mpn","value":"1N4001-TP","unit":"","showOnComp":false,"userVisible":false,"required":true},{"type":"string","name":"manufacturer","value":"MCC","unit":"","showOnComp":false,"userVisible":false,"required":true}],"componentVersion":1,"imageLocation":"local_cache"}]}PK
     B"BY               images/PK
     B"BYP��/ǽ  ǽ  /   images/0b351edc-7875-4477-b820-546ce15be531.png�PNG

   IHDR  u  v   ��:   sBIT|d�    IDATx���}tSwz/��$۲0���Mblc0fB��3���@��0�b�!d�qN�bν'�tAgڣ�rf��i��Ճ���M�8�Ms�z��� N�`L�~��-�/��ClE�e[/{k���Y+kY��O��g?���S��ҡ�D�P�C���{HDDDDD�;����_��{�R�=�p����V)v9""""��Ή�:�t(I�R�)xZ�Q��5�cR�GBנP�@��x�1�cR��+o6I���t�|�&�I ����W��ǙM~��<>/(�^h�J""""
O����=�p���`T��F��:ix./M�8�IV�0<<,�0������ ~�}�M�Kb�J�/^:���Q��)��ӣ ]��+���!�L-[�,(q��~cP�Qx��+u>HT�*�GT�K�N�F#�0�����BN�T���@{��c�NQ9*���!�S�=�p�n�DDDDD��abg�{�aR祄W��="""""�G('v�~I�v|b��
[�M�6ן)�B�;JX�&"""�^�N�dRDO�f੅�`�b���y��A�����DF=T*~��"�bb�������_��g}� �L|v;>��f�@�|y`��6��~�PN�JU�Pث�B�GIDDD^B1��^Jx�PI�g9������~�1��y��\oo/���@�Z����80w��Y���G'Q�f
���c��	��0����'�C
���䎈��h�P�:�aLv��0�Ə��8��/�ҡ:m�Ҡ ^��٨���w��cqyX˸�˸�Ըb����q7��
B�b�J��X���Z���qu\e����MRʕP��{`<�}���R�a��A�<�,]�q��G��s"�������m>=?*v�~I��v\���H�����_�W�J�@�g�DDDDA
]1���1!����(F~�r;"""���N���);`W�*���	F~�r���`�#"""

�r�f��0e�tk�f����봯��f �S&&�ݮC�RA�R1.�2.�W,6����O�P ֋�y�q7��I��f��b�`xx `�Za��  � ��������"��<x��:�����e�?�S `||f�FGGKllRSS��!�2.�2��q�b��1:j���H��R*��?���\�e\�<n8`RG����`�Zq���ޅ��?�6�������9Z-���/��#�uB�)�o�<`�P�B�|ǟ_W*�P��D h��q�?>�v�Wg�˸�˸���B��J�9s�tA*\����xu1ʸ�˸��L���������z��c;Vcn������ݻ���|���>�����ݻHNLD�R	����	L���X`������͎/&&�y��]�����BZf&������(�k�Z���?}(��"<����8f}��6��1���F�oV�[���pa�P(`���q�q%�+�@.H]/D�q7�qCYd���fý{���ڊ�`�Ղ�y�H���%&c�}p���� ��#QJE,���0������F���`Q����b����ܩ����)lF��� 7&����q�q7Xq������˸��	���&A[k+�:��א9/��x���`��8J qJ%�J$ƨ`�����������'�=�RRR�z���.�Z��ƕ6c�MPR8.�ZZZ�~�ʕ�D�0c\�e\ƕ�J����;ר�fɒ<Q.D�q72ӟ�|U��Ʉ/._��cu��j��Q����qc
̍�A�J��]��f5z�菡/-EFF�#�"v4�=W#�x�I�ꛦ@�`
�����&�)�e\�e\�X,V�_���~�q7��"��d��_��G���I0wv`��W�1
t11xT���}�O���B{{��1"�ݎ�oa0�K4������:��d�o��a�ڄ�9��&��$�� �T���x�_���＃��nIbE"��� �&�D����(�0��r###�M}=p���`W�A(M�*H���D�u4��?��ݻ��$""""�DLꢘ�f���1|�7��SWWP�����k���gQ6��t��W��!Q4aR��Z[��#;I�� 't�X�ɱ1�{���ٳA������(0��R###�ZW�m"�;�2�r:j��qq���Z���m� !�r�a2�MY"��������(����B�sc����e��F��vxW~�kV눈���|��.
Y,�7��|�C==r�c�����~�vÜV(V��ЫE&uQ���Z�#���N��,N�D�݆�S��J�
�J���@DDD�b�@4��ݥؖ�,�Y��5O�C��`���54`�ܹ�Z���
�����s����{H�'��9?>T��A'Ʊ��ӽ~nll�!�q�qe������u			�˸�BqC�� �L����z����_H�X,�tu ���m0�X��!t~�%��^QJn
@7��C�^�N� @�MY!�q��Ұx�b�~gxxV��7H�q�qŌ+�����;V���Ì˸�+s�P��Q���/��T���/�P<�Q*�Q����,�PB��.N"%��@������D�/!!j��q�q7hqŒ��������{j�:�J�2.�7T1��2��혫���phn���cm]��~'�PB�B�����=��WU(��K/��^�1.�2.����Q����˸�x�P��Qftp�PȾ��LT
��^ht�Uj��h����^:��P(���u�J����.�			���^Mkf\�e\��5�X
E��!)�f*)�2.�70��2C�3�'�J���.���(xZεu��!�*]LLFGG���+�x�v;�2.�2�$qŢT*#���q�\1��211*����ƬT
�G��P���P��/^n
fܹ�*W /r�͆��Q��ĸ�˸���v�,�g\�e���5uDaJ�b&�F�t()X1���P�Jc�����E�ؘ�(�*Y��B��J���nΏ�ؔ�6G!""""q1�#
sBb7�Ǉ$��oʙ����(ېh��j4rcF���,��B�@A�Mِ��������])�x�P�æ(~�����w2�����:�<�������a1.�2.�J�A�<|�rیω���q7��"^9{)��C%1P�	��K��?��Ǽn����+z�իG��~��|y��	Q�-���	Ld/Ď��I����%9n����Ʉ�f~��@���ʡ
�BiP EQD3���,�+uQF����/>Gl|<F����G�v;�͐{aK���1P�Ѿ��'v،C�Û/x���ĩT�
����Qx`Re2�z|u�#h�ڐL���vL���Z�B=�O+�|Z�w쯼��ݎ(lm6�\����

{�(Q(P L�%"""����.�:�ڝ^<��>�R?O��&��		S�#Y����;�?P�v;,6;�=���P�i�Oʩݑ�8N��Z�>��  �ͷq����#"""�hƤ.����M��ۛ^=�؎՘+�ǳ`u�?�-�B�Z7f�#5�		r�h���4��� �Ä �m\���.�2��,��`�Z�����Iu46m�5�������CDD���A�{�i�3����*�P܌���۠��?�{(DS�4jԾ��-��.@��2��I5�v�PV���t�ㅙ�0���/+�'""���J]R'$ ��߃��fHU�6�s�h�j��B4E�~1����� ��q ���#;E���AY�竺=ې�Q��ݏQw���gBbW�gJ�����$�()�%i�����ꛤQ���#�����U4��`	�����I]�Z�y3>�������H�6F�6<U�W�y����6��Q�� P�w�3�[�� �a�ԕ�03�oECKǔ�7u����h����X��3Wd%��$�U��P���V�0[��kB��IΧ$�Ez$͉��B3�zM0�;Ө��ك�O���G�؁�Y}�rпk9�:6?�f4�t�� �9% Z:`�o�}��1���P����(�#'U��7�a8�i�n(5T� �T������R�π�]����Iա��է/OIn�vJ���Caf:*��(�L��A��I]�R'$������e$��b�����2a��j�!q�rV�$�؍ӈ��t�Q�|��4�q��}�^??ntK��J[`�1��[U;a�o��TI�03M�=��.�"�@W�F� �]��8V,q\��t�$/��b�����9�Iա�j�󮼐 U�_���-h�Daf:��lsܬ��.I�FyAJ�fKrq�� ��B3J�`ܽ	m�&�w�|��+�B�!$��bT�_����]��$�%yYh�ډE;O�d���1�p�ؚ<��_��B�]Q���B���)�����s~�m�&g���HҨQ��.˿CR�(ңzG)�zMh���o���AR%�rbR����p��e��Q��`�b�� ,6�J��/�"�����'��^�Ռ��x�I|��Ը��� ��+nt�>���:���˜�i��P�w����[��:��iҜx���L�<�ԫ��:	��s�*]����b�P߈���h�쁡����0�����fA����8Ū�+U�IS���ls\ؾ��(q�V���0l~ʭr"er'�o%�G0`�¸{�:{�>��ӗ/m~J��M8\+w�k~�><-J�$�U�W�����g����U��r$�6!�5�7:���F��)��5l~����`��*�^�S��*�����2�Z���|�#�%��(�����?�	]����ڂ�ؙ'&`��P��͎�+����^%vb��&�3�s����Gб�ȹ��5����h=�t�^��4���gO�	�J��=DI^�ǋ�����VSg���\����k�����f���:{P��%JL)�XP��Ǩh�pT�&�-h��ASg���sRu��v�y��1����vK��-I�vN��:��B3�o�qU�v�#BE�����b)��r;?��\q|��r{�����Ϸ���oEݞm0��$i����9��k
ڍ:�����^�O��o-��(�NH��?z	��7�@F��:����Yl6Xl6<��z}PbF#�+�l��TqgJ�H��wocw�_���6�fck*��=f��4���#p�J'֜T�E}��V���rR�n���z��
����sKĎ+�f/4;�r����V �zMn�[CKrR�S�����dm[E��9�q��b^��A��M0���V-��b��n������3��{1�}0[Q��ǎX{�IV}5�7b`Ă��U(������0[��TeMҨk7E�Ć&u�y�����������I_��yX���{�R��g���J��%vR����I��	�_b�K?F~َ��|���:bO���iHr�<����6���]mA��RwoBCK�V��X��<����C��R��e�����ݛд�nu�;J��ԕ�WjBr��Q�di�#����B3��ls�w���>V�_�;'ޙX�y�?0b�m�p�w0[a�Ќ�T�֯���j�5���0��PV�ܣS*7�a(+F�ي�3W��h)/�s~O�|�B\C� n�;oX	�_��I����Q	��N&�$�I�:*ۓ�/���(_����Hä� 8���j���~�0��+I�q��	&�
<��V�$$ub%���+�kb���5���Q/A�`�xu�t�l5ቶiH�;J���O�i��tęr���	�/��W����3WP^���-�><-�U��T �)�U�v$)��-q0�7��܀�*��.W-�u|�;���*li"�6�7����/4;�f��%VBYx��VT}x�ys	�d7w��\AҜx�t�����K�r�|��g�8���,�ñ�I���ZQ��<�B(܌��j'>����r \$�z�$�3��wl�j̍~�mƥ�%l-7��h���=Q�����0n�#&�Q���	�����{�3u%�=v�44#��[̔�(�FG���#K��ێ�1K��v/X���&i�h{mϔ��+�d��<%u{�9�	�֯Dݵ[nI�q�&$͉w�o�".�m���ׄ�w?F���:���H�`�-�3���>(���C��{��J�4'^�q�$'U7�1�	[P��3j��A����_�
	^�>/�r/l{!��TF,S���3.0��Y�~%��e=�� |�#4u��|6���,�+u�F���5�{��܌k�|Z�s���N�d�f�æV���ǲ?�C�Nn�>���1Y�&<�J��S\MW�4�����d`�"ZBmӐ�F0u{�9���0��n�6g�W9)Z�,�FI^�dӢB�1n����dO8Z:B�
�{������ӽ.�_�lǏ��P����*ؘԑGz=2~�:���q���	�qq�%%�n�atx��a�'<_H��혰�a�c:[|<����d�ȅ�{�T�gm�-���<�8����g�8�)��t��>ga�]�$_DDN����/����S��e�����`�b��4�S������9|s�"�{�C��F������v�Y,Ǹ��ݎ���1O��%6bޢEr�I�R����bb�������_��g}�߿/P+��C51Ԙ�΃�l���-�Y���ʊ�����$R�]7[�Nh�`Jw8��G�4$O�w0M6\�1���(Zp�exj�#���{cc�]|����LR������ہ�۝�u7O�뜺hQH�7�]˳�����s������ΰL�����q�g��{}&��[�M�x	ӳ�O��ݙ�����~��;�q=6�u]�S^���M������R�]7ݴ�$�ڹg��Y�S��q�X��|%U����g��d��w#�N�F~Fηv-f��'��z)��ԑ�ع2��$�Ŝ9j|��9ѹ�g��3l6qo8���0G��Wmw<�������fO��!n�(/ȃa�S���"6��tp�:�.@s�}��|+�!/?#�+� ���j/ݐ<f��'��z)���E����P�Th���x��=��B9?]U����F��U��u�~q��2�&���q��Ձ��w]!6/_��Wc߱��� q]ﾇ���b�'p���o�-y�q��E<��2<�jYT�'�ߋ�[ס��)��kr3 &�U�}]�3�P�w;��q3>��ɋ8x�d㐋R����j��s�O����R�".���_$�E%yYh���l�!eB8����$��q���|k'v�s��B�B��lE͹&�w� ���ηv:�h8O\���Z�G�6����gp���{�9g�'o:aL���:"�($T�=ڂ��J���|�ś�w�I|k���E�yM�7?#mJU�sּQ+I���ϭZ6��-���Lꈈ�����FU�WN��^�y�h�ϸ�$u{� ���,Gv�Źp�s�^
��q-�I4}/jvn��XVr�dSm���2}�պH��ʤ��H&����=�$�;0b	�F�MXrRuAm�ϸ���������}?**�b�êJ���-�[�,jΓh�^�۸��y���Bo�-z����A��8�uݴ�9��m�7��7T0�#�r�� !�}Ͼ�ix0<����q A��i2{�Ed\Wf�Ǥj��DW��+�����\�578��uT#��L���;�F��V-CG�P�.z��<����i��dRMì9ׄ-�\�.��A�h�V� &uDQ����T*��
T*�����װXş��so��I��TJ�`�"\��+H1�]����T	N �����T�����ͷe	y���,xU�h;O���z�v9���0+?8���2��ȩ��F�I]��Y>���Gg��y�wa�\uF]������סP��P�����4�Q��~�l�	���i��$g>z�� ��>���mbv�j�������Nː+n�JҨQ��9�:�TA�F��Mn�ih�@��Ge!�3��q��ͬ���nv�:�:(��z�D��n��d��|\����4�H�v)`RDm�Ch���;��G֜�ٟH>��l�|g@�a����<����<���;���6H Q    IDAT,$͉��}2I����-�v�LҨQ�g�c��ӗ�~f�oD[� rR�Ά*rOդ�s�l6/_��Ϡ��e5�=$����{hl������k{���W�'�v�8y���?�_ock��鏮-��w���Ps�	�cZ��#�:""��`ܽɹI���R��}Թ��� ��O!'U'�vEz����	����J�f�di6�:����N���e�;�1��j>B�>����?(y�h;O�����|4�~t���h����D��:""S��0[QQ�w$y~����(ң��G��K�f��f��0n���t���)z��F�EU$�on�4�h;O���F���PŤ��H���>}�Y6��۳%yY�>sE�΅I���n�lE��+n���"I�F�F͆)�N�bתe0����|#���������o��cDD<L�\\\�^4	�%8���&$Jm.SO�d�03]�ꜧ1L69��9&t��N�:[|?���X�F�,����jl""
&u!*F��J5}�>�(�ʐH�
EP^/Q��>}Y��j*���>�$/K�M�#���N$��ߢ��-ؼ|1��fmz����i��1Q�aR���P��������oJg6��9o|�	��A$�6��@ݵ[�*]��������T�_��<T�����&׺�a��ŲĖ�)ɇI]����\�+}��K]}���F��0�o�Z�aE��^�O_���%yY0^hv&�9)ZG�ˇ���y3�=���  K��L��A�(�tDD�I]���i�_���AsHT���j�JT�_9�c��FѧdV�����AT�a(+v�Y[�	��Fne �5���JN��An� ��\���D�]�����:"� 0[=�U�����-��ڂ�T�s���^��Id��f%��?�ڿ���IQDbRGD$���#^=/'U��i;ö����k�4F��i�(�]�����O��HCVr"���s]E�.���řIQ*/�C��%�f%\���3�  �]�"�u/l�MD��03Ezf�;g�q�zM����K��E��<wo���-0�7�M�2�ބ��[R}��w�֯DE�9��o�s�ٱF��n���S��L&��i{m��}�\5u�x]� 
G����d.'U��^���p�]�Q��w�àe{�9���^���Y{�#��uO@�Q56E'9���"=�w�:f��N9~I^e�(/ȋ��I&u��̕)�f�ø{��lC�ύS�����^�=�۳9)ZN|���P��U;QR}d�4.o�9��۟�^ۃ�^SD~�&�Z���qpL�du.���V�;�	n}�6���֮�%u}����)YbQ��+��(�;�a�a+���,��ن��+#�bǤ.J4u����T�(u|��8�K�P����O�]l
���v::�M��}�$/�Q�+�C�F�'͉w��Ä.��^���K7�.6E9��$�������M�=H�p�Pä.��8Od��<M�l��Aҟ����#�"I5��ls�l9}u�n9+ܳMY&""
Ur%Wf+�Vf��xS4I�v4 ���L�HN� ���p��Q�++FN�M�=0^hs�DQ������>IDDaN���x�U�W"'E����M�f^����K�ύ4L�DyA*����������﹖��VT��1eŨ(� �w����-�>}��<��M��.f딵tD�"��FE��y��Q
CY1�Qؓ+�2�7b`����Փ��-0��4"�8`R��֯D���S��D��QJSg��>�$�U����Q;�U�Q���)���g��0^hFaf:J�]e�VʊQw���QX�3��>s�g� 'U��usĂ�Ξo�"i���1��@��/sRu0�ބ$�zʖ�0[�1�><�ܾ�zG);V�������H�Ҡ�H���+��ك�w?���DD6�M����t�������$��?���+80��p���?,Gݞm+iު۳����LV���l��w?"ѳ�O��ݙυ{��ۯ�7w7Hꮶ��j��
^^����t&uDDv�K�b]3&i�0��03U��x̊"��Y$΂aR烵smXk��ܤ���VǨ#�N[�ɱ��mU�n�;۰{��!̝fBRRt��Q᫶;~�����f�˸20[�w:���7��]1f�U��B�_V�m�%$|Ez4�t����y��I��~�j��Z�q�Q�R���������!��KN��U�(EN����MҨ���P��Q��N����*F���>���	���䬘U���hܷ��ݛ`��r$q�W:�Y�E"&u^���~�slԺD�q����Ά&��#���%�F���Z���	8���T��圮�%��2s�����7w{�S(����|#w�L��4�;�W�zM(�(Z:D�j��yA�T�(��Qw�I���''P�~<ܲ�[�N	d��: """
?rW�\��������C��l&uDDDDDDޒ�b�:�L�V�(u&���� �oq���*fR��Q���h��A�ύ0^hƀي�w?v.Aj�ډ�"�dc�+uDQ���Hиw|�^���C�0.�$�3a C}�ǥ?���)��;J1`�F�>u��E��{C�J9���:(X�	s������&G�l�lE��Gg�� L��ԭ�X�#�R�{�`��ݮ��9K-D�o;��H���df+�O_�r�iܽ	%K��4+/�CE�%yY��ꮶ����.Ԯ�_�~�[�jO\�XW�(����(�c��U;a�oDCK�v:��=����F4u��j�JT���������nݼ���
�I����ԡ;'U���?���᪢H��<Y����b&��+��BҜx��MҨ��Q�/�0�#�R�rL�;U���h���PyA��BN�n�}d�d�P��h��m��9m#����^���i��䡩�Ǒ$�T�0�����6>O���7��{
�M�=HҨQ򰃢�di6�V��e�%u���h�5����L��MN��W,���q�¾�Ez��&��\���i�#T�f��૜T��>��(���sw��E��K��/����dUw�����H�r%(�LwV�\-�B���U���0-�P��hn�R��P��&A4��9�:�䡡�f���"�����)�7&'����4կ� o��#�g����-��܎���&7s�sv=��1�����%i��
�l���&W�;J���s��p͞��>���
�4�H�ހ�:""""��]mA�槜2O*��h�왶�2y/Z	chh�pTU&W�Z��2�q�a���,�v&�B�Vw�e��?�ꐓ�CÉOݎ��ҁ�<f�;�ϭ>s�y��wor����Kv��{�C (�<�j[�p�\�[ ϯz��O��b��Z'���t�i�m�&��ن�=�7$�OnL�"Шz4#�݇e"&V���sS��>�jb,�q������3c��$/u�nI:�
&L��vE�Y��Φ�H��؅����4n��U�
3��p��m�eCKJ�]�Uw��m
f��%�W�������2%U�|1��q8x�"���]O.��Gq��.��e�}��g�CG�Z��x>Ea�\[ߠ�1�.�L���+&uD��e�x��$���ĳ�p;� ��w^�,���EX���Ci�j\""�ʹ�+�C�^O����zf�_�ufBu��f;�֯DyA^@S���{la_�~%�֯t{��j�]�Ȧ�geM�
UɆ�gϵ7YCK��rVq��®���Qs�	 P{�j/����L�]W���;�]���'��|�Y�Z�b�W	��B�䛁W���	���(b}���˪N���A��;/��  ���������5.���K|��t�,y��r6Ez���9s�ʖ7rRuHҨ=&��L��Օ�e�-E����}����n��L7ƺ�-0l~
���0[��2��j��
�d�[;q�uj���}'�㍀`��}m��<�s��E2&uDL�krB����`$vL�HJ9)Zgh�!L1�JI^rRu�H�Mi,�4'~��,ꮶ�03I��4N�6�9���칾�%���.���S �����E8���:��ΔXI��1�#")��9�|�0M�x�ٱmA�S!gC[�	�~����f��$5m������kKա���?{��s����j�w�pt��$����*iN���n�ȑ�y����1a��H�����r !!a,!!!V��^zD?2fW���#���?|D�1�;����7��N�fK褊�Mb%EbǄ���TQ�G���0^h������C}#��7�:3�9m1'U��Ι��~_LO׈E��:��K@M;����w���vT��������E�>e�	d���������P(Rl6[�7�x�b���h4���[
 q
;  �_(�a�4h4J ��Ð���x��i�YG:Ψz�\V����N���n闟�������ݛ���g�J��B�W	S��+h�t44��9���2eSs_�����U.��l��p�d��:]zJRZ:`(+�j�_ݵ[���t
3�e�|���G�
�X[z�+�O���6��^�����INN����Wm�
7�Lꈈ�䒤Q��/+P��Ѩ���E��N�JK�3���,��r%"""��!l�0ymI��������������I:Ez��):peE��{
�f&tQ��:"""""�0�JQ��N�";Y+�0�����z�=�"l�s&uDDQ,?#�{�C'�P�������>�j>���.f��#J�|�0Fu:�l�)���f��A�j_������>cn]��#���hX�#�pm��A[�i����T�sASg�c�Ym�+��(/�s�Z����f��n���z0`����e��'i�0��mJ[w��������&��z�8+uDDU���c߱�rCTLꈢ��x5�t���/��S���0��03�~�|�𸡾�ou>nܽ	�ݛP�QO�e�o��
��Iա��� ��=� 8:�5u� 'U��M��a9J��` ��F�������Z��#"���5uD�rRu��Q���� ��\AҜxT�_��k�����U0^h���U��1�2�Q�~�W퓫�\AyA��P��i��03U�FSg ���C}#��l��A��7���A��ADDD~bRGe�֯D�F��ӗ=�|��I5�4j�z^�Zx��>�o�5�03��騻ڂ$����:�4'ާcE#&uDQ�$/f+Z:<�|�l������-(��Bݞmh��P�,'U���Y��03 �������LꈢLҜx�X|���<����F)��b���&)3%h���z�I��xEz������IDDD��Ѭ�VG�w?vLߜ��Y�~�Ǧ(��bʊ����T�3�ބ�Tݔ�~DDDD��:�(30b	h�����Q^��槜�T\;UΖ�yb(+FyA�����?"""�h'߮�D$��k���Q��77YyA�s����+1�7?r�ss;��/4;��4;�qwoB����x�c�}��hfLꈢL���0[QU����'o.4T)/���|��I��v��S�����?@��l�TaBGDDD�#N�$�2f+�><���{�6��SeŨZ�-Ω�M�=�>sŹ����9Ͳj�JT���EN�ι�x��G9咢Nv���Zd�$�m �67�c�\�e2[q��>���k_A�F���4�g̃N����A|��=9��u��:�(Tw�%�&GW���xSg��'��h�5�� m��q>����H��RYQ�G�F�8��8\�Y���~�(�g��L�ks3�� ����_��`ڟ5�v�\k'�o�z�=��*�F�|���f"+9q��)���i�2��8w��[�"�=��������BZF���'��t�,š�Өa��#��_]����4Ծ�Yɉhl�¾cgq��ޔ�w��d�bד˰c������w���[��6>o�k¾cg �6���uO  j/}�|�u���~��'/N;v�F��[��U���?�'/8��؂����®w��z�=d�hQ��)�O�Z�)X��~#b�J��V�|���������O�?��R�@���_��ɏ��DRQ��Ԕ(��3r !!�k�N�P���~�t7�r�(�}�5j�,r{lB��X�bUP)��o�u|jK+���bhb|O[>~���H��u�(��Κ��k�2���V�w�ηvJCj��\�-�\l^�X��w������5Ed�L���[׹%X�V-Á��ܞ����q����P�q�����p�'/�%э�](�����E�s���7p��E\��
�c<y��oLy|�����}�+�q{|��  ��������_!?c�Ǳ��c���n�����7��s��9��"��o���-n�TG���δ�����
���a��_���]n1�q�o~�L<;�����Y�7G��e���/)f��X�#""�'����p{,sI.�sf��x-!6�w����o&�P�%�ZŐ�6>ϭZ6�z�t5*�b�'$KxYɉxqm!^\[����8|x���ӨQ�s��=��������Q:n�L>W�s`Mn��&;y�X�1m�|k��Ǘdz��c ���X� ��؅�ɳ�G�5��Sn���k���@JB<�-��X,w^*�O��ޫ(Ê�#��>&uDD��AF|U� ������^��B��~��I�t��q��8��i���9�$�8f�d�}�<~v�o,
�ؕ0��d�����p������xs딤�d��d�N���*�k�s���8�ډA˨������?5q9���qJ�[���}�㞎8�E��V�c��}oʴda<��p�鷍�]n�����Z&�6�}J��쭎)cl�?�-��)�g'k����޹�N�tR")��lْ�P(*�@\\�)>>>I����}� �-�r�HU�W�_��?�el���}�G�M�&���%A�Pa|�
�Ō����A��>� �`��c�{�F�W���f�~�v<S����Á:F�?xl!��q�����_�!p$��/�������O��{�!��dMn&�� u�
:���B�~��wܞ�x���"I�ƪ��`�2��?:�������7���Y�����͆�w7���|k6<��F���.�?E��.}������څ�N�gh���X�$�[����;�L����:ׄ�'/:�ҝ�:}׻ﻍ���˨�|�ۿ�8�K���;�S����|�|kηv��>��-:�����_��?���������9�������}/t=C#h�@Y�b(
��@�q���.����Y�P(�34�m_�F�5�*�����q��&H)Z���t�����?����#.��Q��:�dU�W�PV��fﮞH�\gw{,1)���n�����I�Z@��a^�b�'L��;_��2�r�G��	SߤZ&���F�S�5w��HC���g̓%�7��%����۸zʚ2!i���63!�6g����MY;(�ף��5uDDRF'�KY�R��Xb����p��-$ν���ˠP�_��K~F��n�m��/6/_��?y�GN����D$�.��Wv��MGX��ӨQ{�\��ų���n��4�pg2[�$k�SovonŮ'���U� ޻�?+7'""�R�e#!1s��	 �զaђ����t\�R1���8�Ņ~b#�]O.ùW���N����{e�ٹa�'� ;E���
��N �G'u^�Cv���݀��Dh�����B���x�e��[皘 ������>���.��5���m�s���L�$
+uDD䗌��ߊo:�����FO����ڧ���V-s�W�dS����n�͋k����uʪ��[��(��ȹ���}�κ}>�nj��]�ۏPhb�����6���`6[1<t�c#r'(�=��3���O^�8],P�k�^EY�&t�����r��v�R��HCv��c2y<D����<u����'��X�#"��d-�.���u�:t����=$�H��]���e�}��kr8��J񼷗?��q�߻e�?�uk��!�{d2[q�ս5���,L�B�-�    IDAT�Q#?c�3�DM���P_�]Ҫ�������{���P޿|��9�2��^���������?CaSw6�!10�#""�`||f`�L`��M����3f(�\[(j�r���o��ý������5��آ_�2�d�J��N�.�׻��K7P����_�b�G��y�ٹ��9�f�k�2�=՞[�Ǜo#��oI��Wy�*�����\���Jvq�ܺ��s"0�#""�%$$  t:Gu�61�ί?C�|xL�l���mA����8 B���A�^���.}�S�⪣�_���/߀6>{�=�]��T�4��iԨ��.�vR�G��|{������qp�:Iײy�0�g��N�$���4����I�F������jo¼�Q�5)��a���m `��)F�)ڀ�E����ɋ�iWb����ɋ8x�"^\[��W�=�0�Į�bK�	����[��ֹ&<�j�o\�wr���B�k�,�:�b���'l*��1k'u�l���}�7<������{���%v\cG�bRGDDS(Uq��O��wU1j<�Y�{�����;�Q١��nj������lE͹&<yQ�QM�hm����k�:�?�]��nS}e2[q��E�6�Ry��c*��uO���B��X��=�6(�i�صj��sq�������w�\��qn]���f߱����t�cp$%�T,'�^{��hS�3�ܶ��vL3Y�����
g�B\�o��A�(j/}���8���#�pp�:d%'���7�wg?þ���{�*|��%""�hS�C��sal\<2�W  ���a}��v&�h�e��B��������~O!�Ǡe������V�<�����6>5;7x�$Ц(�ͭ�<r
��Q���+��y���[|�lj��pp�:���ܺ���.���oL����in窘�b���~}&�^1�x�mQ*�:�:��	�����	{���O^D͹&����7�:߇5��h|e��gϯzܯs���4 "� ��b�͏<�W����q�����ohԌ���qv��C��6%���KG�Qc�������K7������йjl�7j���Ϙ�ڊ-3>'��1B��yc}P:W��]���;~U�6/��)�a$l�1�����E�L*���+�� �۸�����"d�:��zq�I����J��0��Q���z��;��>�l������ߙ�L��G��;�T�o\�״�}��e*�l-��R�+~vv=�{� t��4�mד��n��7�]��hvٚ@.��Q���{}�?�u�(��k��Jr�E��W����bo��Ϙ�׺T]|�$�������3WP}�J���f��ɉ��I]��N��E?֥U9%z��@������ZC�1�c���~��z�=��(�!�;��.���f%'bד�^����'8���?G���x�m�+�bp������o8��:�2;E�5�����=V��Y�z�\�۱�����:""�Iv�q���ҍ�K�B����Pvx׻�!?#�{��U�ńN0h�.�q�Wn�ij���E~'ukr3�������T��P�,����uX�F�,�����޴9��m�;vv�ϡ�o�}�f&kr3Q�s��ݞ�˺T���nKͯ�&wLf+�:�aMnfT�8��#""�d�'|z���N�� �7>x�_	�p�*l�i	����>�إ4+9ѯ�ukr3q���۸�6��?���z�x5Á>c��]Z�Ө�ݢd�����^�[;��Z�S���߇�(�[;q��E�X�����v�|�_�ŵuaH��F9�2�#""r���e>%.Bӏp���S~��g�õ���k/:���[ס�r�����1<����)����^qͤi{��8����f�9���Em[�y�~����_7=Lf+�j>�ؽ����)Z�)���8���[o�|��H�����c���ɋ�u��G�SA[�c2[E�н�p{	O����q:�&蛗/�����]+�pv��gn����I���ǣ�S�����y�K��S�6Q	Or$vLꈈ��i�3n<<Y{�`Ht��Še�GNy����f��e�C>_���?g ��������>�o�t�pt��k��E��!f�)����yڭ'&��c���V-�Zw��ޔ��q:��<���1�#""zhMn�O��bP���%�2���ِض�N^����VwMf+�s��yc=�7�c���'١�Se���uAٻ�S�x������K7<V�}�Z[V��������N�&�n��`&vLꈈ�Z����}�!���'>���)�P�ꍎ�!���r3`ד���k{���#ܺ.��� BE�}����D��)��L�;e-ݠeT�
��)� ����{��&�O^Ĺ[�x~�㨯��J&I#X��:""��|�8��<�����s&�}����{>�/��8���4j�=鲒��F}s+NL�����P�N��n��7��^!��p3#+9ѧ�)e�\غιf�����7�!q#�cRGDD��/�߻�#	�}�>�qJ���n�''>�������OIK�6¨<2�<�n�1x�as\�u�&�����Og����2��Rh�:����DDD�|�=���A�׋��n�&����Lh����۞�^���֮���7�M~F��]=Ϸvz=�-;y�J���Nt��mV}��-"��lŁ��.�/���XG�醍��Wx�xs�xޜO7�K��{��a���*�>6�:"""������rm��E���7����h����ـ*%�u��V��͹W���g����+Q8���uR�671��]���﯆.^�s7��V5皰E��b�*������ۢ�5�tS��H��4��S����8�p��/o�k
�6$$=�;N�$""��)Oӹ�g�N���ߓ�/��r���ـ�]J���{l).�u5�u����Vv6�c��+)�����K٠��/�}+��@V�܈M��)�e(�I1�I|����w���x�N�ӹ����M#�2}.�W>�}W���u�����"B{���je0�����J]�ߚ���sq��]���lG�{Q�&2$�;&uDDD>2Y"sO����~U0"uj�/�G�ur�ٻ������y�X����5�b�]�I��k=}�&o�0��[�9G'i�����:"""r�Te����Q��Gܧac�P6�&�/�y)����1�#"""')׶E�Ó��5�vEl��W׻��I�X{�I�EJ���N�׏"���:"""��s��\�ʛ���ͭX�s#�����BY�GAY�8p�":�ݛ��1��S%y�[����]��8��m4�v���7�T2)���qK"""�g���������� �"l��c�_��&7��/��0�{����u�ZG�д��}o�Y''�J~F��s�Ө�����-&3���<r
�+�q>&��uR���[�0Y��o���F�] �0�#""�o��z��Г��V����Zq��zr�߿_�s���������4j|�ڞ���_�z�����WQ��󾍫a2[�*a����N���66/_�|,н���F�씩7|i��Өq�'/8�4��������E	;N�$""�o�n"m��6>5�6�M�Qc������ƛ�F�^_��y�`&;yj��E����|�V9�vs н��F)v�.X�a��/۠T�-t떩Ϙ�]����B�ǟ��Lꈈ� �6���H�Ey(�ٹA��ʵ�(�db�2��ٟ���^T�<%��C�r+'�ي}�>q{,н�<M���ٻ���;��H���e!"8�Xp�d0�f�T�2"����=A�dfrj5�����`������cMrƐ��(g-r	V0Nl.��E�`ld���ڒ��R_��;�����[?���r�~��<�H����<�'Q�wK�_P!ъ6��  �"�bf�y�g������+�,��mј�#X+y������ӽ:`Ц��X�t��e,�^D���'��x��We4��Eya���F�;9c���P�/��h�� �+����;k�~�"��Ƶz���*��灻�g*<r��:?ҭ	��P�7��;^xY�O�;��������|v��dT��<sf<{�S,����7|�p�$;�����=�Ԗh��Ǵ��c������"v�:  �8�L3O5�)+�k��BvݺV�xP^F�v�yh������*~�a=s�����zC>�Gό*���3򔌑:i*ܼ��3�źw�ۧυ����|5��=q����w�=֕�ЁǶ�ÿo�-�Wh��"
v�:  ����}�����0Wm���Ѝ��<pg�ih�Z��f�7��ĝ_��o�ᕤ'f��3 X�蝹f+/#ݐѺ���z��>l����9k=Z�{ׅWO���
��.p"M}mF3���c�C�?��zC����p�`G� ���'��ւ���I^F�<�=��N��h��%���myံ��i�?[^8`�3�����Ϳ�k̺�x��4'�>�A�g�q�'"�jj��oה��4�y��9}oe͠ue+�Nen�<�(�����k�`G� `�h@�����*��{]o���L�ڞ0&�u:���sa�9=m�C�Dx{�F�9����!��}�v����F�֕��3�6�,�軤����/��3��̙��W<#b���ٜ�	=3�0N$fO5�kK�|��P �4m�����i�� /}垘*]:��ㅗc�s]�
Â]����Q.	�f����HK���~L���-}�7�nH���_?6�㼌th�mT6���j�H��_?�����;��>o\S�[W�b�F��=�ˣQk���hb��hԡ�C�`G� `��_?���n]kȺ�D��;j�+��x��ԉ�K��r0����6W��z^�륦k�<=�n��~����������״��A��������"��W��{oW�_�3���N��hǈ�3gf��ٵ�`��޸Vo?�+������S���#�{�o��b!�5Uj��%=���k���*������I��
��l۷o��X,�jPzz�HFFFA�������1����n 9�ׯGn�|T?`�}ӵ:;�S�a1xx�Z5��ӵO���P�ק�O�j�>'���}�����7]�W?�X�/��$JMY�~��;��f�꺽o��_��l���u�Z=��u��Ks�tq����>�=��>�{n�TinV��nS}M������ڕ�.-TEQ��33��ժ���#�~^�޻I����-U�s>�=C���r0��ݖ����{'㪜�=�ԵEya���F�/�^V��3�uin�vݺV�k��۔�f׈�#�קue+t뵫����ڻs���s׆�{��ׯ/���G�W[�����>���<U�j׭kuནQ��a��H��?��:���Gkt�z �L<��Q����c�o�lІ�Fx�+��<B���:0k�ቾKz�翉�o�?���~�E~k�Jb��tOD5N~��g�[�f��Q��Wն�Ks���e������z=��=�]�.������R}MUܣ�������k�J�|T:��U��ը�jK��Q�o�>�/,WF�~	 @8�=��}ݳ(�h��H�+�9�;�z��Ԟ�V�+[���_ZU�btRl�fk��̜j�oP#좩�:�ξ~տ�ꢙh�4Li��x����%�k��:�I
{~���|X��a�%�<�_�Չ�~}m���Hm��REa��>����5e%:��v�}ӵ1]����O��;�j2����nԺ���gS�Go\���ᾘ]g_����1�~����L��ghT�>���rm��ڶQEyq<�קW;>�ۧ{U��PuiaT���������z��.�^��FO�:uqHwT�Ϩ����麇����;��y�1W���?����~,��-U����Θ2��{'����bj�/˾}��V�T5 ;;�l~~~l�u�<��N�R� &�̽���*SS�JjY�x�+MM����bL�,9#.����[I������g�rS�{�9�	�j��%m�6���;�~���Ж�r�++�-�W���y���:���^C�_EQ�*
��N�]ZS8�SQ��'�U}M՜"1�t����̙��-U�:��v�e�����W���[,��0B�<B�x��a;Z�=��_?jHI��l�Z�}_�'�}�b	,�M�g�ߊV��SϿ~,��Έ>z��o��C|$����3>v�'T���'�YXغ�Z��dF(
��x�xlFp�պ���|?�B)  \Ů��z��]��>������h��I�t�C�����z����W�-���
sD��(O��G��{�^:ܡ��ް�N��V��{o���^~�d�]8��> S�e�1��oI��� A��a�c����k�D�%�u�����1��U����J�7_רS�S
������v��ۧ�E=ʹ�0�J���1������^��{5��,d׭kC���	}󧇴��
U�{ȩg~�֢�����+[��L�N�]ҁ��3F�������P�%�P\�#�tך?�������望�R�����ŢQϤʬ�����������d��D�����=8��!��]�᪢0O��)?ӡue%q�6�f���L��<pgB�v:������#ij{�[V�PEa��T�6$��R�>V�uh'�.i�C��X����5}���=���?���z��	�0�/$��;!��`���4����nB��Z���2?}l�IW_��5.�<�H�J�sT�]���옟c�Xd�X�i��б��9���co{2�軤��^5<�m�*��pF�����vEy�(��at"%3�IS�58�rv�x�u"u*��f/��H����v�?��g��7�r��ict��H֬r���d�Ŀ����gҫ4�'�j�ߍ����?�G��0��A��x=��H�O�����jo|(�s;�]T]�+j}�A�U�QS�5���
2jo|HY�k~E]����}���˞�#) �,�H�W�#�u~�1�R%Q�.�^��v��FB���W�����bڠ|1y���)A��SL��(O��{�*
��o��>�k�����:�w)l��p�G5��U�r�������{����g���{���W,�=c���@@���# O�P��b�U@u��'�-�: 0������oPS�fu����S=3^o����,�W�Oތ9Ѕ��9tV�.�QFf��)�)�[|ۦՋI0�xl�)<���pGB�q�ݓ:��o�>2r;�X=���{Be���[j���Pn�Z��¼�7�Gb�^���7���?c�����ڦIϰ���~`O�UzF�����R�q���X���5�c��O���O�z�Ԝ��7�q��?���"�=[�O;�W���u�����KW���-�/<��EO�-ȵ�,�@�EJȲ3B �Hǹ�*���f~��Ӱ�35J�s���7�����k�[7��z��O���h�!m�Xm��3%I%�*��9tV}���▘��L\Y�d:�wI[^80���b��ׯݯ���}��}4{m�b�!���t�����Ӫ��im�*׉�KZW�bN@���\{tL�n]Z���]j�y����e�k�w�~߫�փ���K��&<����I��ǆ���#�4��{2d:����g���뫵c}�Z�ר�'o��~��j�'�%C ���,����j������%5�>���b�6�u `2-G;UW�F;�W�y�65��MՖ���~��F����yNN���^5�xኛ�;ߩ�K��h�u�<ˬ���w�Q���3��YО׏�dDg��Ѯ�U_S�=ܹ�G�9%5o_�������ۣ=ܩ�����-e+B����:�}�o����GN�jW��9Ӳ��{�Zo�
�W����5��jxxX��.�ᰫxE���	oC0�u���h�%�[7�q�F5l���x�`�t�����n'�k9 ������l��F_x�EO�mͳ[�,ғF�S"��)�\æ�?���͡���fW|�Z]�=���ߑ=-]EJw��n��bY>�)����ۧ{��;ݨ�����K��gm�����s�}G�����j=b������E0:���A�^~�d���=��yL��~x�ywG���،-&��	�{n�F\�P��ٕ�?|����Ј�3c����B�XW�B������p�{|�����*=q% �t�#������d�    IDATu�Z=���q{��/��F����v�QU>���!g�k>?ӡ�wԆ��{��A�=����O]��������Lӛ�Vk�Ƶ:r�wƿ/����S�?]o���3U�����\Ymv�9/�\��UPP���jY,���,;�W��zMh}�l͇ޟ�~�?�Pæ��3[��T�Ԛ����>�:��.�)c�V_|j�)5�|co�U��w�&��	�<jz�jy�>�>����o����%��b���Z��z䛼�1���̑�jU 0w���D�%��{U�n]�g�ݔ���>:������,#.���~L�wLMI��Ji�s�'��[�jM��W��Kou��;qy�tO��G�{B�5��XÕ����w�N��N�vb������{u�T��U�umQ��T�Y����_dL/��j�F\�}t&��	�軤k��gs�jm��SI�s���ܢue+f��RU�-/P���Ϩ$���\�ۯ�wԆ�o����ޫV+?ӡ]���V� �1����{�O�5��j{�Ka�W޲z�v��S-�`�
K箅��[������wy�Z���Ӧ���z���{~�8I�����ڱ�zN�kj;��G��23���w��uz�᫟��~�5�[{��~k{��.��� ��h=~*���k`DMmG�ކ��J]�N�I��^�vISB�=�_O����7̎��=���;�[�s�v�?���t���=�_{^?��~��?~C����]Љ�Kz����tʗ��`��/�����go71=��>o�u|��V�	��k�TQ�7��#��ծ0[\l�Z�-aF�wm\��53�`�e���0O�gmi����ue+tǬ���j]ي9[`��^�k>�aij�qKUy(�Mn�鰇�|^v������E8�7�5���]�=�Iψ�3.j�K�50r�"&�~"Ia��I
��;�ھ�B��������}��k������� ��*��UwcE����	M��e������}���'C0�m��ӄN�
�GZ�T���k�+o�|�e��#w��)Q/�Ow���=�I���1m����m�茜�ۇ��u8�����>����u|�J��3��{/���+����<a��=�Ԉ;�}f�]��.�uI���z��M�}��՞׏���j����[uy삡�-�t� ӡ��]�Ѱˣ����V�B`����eFH#�G2]���>�ᗿ!�{0� L��������Tæ�P��. ��Z��e~}�{R�%��ͻ&imX��>}nj-�+o���JwTMM�="���Q�軤{/��ӽ�v4.Z�~���#�u��aG�"�tO�����a�%�u�IZ��T������-/���u�	��[%L}���g��qy�ďߘq<�����;Bk�z�FC�ئ�������{d��C#d�}����ȭ��}8r�W�=���33�����I�軤�_?�-U塯���P��S��r�x�==��7B#fӧ�N�{�k�v�릿�g~�������N=�ũ_���/���J��^�k1���U$�?���)+w��3c�w*��ڎ��z��nP��݆O�����y�.Co��~�5�/�k�B �PS�fՖ������t��M5j�����%�~�?��m��Hekn��s�9��V��V�#[nט|^��F�~���p%�}��� ו���Iq��3�O��m�EX*�jN�]҉�K3ʾ�*�_���<:����S��{�vzi[�i�{�\hs�`_x���:τ=���^U��8�����K�;TQ�7�ks�+o��׏�9^��U�+[!I3B���9>��h��������R�=�{n��\)|�'�.����{|�s��~�O����zo�{ZJ�N��is���3���SZUPF����;��L���݄}���B�4��)���O��f셧Z�a��^S�����:B �L�7�]#�@��YW�&T9,�i9Z]�Qc�^��=!ɮ@�+�-���IҤU�u�O�ե�C������42�*#.Oد���wΝ����FL�;>�ߍh�'��.��ْ����K��>�Ν�@��(�`�q��ר��t��\Fp�ѷ���z�ڱ�Z�[7�ն�<���@��ŧ�O�m�X�����5u `"�������4�o�w=B2X,6��W���MZ��Z�y9r��]y�*i�my  fc��U~�t�����+��5֫��Sr|����l�E���;��`�Y	�׆G��x�Oޜ*f���@@?OŴ��F_x�%��)�: 0����?�@��Ȝ�d���Q��g�TKs�++�L9y�dO�Qzf�` H���1]g�ٵb�M��s]�kt�3y'���M\��i�[Ԗ����9�k�[7���!U�ݣ.�a�'��ymyiT�	�o��}�D{�/�$�nm��F6[pyp��|�E�b��]�:#�$t/�ͦ�K��
 �Q^����^���Y�Z]�^�44����S�P_��}v��gj}�����WN_'���������F��9uk�f�Z�-i~kTSu ��4��w���C�G�bY4��e�Q8s���>Y'G��d���2r�W^�_���r����'$���� �����ʟ��V����r��S�K���l�Z��R��oC��?Sæ�9A���)�~�ID�.gk��k����y�uF$���/6���>Ց��G�)�B� 蛿����v  ���Pqh��O�d���ҭ�Ϻ�d�ov�+���ۡ��٣���W��Ψ�y-��Nijf��A��'P���J���e���N�   ��o�98��')i�Y����T�a�@@B  @d�wnU�j9ک��|Ֆ�������8w1��A��P�  ,k�?yS��^h�W�7�*�P��Ў�Ւ����k��Eiܻ��_F;zH�  �Gp�dI���"�R� �l�:  "P����?}]���uu}���T燞o�nij�)x?D�����H]æ����Xܲ�Muf���uQ���f  ��L_s5}J��a�G]#j�߬���<�n �A�  ��~�g��f�~�G���
���T7�T�O��q�F�%*�Q�d�X�=$� p�奪-/���~Iu�kTY�0�`�z KK�*),���t�4  �*��r��O���Eu�����R5l�YpS\�K��g|<}ۂ��fǹ�Qm���P����������!� �G��5顏�'s4�cW��snN K9ʊ�A�F=�*��:q��y$��%Ip=]p���������M5j޹M�z��vD�;��F�Z��RÏ~1�܆M5��;�]T��筴���y�R�^k9�*�_W�F��?8����FT����q�5l�	�D�<j~�9�g���HS!)�`��H�9�ػc쟟jMu[$��6D}M� 0��֤���B[s��W�y��*�,����Ue��(-;��X,Y,}�y4t�du��e���r;�WOU�tyB��Z?�DM��U����d:���}3�Nנ3���6��-/Uˣ��dD����T�,�t��~��n����v��ᦢ6n�0��'o2�`Q���E�����: �~߄��㲧�H
�/�2����5��f��$I�w�*v���T���h���Kp���G���G���Q������7�	{�VY����|��TS��<�,�W��m��^z��p;=��<jj;���ҩ X�F�;��� ��X,z����JϋOu���O�m�(����R  ���:����х�?�u��ώԨě�uA뇟�x-P")���v$t~pM^A�C��6J�褩i�;~�3u$Zjp��� ����BO�ӧ[����f�ێs��?M�l��ϓ�  &��%�xro��bm��RB �X{�C����io|hΈMp�g�f�M��n��?}=��*�M���;rUZ�N�׮Sz����a���N��|m��=�(S��S��s��pU�n�}��|o���.OJ�,�{��
gӿނ���h���a��8F ���b�]9�ػ#U�ϳ[�b��u ��Ֆ��Yw�~�G͇ޟ�*����\���q�b�HF�r
oP~�-�)�VNA���t��*\q��ӭ��i���,���٦����p#n�Ey��F����:%��g��CA�#�j���f�����*kKַ�&}���o��a����z���"Q��~���`�kܺaF�hj;Z�4�XGA�#4:��r��׬Յ�:{����UPT�tG��v�,KB��l�������
����N�,9��^K������_v/xn��{�0��o�Y[���:���p2������V|S?��E��'o��TO�����$��~s���TY����#	�XlZY^��kV)?7Sc����Z�η��(]�� ,N���٬�zroA�������v��=�i�A���	̷n���E5�QS�f5�ܦ�㧴c}uhzf���W�f��y갼^��m��iF�R��T�Y�[7�
�DZ�$x�|�۫�v5��>:7}�n��,�G �.����p��Ou$�9�ػ�귶��$F� `Q���-/U��H��ܤzz������v�,�����^�ˋ{�H���¯��n���lAܫ���t��Ia�x�����)������0�E��~k{���k4��O�-��Ƌ�6YfD��u �ht}��9�/���xhZ�BO�����{I	
rd�PY�M���I�:/$�ىڛ�T�UGނ{�Iх���B�nm0�|����)\x�Jiz���BdS�fISm&�0��o���=�b{�7���{�ܧ�6�٭�E	�P �\���5������a"�k��~�&''599)[Z����,�P�z�vh�3.Ir�����}Ѕ�?�;�pQ�T��7]��eO/RM�N�mܺA�;���Xmy�Zp�)��+f7jܺA-��q��r�30[p�{��`�kz�Ii $�Ţ���{���ܧ�6D�������ܧ�ט�����~�t���cM ,ӫ_�X_ڬy�=���@װ�&�~]������5u���rTV�gs��|�	Ym��y'd���3��j�Hz�����t�i=~J�WBَ���/�r�S�5�o}�k>�~�Ѻa�G�o�*�����3^�0F0c1���G�Pˣ���8_�;���q��� `f���zW�]�O���@@����uM?���Z,�JTg�h����}�: X��S�ZP-�ާ��aGꂁ@���9����u����b�)7�B����h��#��s�5��Ž���Q�h��CV�`J��z_]�N5l�	��u��Z+9��p�u���h���צ���8wQ�����nPæ�ｩ�Z?�$��1 `&��Xt�d�;�1��$}˳�۷��j�J������>���o�$�\�g:9�Ju3�����Z��z���4��}5���Rmyi�}��nPS�fu�����9��>���F�mGB#s�jԼs�T��W"j��}�Jݔ�ٌc���O٫bzO�M�����^������ׄ{0�z�d�������  �+���"�|���u���`�����T��Ֆ��=Zc�Xd�Z����U��5�/�I�E7�jK��M  `&�_�"���7����6ը�T�Z�����2�n�������oPæ�?u�i�N_��kg;?�urT�Mv�-����z���eM_)Gza�kpBҙ�� �rE��E�k`$�^���?W��ݡ���~v�װ�35%�J�pS7���/Å�?�  @��Kk�R�5u   �ǚ:    01B    ��    L�P    &f/))Y��������8��=K_q�D�   ,Q��   ���    ��u    `b�:    01B    ��    L�P    &f�t����1U���^��>UϏDFFFaFff��?�����⾧;@�N�7�M    ���/�גnJuC��>���������z�����O�    0\    &fOu ,]��"��ޛ�f   ,i�: 	㷧�U�2��   XҘ~	    &F�    #�   ����   ��T��@C�o3�*=_�P�j��G�   `g?PqW����Oߑt�a���    ��q�u}��[
�.���wT8h�h#�   @�4nݠ�m��n)� ���   @�d:����*��P���Q]�]���P    �wn��e��ڎDu�RtA�;
�    H����j?��5e�-�@T��;�H�S�9�Q_�H]��Ҿ��6    fm������d����:B]n���Wz/|��v    �lL��P���5����:9�Nus    \�V��U���7n�G�'���>5�E����f����T��^��qѰ��F������댮R   ����1�S+W(=}n����ٳ�
������46��ʕE�?�T�~��ϝ�P   `	����a��:k���w���+Q��ΟTaav�����$���    ,~������y���|��~6湉t�R    ���   �T?�E����0R    &�H   �%��%τwƱ4�_��i�}���<�3�kKK�s%B   �%⓮:qp�q�զ��I�	X�t}����<ע�Ң�<s�s�    H ��:I��}�8,�w2��1?�2��zn@}���O    �����#8�'����3#�>���:    01B    ��    L�P   `Q�_q}���4~�M#��b��P   `Q*Z���nKu3�o����wk"=+��	u    ����t�   �"�T���N"�   0���
t�   �I,�`gd��$�!w   �$*Z-�6�\:�����ut�   ���^T�k$�͈Y�ؐ&�u    �������+�͈K��H��ʨc�XS   ��B�����r/B   �Eo)� ���   ���]���P   `�Zʁ.(�`G�   �(��~��]P��({l �k	u    ���T7!��Ƈc��P    &�>u    L�s7��]��d��o�n�:O�׻|j���F�   `j��4�tj����ύ8�=:{�W���S���u    � �ΟVaQ����!��w���+1��R��?!�   X"���;/��?��?��f�
�    ���    ��u    `b��   �d�����8�f�+==mI>W"�   X">麠���Zm*+-������熞�л   @�Y�7XI���S��ay��K⹳1R   ��>>}>��|RO�x�l��   ��1R    a��7�aS�
2�Q뇟���H����0R    !�wnS�����sU���ƭԼs[�[��0R   �p�5l�Q��Sj��/B�ZP�j��vD�.ς��_q�r����ܔ�[m)\ӵ��   0\ݍ���?	vy�z�Ԍ�2T�Z]�ݖ�."~�M'o�[�Y1]O�   �4]�Ψ�_��.�@'�    ,rK5��$B    Xj�Ψ@'Q(   @U�i����;.I�w/X<e�h���T��;	ik��$B   �j�����"THe>�`Wr��K���m0,�I�:    	�q��5���h�V~�Gu_���G�   `���5�1��g?Pq���M���.y���[}�!��P
    SX
�.���p�א{1R    a
2j�T��?Q��H�X㶍��^�a�G-G;���n)����/�]Y';B   ���-/U��� ӡ�Ag(Ե>��j�KC��U�QSQ޼k�b�2"�1�   @B�<z�$����?�$5nݠ��R��T������W�q��mTA�c�=�r�������b�    n��jU�����|����su7VH�������P���4���z?Z�.���w�=6ӵ�:    �N�l9�:V��P]�u����))4�W��1��c�Ih��5>�u�:    Iz�zRܒ��B)    7|�-I�,�m*�c}��?�������nX��6W�f�?޸�u�<�w?�4�g,���F�   `��h\��jz�*�th��ju������.�<@s:�re����F����=۫@�؉��z�l�:    ��8wQ-G;հ�&4'MU�j޹Mu�kTY��+CL    IDAT��������u���
��e��Q��[~�_�Y}����	�   @B4��Mu�h��j�<j=~*T8%8B7�����3�^����;/��?��?��FI�s��    $L���n*>���G�P��S)h��B�K    	S��PS�f�U���Z��j޹-��#u    ���T-�ާ��|Is�T競�T;�Wk�~皺勑:    	Ѽs�*��`��ޜ�+����vD�5��f�3�]�pi|Ɵ��IC��+1R    �ר����EP�����5nݠ��5qmL�I���88��jSYi������zNB�   `Y���B�B�.,��&Z�V�����wqX^��#g�z�l��   H����50�3>>}>��|ROo\�Y,ϝ��:    ���`���ω$ b.B    ����X_}�s��P�26�:    ��8wQ��O�q�5n�0�y���O��U$e9cM   ��h�ɛ�,�WS�f5l�Qǹ��tJ�*��T[^���|u�����6����m�ڏ~%�ߗ�'�Ǒ�K�T�t���,Y���[g��P��   �IA�C��6j�-7�Y_�50��?Q��i��	{}���%�<�l���ޘ�'�E�P   �'82'M�H��-�`o���~	    I:�]���Dz�N�|��vF:�P    
2Qo&��q���0�Z�3*�I�:    	Pwc�Z�/�k~��?5��K%��$B   ��8wQ͇ޏ���	����bmZ��Z�r>J��R    ,Fl>    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01{� s����5=�RZz��2?�_#���T�   0�q�8�У���T7e^�/_V mT"�  `	b�%�666����T7#�˗/���?��    ��:bllL�������������@��   $��SZZZ��2::��&    	G�ò�ZT�e�l�,G�N��   +B���4�ʍ��YRR�����a�   bE�    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &fOu��
3��ސ���C���ci�����|�c��n  �]y��+�R݌��,�zzc�k��
=���X
c�����f  `W��T7!*�:,�>cC���   bŚ:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� �P�f�Ck��_Ia���/v?    V�:,�t}�q�%9��   ă�    `b�:    01B    ��    L�P    &F�    #�   ���    ��u    `b�:    01B    ��    L̞� ���Kg\~����v/    �:,�~}�g¸�\2�^   @�~	    &F�    #�   ���    ��u    `b�:    01B    ��    L�P    &F�    #�   ���S�  rm�Zlܗ{aN��߳#��   ��n�������F\~C��?i��%�n�=����\B   B�2qflB����o֐O��   @�XS    &F�    #�   ���    ��u    `bT��i�|>��n��~�l6eff�b���Y   @R�`J>�O���
�$��+�׫��\�   ��_�nw(��|>MLL��E   @j�`J~�?��   �RE��)�l���   K�����)�u�oZZ����S�"    5(�S�X,������D��%�   ���e�X�p8":�������۸�|θ{   q`�%    �#u0����R݌�ݮ���T7   H(B1>>����T7c�ϧ���T7   H�_"n�5�I���S�    a�C\&���-(UAIy��2��_�Y��n   ��:�er�u����W5��    	��K    01B    ��    L�5u �����A����n  �p\��&D�P ��seU��  ����K    01B    ��    L�P    &F�    #�   ���    ��u    `bl> �jJ��o�ָ�:����g:�t/p%¡? X~u R*7=M5��r��c��e�m)l�yџ  ,?L�    #�   ��1�@T�\�*�՘˘�YΡl��������\.��*��D���ONhrx@���2�{%B�k\�?9��˗��Ŏ4��o[���CǼ^�F�n����}�I�Kc�C�>�x��  ư���r��VZ�����+*��\Y�7�\s��ۍz<�(���u�~-��-��<E7����ؤ���T7e�  a)��:��~(�m����T>0���n���oVVV�$���L�C.�K����$��ŋq?o��d�gFF�._��,� ��lY����<���'�===��'�a��7���v�r�-��?�3�p�*//Waa�$͘&8��������&&&��ե���9sF��c
&�%�,������ٳg�D ��-�PW\\����<��?�?�KA�$##Cw�}�n��v�|��r8��H�|>���kddD:y�~�����O?���"�'  0��`�C�xV�������l|��SFA���Mx������!MK�XȪU����k�ƍ��Ϗ;x,dhhH###�����~�;���Gt]���	  �Pg����r��p�je���z�r�\���]�����٣_�V2��4��U�V�G��͛����@ ��VNq�\�������~��_GF�Db��G}T_��Sڟǎ����z� ��Y�.Uk���Ҕ��-#u���x4::�����s��r:�S%�P��&�dggk���)	s��\.}��gr:�:x�;����
"�'  H�e�R���D���JKKKe3�˥��A�^�z��������'�۽dB]��n�����׾�5egg'tZ`��N�z{{500����/X$�A$��|�ǔ��C ��-�!���C���EVV�#u&�~�����y�������D��$�.q" ���z��'��C�f��t4)�á�������v[(��SPP ����ߖj�4�����	  �[�i�P�x,�Pi ������|G��r�|>_[�ժ��Y,]{�*++����Þ�� B�  H�%�6u��ru����K�>������h�|������)�á�7�>�����"�'� �d�,#��E@�mۦ��~ZYYY�	 A999���T~~��y�egg�=���R��O���b~��'F�'  �:B��E@�|�ISoϑ���믿^iii	"��\;  ��	���������T61p���ʕ+<���������Ą�_.� 2���ҙ3g499�={�h||<�y�Vq�?��O  9B]�|>edd��΄&''5>>����ϛ�������7U��4��]�V��������$�.�Ad``@���w�=/� BN����VSSӼ��  H���b Q�$���g�UVVV[����*++Sqq�{�y�N�����9՟��'  ��X�2�� z��'URRb�"�*,,T^^�jjj�iӦy�+..�Ĩs�{џS�YXXhH ��� �q�}���n[������L��k׮y}a���5�\#)��	  f"�����Z?�pؽǖ�ͦ��2����'�H�3�[�Y�&��	  �"�����򗿬���T7%irrrTRR���r�[���{/�����LX ��u B6nܨ��k�O��k����Z��G,�Oc�  �G�K �Ͷ$�X,Kv'�e-##C;w���MuS��f����D^�W�a�=�Oc�  ̏]��b�hrrrɭ��Z��X,���,��V�|>ߒ�����jݺu���HuSR���D������ׯ���G۟  `~��
Kr��|��n�+==]�E�@@~�?�-C��v��o߾,G����K###ڴi��=��Oc�  ,��0�����˗5>>.��#��*�����5�\�[n�e��"��n�q�q݇��bT ���>�/�$��jbq����+�����)������<]w�u*--��>����  ,�P��
r��r�\��wX\���USS�$�
�"??_N�S_��c����)��  W�O�H
��/�˥��IF����UWWS�押�<�|>�_�>���ϙ��O  pu�:$���._����ȝw޹��~Mg�ٔ���իW+;;;���ϙ��O  pu�:$] ��c:fj��v]{��Y����v��nݺ���?�������X��	  "CiB�������f3������:+oKQk"������J���Ѳ��u��]��Q_G�k ���R�gI;�ͦ�˃�nF�


�f͚e�A�|rrr$I7�pCT�џ��ڟ   2�:��R	vf�j�*
z�#--M���Q]C�/��  �aA�ǣ@ @�$#����p(///�k����ҟ   2�:,���<�iq�+--M>�/�>�?�K ��갨�\.��K"*5�/==]n�;�u`���b�O  ��aQ	r��
)�����jrrRn�{��&''�!   )E�â������NA   ,Z��~�=`�w���Y��X��
��b��D��P�EirrRiii���LuS   ����7�����w���?��X��m$�ٚF��,v%j��P*vQG�W�΋�焯jܽ�(�!,��=lv��E�[���L���oþp�C�2��]j_%G�nD'e,%��&��-r�^P3�(��ΐ�~���4���cZ���{� l&r���Ƃ�~�踽�b�
���Cz��I�;�Y�2�eɿza,\�/�ŗ� �@ۙq� �~��;&udZ�t��:"�K�����n�0��,�?�����x��/����u2��u�_���Ů����,��?h{��X��v���Q-�`�K2�Z:��j����Қ��Y}��E���Ç��Ԅ۷o��1���ʙ�z������.ڛ�����8��gB�Nf�g_�_�y�,c:-Jn�:�ű���Q_�	Hh�� S�d25q���ں�k��L�ϬVVV��imll�b��4G���ʙ�zu�DU�?w�/!��2z �^'s{��S�1�����WǦ�����PZ��Z$v\~I��N����Oj"i6B*�*yo'糰r�^��_�k�o����Bu���y�4I��dV���+3������X��EI�:6�rn�m�İ t��<L�X<G*���e�Ւ�d����d2Y��8�;+w>�ٕ����P��ש��@"��<�H��WǦ���Z �U�s�#e2�ZY�Y���8��鬭e�A��Ζ�8���ʝO""�j� ySǢՎ�r~,$�}<���2�,��èK�D�h�Is���U�۷��~I��|���$""�&YƵ��c!��/�%���x�A����_��IH���U������|����<�̧����=""��TF�:��cqY�|�<�wT�GI?��կx`�L&���|��Ge=�����|�t>��v� pr�β��Q�e�̈e���/�˩�1�#jp������e�iii	{��){�W<�|�t>����A���c�,��~I5A�$��P�VWW1==�g�y�t���.�H������/�z<�s�T4�fao���œ눛��<=��ن�_���{��|�'��}������� G��� 89��cO�  x.mm`:}ng\���h���'�կ{���:^ṕ�7�r��u���W�cj�����ف��_B|-�_\�������9������?r���7��Kptv�s�-�#s[����q�?�v�^Ͽ��焫�K�Z��M&n�<u�#��R��ւ$��K�/-J�=�8Z�c��QM��V��������6|uiccKKK���X]]-�y8�YXYY���|E�Y�o��#��@;:;��4k%�{�����\���y\җ��w����7�:}����������7��<�^��$wv��:  <{��mq\�]����9z��7կ��=�n�w���I�u�f�/>���|/����aDc	�[���-�,N�xsW��v�d���x����W����z�����\���Ww�#��� w�͒?�*�ukFF���K�:6�~�b��s���j�,�쀩�{��arr�����/���}��������|fi5��8:;��߮��;ث~R�5����]�(����w5�I�_K!89O�S�R�G���l�;��0p�&����V) `j~!{��G��;؋xr���G�_wtv�7�Z���:�[��(�����$��������]=��ȅ�#��QJy��d���ϏB[ө�x_[MZKQ��֊,c��w��D�I!�N�ʕ+��d2<x� ���wiT��jm��ZΧ�n�Fpr���7@T��k)����-����!����a���M���ݥ���~���A|-��{GIDɼr+j����|�X��7���U�>'³w�u�f[Y]{Ky�+�'gv\�,-ͭL�F��[+�(��l�JM4�� ࣏>���߰��!�"���I���裏��{�5l���|U�����^�g� �ހۛmE���g�l��M�/l�u;{05��pdnK��݅����b::;�Pc�9y����jUMY������E�Z����lC��mDc���BJ}�k]iε��M[5���TSA�:��������7�7�,��`qq�dR�$d}}?��Op��Q�g��_@pr���C!O�n��$ `oi*�9ów�*���)7��X��.�#sp;{v�KUh�f~����S���yy��L� ��f)	X�����u�N��o���5��K�b����Nv��A���BU��_����������uki5m�嗒(�E��u��3�������D"����w��d2��S5��9�����D���|j;�;��4!pr ��H�^%1+�r�U��H���7���F)��I�J���CM�����Dpr�`���F)J�{����եQi#���MG89�Vn�#sN��7<��q
een2�u[��۟K����L��N<u��%��zݴ]c����ӨKت-�N�ҥKX\\l�����
���055���/Χ�{颱��u��=�})���%�?+�U��(��q{�S/��ei��d�ꏲG�X�����rM�1�����-I���N醩�2��Z*۔�ن�<?�Gm���K������J[.�<�xr]�v�sn.��V�s�����J}�Gc	��b�[k�V�tR"Qݥ\�J�.���X,����A,3z8������O?��������|�'p�fիc��&8:;ؐ��'gԆ��	僃��������V�$N�����Z
���E��q�G�mk;O�S*j�+׷��
�:���E��|�':}b[�47�*�� ����RI+t]9˗�zݴ�:�	�R�0�p8���Y�����O>1z8��x<�믿��9j
�'Q��_��M�N�@���-gw���|M15��=�+����=Ww���J+��BG�7ԏ�t������a�Ȍ|���N����Y����t)	���+{v�G�($=}�]�J}����.1����䌚�z����n[Z��^�6�ba��AJ�2�#�mdY�ݻw��3�`qqKKKFIs.�}}}�Z��/̝�D"Q��jΧs�؞(�P���\  BIDAT�)���\z+[�x�Y�#_82���;7;��t�������#�N
5J�M�	��	��4��f*JI�vJL�%������<�_��]R�YS:izLh:�����;>�����^���|C�p9��1�끫7�<����׭�R���.��:u��!��j�j�8�r� @Ū6�H��X[[C[[[��666 I��կ���s����E��{wnWl�o����G^��ֆ��&���u��9���Kx����o�vyy�}�[XO����p>����
�����+�������������/!�+��b�`o���+�!Kd�[��|�'���qQm�����Q���P��w��_��V���,����hH���hii�7��M������0zH{�'��/����ʾ�\���ػw/�S'�f[v�[K���t�;jz����� "�mб��g��X�� �U��>��/�����X���Ckk+�}�Y�ٳ���T�'����Eww7~�ӟ��+�q>kH|-���f4��c������Sy%"jD�\z"�#o�`��L�	�9ܻw���>[�&3% �������B��7��>rP�6:5��{#b��߷��;RǢF���̸W J>��I���j��ޝ�����~�ݻ�������n��	s�\�����'�|�4	Ƚ{����Y�����i��ԛ��R��WΦS����g�N����v|���|�'tI���ID�a���JkP���q� ��rʤ�L�V*u+++��ں����yҠ������hjj������֭[�����\���nA�$�A���E,þ}�jv>�|���z��&�`Z����o����y�Spr��j�o �'������59H������}�`��{N�@��'{.���\zK�$ˈ�Dd.����[�n��T� &udb{��a�Z__������o���|��)��v��N����x���ҎVVV�L&100��,Q4�@<���g��r�O�WTEs;{�9�=�|�\1�ȱl��Ko!��B��	�G����F\�]�N�;Ҽپ}�Ͻ��V|��1�ȜD���s���cSՌ���G F�}<�:2-A I��àH��h4�'�|_��W��_��Tg���v�����~�3�/�$	w���|�(p��p���D4�P�y�7����BprF��g��?r��.�Ԁ��5t���ߏ����lI�k1&�� tX3b��n\�W#f˹q�(��J��I���je��ܽ{�(��v�Ν;����L&������׿�u|����/~a�X���ԇ����%s�{����;�״>>����%�k���*$v-��]VI���R���Licc��q7J�LX__/z]:���b�Ҩ�I�ڵ��bdd�H���UMF����tbqq����*��,���	�P6��;d\�����X����<G#��ڒ$���_K!�,��B��ē�L,��4�$v�s�^��b�;;�%1XiB0�#E���D#Hg2�WCWWW��'�����'�O>�sss�{��f1r555�駟�7��M<��Sx�����Q�8kkk��Tr>wo7�[ng����-�=}N ����b��U�D3t�6|��>�ݯ��H#������`/<}�-�5���ݲ�3x긚P&n����|ϥׁ�F�$"��Y%1�v����~XVW����7�����.�:2Q��5��$�i�^]�������������a�Z��"�U��455��p����~�iX,ܸq�n��h����q�=t�f�Z�900���fD"ܽ{�n�s��Gf�g�K�#��������	'g*��4D�S*e�/4ѽy��|C����9�Mb�Rj7N��1 ���.���b�<�݈�DT�C���3=A�W�|mgƽ� ���FC �F��2:t�m�Z�=�=A�N�M��/�� �J�����u��˶�6����������9Ċ������!<xP�f4� �w~�w��҂��%ܽ{���H&�XZZ����n��n��'�@WWzzz��ގ��ܾ}��_^^�.�����c_)x�Q���c��/����l���`�����a��=p���l%+pr���o��{�Ww���SO�f��ܫ&�J��WA�:<u��v�A�>'��?�������VFDD��2�ɐ���v���6:��k�xA�i��)X�#S1CB��<�;�{�H$tODdY����YEtuu���v� ��������b�ǿ������}�>��3]ǘ/�L"��m��!]$���OeNͧ�b���>|�>��ABWL��M�:GgGv��?e_�w��f�nU2{K��6�5�#sۖ*�A��Dc��؛mjsV	��A� �+~,��xM�� E%���D���nA@ �:.&ud
� `mm��a4����o�z26����ê!������qUc���C,..b5��M@�������AI���:�sS��Y	-����=�F82�m��lC���o���t@�b�v���Ec	u�`82��tD�`˾�z`D���jY�F>�c���<"2� �9A�s�q�77��*��dRG�cBg�ŧ~�O����֍5H��t&S�18���G��e?���~��}�6���#����@ =��.y���S��Ep>���n�[�89 [U�7���_�xo]n<GgGիb�+�|�yO߲����D��0����߈ʕ��e����VM�}?
��C"z$&ud�zI�������o=��-xʰ���_��aߖ�#��8���(V�W��많j�4��M�g!�X�����;5���bGg���������*B�x7��^Q�2K��7���@��k�臈�:2� �$���ՊL&����F����ެ��T1ng�#�Ԋc�A�z%t���-q�J��\U;���Tٿ�r�!��7�`oiR�\��S�LIGgG�^�Qg[*��Wy5�Y�L��,R��.�߉�1�.������S7�ă�3�7���s"x�8��?�M�n���FШ����\U;�����lSv刊\�X�n>����;ػm)s4�@pr�n^�"x�8<}N�g�����I���z�5��]��=��9�f���}�M������D��_|C���;7��*����	�8z�hL�j!�S4�LB��� D�c��fXͩڮ�&�LWw/Z�h��TZ���*�ĵ�x�����9���8�Z�J�����s�7< �� ³w����X��Q�2�ZO�#�\�~8Q଼hgG]$;��~�G�!�C`�Ɩ9v;{����K�#�gD!Z'�~��TϷ��"�{�������c6϶T��*�� x���:}���۾noi��ϩ���~���^�瑲�AY�`o�m���^1���`u�
�YH���F�n4�|O���A&n �S[�+7��Ύ���t(u4��c���j����_�6E��O�3{�����MGt��f\#*WFV���;eI�N�.��3�*,��=z�>�#�S:�j�;؋���}�u�x89�k�LIr<��R���7���^�c�ów�9�mń�ϩv�՛+?�����f&u�+�ł�����;GD�|�}��m#%		��<|C�e߈���[Yf���;���@��M�JN��Q�j�j��r�\,v���I�J�� �U�Bϭ����X�X�����v�Ճc��s14�.OL�4��� L�y\�������͹��_���S�!�֢���oX��k&L�Hs��$1�#"]){E
-G�7G�~#�v���P<�bdoڪ�߬q�H��L�]�]��>�z�S�u;���P�Z]Wx��w�S��$W��٥�:�+�/�SϑT~F(U�����ȏ�z�5�{ng|C���sh:���F��	&��z�;ث~ �,�MG�+66_�s3&uT1Q��(�2��4R�����r�����rtv pr����_���zc���ܛ&=؛m�A��.u9dprF�O����/�8�ju��FLGgǮޣ�R%�_���q�i����4�k)�.OTe�Bٓ:}b����t����^/��_|��
��]{�������h,ϥ��9�.�ԓ�G!��=puw��ݕ=Sts�|��[��}�m]�`�*�q^}�r[�֫F�A�$X,�AH��l�,�2$IB&���$.�� �J�����u�t��(b�?�����vS������>�]N�s`w)��6L��7�\�u���O�7<�h,���}⮴�w9 �7)1:�"prX���	RDc	]MSI빂��܎�
e?[�+�
=�*U�|��l��Ko�����<}N�g����U�yV�{T:�V��7w�`�_�QX�����2��٣V���H;��|�o�Om+Y���tz.��pd�����g;�uv�]��v�d+�U����N�����}Z��3"&��B3��ԃҡV�_֣��N�7��5?�^{��6ڛmp�oG���sh:�=Ba��g5��V&��z� �1�#"������P��ܮs�P�JwKe����U��[pr��5=.Wi6�׍��g/�S ��<e���/�Sa�� �����+��_���wt�˸�B^[:?�eRGDD5���;�޶?G��f���;؛Mb7�f�S����B|-���͓{�m�YO��3�:(���Q�J(dj~�>'��ܤ3�Q�I�R��=���O��~v�2n�Q:��/�����.O�庺T2�|$=T��?r��~� �h,��郒�j�`�[��N�S���g�s�<0Z��s�'�y��LUc���i�9�������Ҕݧ��Z��p�e�Z�k�܄`RGDD5J�\�$����W����-V��(�l7��	\�	���j�,����ϩ�M�!�@v��w�WӤ.K��YT^_4�@0�:���P?��՘�u�����S[�+���
θ�k��F�O� &uDDT������r�Զc�����vـ����-M[lG�%��^B]���+���[�##�#s������Mh�D24��x#bc�9�z��89�P?B��޻�˸�h�����J$�~Y�x���r|C�r@�w���c��!ttv`�� |��[����&s���e�o�_������j�é��TZ�m3"f���T��z\>���P�V���.O�t�q��J� &u�bRW�����(	�rV�B阨Wg7�X�l� ���%L�����|C��l��=�[��4�<@3P�*���qT�2n�)��L�t5??Q����F �22����+�eYF[[���ˤ��teo�e�gy]7j��r��;��٦&����S�SL�`����^�r��ۆ^�3.��j\-=*������?62<U��?��Ƥ���H�0.��z�J�&� �$""""�0�ƛq�lv���~IT3d�daRT���([\� ; �-�3h�DDDD��R:�I���2�ɐ���pq,^�Ұ�l�㎽�Gd� ��DDDD��R:�I�)�2�eɿza,\�cSǢ)   �vf�+��������L�LE�,��/�0���-_bt<�n�0��s�QG����O�����G_ȸ�˸��5J��3��w\����������x��AU�~�k_S�<�9u5��s�V�&���2��ɛ|ul��'*`��q�1( z<?Շ}ˋp����� �2���D�c���#�U������f��f�1��A�t�,�����u�$��x��饌�ƅ���*�r~,�rn�m��0;""""s�4����j���Ts+���ș4�)$�[�_�� d��XJBW��&���M1�#"""2-:�I��$�3���CF����2�H[$���|�WǦ���Z �U��DDDD��V	� Iݣ��E�~{�Y9?j?{�"���nH��t:���	��={�0.�2n����q�;��L�J�ؑ��2��\)-�ۭ���0�QdY�Ç)$�Ɋ�KE8�2�G���q��Fi�yf����5�:����O?�4�{��w[!^����R�k� .���3�>Al�8��A��bEKKKE�H�_�V�uW�D�q��Fi�yf����%=: `[F"�2~��85z�Ƃ2�0zT�_����ʸ�˸Տk�F�gƭ︕�+���B���c�4z T;��E��/P�e\ƭ��N�h�̸��\z&t@/�$2+H��7n/]��(�H"�ЮY,V,..buuuW�>���(�2.���m[��3��w�R��LꈪOF��!�J�:6�~�b�S���)���n?����q�v5�<3n}�ݭj$t �_U�,��G<��M"""�ZW��`RGTu�(��C>S&�DDDD5��	��������H3�N� &uDU��6_Ǔ�C"""�ZcDB0�#"""""҄	�����Z�p=�|�$����IQcRGTef��	����DDDD�;Lꈪ̔	� ��C """��X� Q�1Y�rn�%H�0zT[�v;���vumkk+�2.�(�Qm�����:�*��}g�=+��BF� ���5zT[Z[[q�ر��J����ʸ�˸�5J��3��w\3��K"���)������ڊ��8��V�'��˸�[y\�4�<3n}�5+&uD|�6:�0zmgƽ���v��_��r�2.�2n�q��h�̸��̸��� 6�L���u��vA�ŧ�!Bſ@6�@v��2.���(�6ό[�qk�:"��3ro]�U��JG�!�"�V+b��2.��X\�4�<3n}ǭL�$B��w'_��f�}g�=0Z͘T�dY�Ç�q�����q�;n-��:"	@�5#1:n�V̖s�.b�Z񈈈�H_L�&�k���j$v-��]VIs�%Q�`RGdJb�rnܥW�}g�=L興���`� jE��q��U��A�M�,��/�P������ͦ(�CG�����7��O����v�e\�58�Qm�����8?jH~Ťn���Q5�2�eɿz~,\���
���C�����
0*�c�K"<g�x����k2��r!\��汶�q�^��#���Q�cRGdb�����uX�c���k��0)*	��^'�� ��p� ٠Q�1�#�������G�f��DDDD��/w�ҽMDDDDDT�d׌�ͤ���i��@DDDDD&$`ʨ�L�J C="""""2��(��ͤ�˙LPF��������C�q-��+u5��X\��ݡ�DDDDDT�2��72>{啡��ũl�x"""""jd2pq�����1�RW����f�""""��&���L��sq,���ֶ��������Y��=��/+�v��|� ������d��$��αfR���q{���L�������|
 ,A
��=�|�����I
    IEND�B`�PK
     B"BY$7h�!  �!  /   images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.png�PNG

   IHDR   d   G   ����   	pHYs  �  ��+  !�IDATx��}	�g��UYwuuU�Q}��P��ò�[�c3> ��L�L0��%v �`� &�{�e�X�;,`X0�c{| �u_�:�Շ�w�}WV����է���f��������������T,��~*,���t�4]М�k}��%��n �-ȡ(�a 5n;*�t����I��p۬�4(�-\mPh �����	+�~'�oQPNľ�i�xcx���Ώo�ƽ]�hvP�i �BQ�vBI�M�O�os[��ǣG��Z��):���H�Wj1
�&�&y�G�P����
l�]�!��kjW�v�!⒥vVjg�/9j�c.;�S��8����������Z�!��Z�r�Cn���]�(�v)��dE�c$ wQ�e]C��p:�X&��ܟb���g�ѳg���ƪ=7�vp�"Yj�͛���4��2�ES��t���#�bzj�u�PU��F�q9�ZU�h8�d*���F
����6X�ǋɉq4��L&O��pX�V������ ��)d2��7 ��c��U���r	>&@e�譼�l��Oc��;����u���F���N��?3����&\nL��C�����!��#	����MG�[�J �ӓ�SZۺpr��H�?E]��e1�Jz��4�,X����n��>�~:��~�K�"���~�z��g�P��Fs��� �ɑ����,l���CMu���MN!�&�"��bdl���̂������ëZ1�A�u445#G�G�g(�NL"TgEU��D*���I�Q���(*�T���pvzfi:�]K�P�6��F��'\��kUĉ�����������D�����4�����>�������sb�b���ghc�&�2�[��_�gn_U�	�-����/�J`�e!s5�w/��6�MiW��������9��V�}E(Ni[o5�vˎ�R$���������Ϧˊ]{��,�S���'X�@M-��ד頾��m;wR3����]]�kE8HJw�|Xu��6L�2�����9��2.zf����ց���Ј&��I W^ú���zNim��Qơ��7�$��Q�Vw��K�x�+aH�/��D�ӊF�!��׃�-f�^�����6�0�
�Ȟ�T�i��b�#��]{����ؠ>�^ ��yltR:���������TN��Ͱ�%V�l������D}b�^ ��P�!E�?I��٭"<S9�G��4��Ժ�ই��E���*8cYN:_A�K8S���������	�T�@8����Z�FLq���fY������̣�e�,�8�����+e𙭝0�a�� Ǿ���*Ih��!b���΋VX�T-���܁�;3q�ܕȸ|�OC'�W�"@��\�7����8hGM����?u��c�L���at��X�ž�!��u蟎b8G[�_��|4��σ�j�ʹ�r׭n� ��DWc�^������Xa���&���i��n�h&b��������p��)2Y��n���(��0ZCU������R�St~(G�cS|t6V#20
�|-ɲ�&��޷wv��K'�\��-���/"569/Wu��yr��ܻ6`Cc-~�IK�tQ����a�������Q�`��8�?۹��n��p��ÉuV�omD�ߋ�Q���y1��� ��"i�A~�D��"���z�H��Ɉ氆��۸�p8���ؗ��@i!JRʖ A~������훘�1��EX&#H�r��
��9'�#�]K�3u��dV��M�B�U�d�tznT�gת:��;���_CX�;~����UȒ�fHz�^?Ԯ �������&���!	{�yZL��Ldɜ�p) K���5֒��[%3�����;G>�FDIҀM�SD��``��찘���!����vS������/s�� p�:Gj�'P�/�&�M��i7�nchb�f�@)G�Dc�Z$�ŋg����I�Tx�:X��3G��O���
4��&ȖO�T�J�w�ā�29�R�f!O���T��pD�3���H
llO��g���J����A�|��Y,��q�LG�$5AB½k	���e�>6!�E�p�(����Dd38�~�)������89|E>�%!a3�-1�+K2䏫S8�y`3����h0i�
=��*ND�񲽎.Ē%FL%��$�f0��y=�U:pa<%���'F��T����Q"3�0d`�/Αy1JQй���Re�G3��q��_��x#fHһPi��3׍��Hr/E��v��}�E�H_�}g�_��H4�
�7���^��&�7�/|�3�r:�����Q�mU�R���J7�F5|;��hO�8'.R�މ�t�U��6���cf�.�Fj=�'��
}�"CIg<���k��i��XZ8M��7�	|90_{�Y&�R��kT��X���cqS�8�`Ma���f��%F�)
�@b��͎��o&~���^��b}R)�~�����i3��[Ŗe�d�6{��2wŹ:?̜6aP�HD����Z����8�:�*�Đ� MQV�� =݃H�zd�������)�T��i���
���0m�n�m�ߪ�yE��ܰ��R��H����,6Al"��EÊ��!��33x���}g�Ŧ�}�!>����^��߿��`������f�q��9��@w���lz7]#g5s�����M&*�)�e13H*�>BG���)��ό\Y����m铲�L�M|�Z67L���c�3��i3���%0[��^[W����3����;���T����.m،qnB�1J݂����&Sf���.�A�b��� �HI��?,�q<�f�M��#�j���6F��$�	_�4�N���_&ЅXɳ%�d�&����KOh6�ia�3OJ>�$if|G<�t�%y�|�d��2��Y%fVy\r�	X�r�(0�����'�e�)K�+��Vg1��o��;RrZW��2ODy�3�¸!��
��Y��̌:��a
(�9�ϻף"�	��_<�,�;O�.�:,�;���={$�LPd��g��[��_O���ޛqφ�T����'��S�"���6Y�_�f�:��x�#V���9��
�6��O��i�_�TpqYy�J��gfwi)ib�T�n7��8�**)y�![�#����(��9�է��k����������ַ�k��6������|O~�����>�<N�Na1��o�h����I�vܷ�/�_ ).P�8�5uAѲ�(9�g�͉a���7v� �Ç����s��5A�����z{°��
�;N�G�+n��+2�W�,�y[�����6&��{_L�*k��g�p����?�߱A�;���Dߵ�_y�5��F�v9(b�r����V�{w�7�w<�OߺYL3�����%ʸ�.'��Ղ��g��˓��f(�v�QM�S�mg�r�;�S✍33Ù��y�1�Ḛ��������a>��w��|��Ib���~���q�??&����;�Dy�NSҹ}U�� 9?!�R����&�Vv�ϝ�~����!��5�)'%��p�n1W�f9�˄t���;���g��`&��.:XӾ�g�,��O`)e��&��9$-w�5b߹Q|���bj�8އJr�~:"�񼝋r	6�����lN��a|����>1�E�*���}��"�eq+O�q��eO�����T�t��4���@�L&�a''j��LL�w_;���s�H�ӽ�"�~/~��$0����>x�����ɡ�����o���i
8*ȇ���,��5�w��sz<�f�O�~6i��L~���)�oG�bKkz��1�|�Qr��n��l
�N;O_5��={:����	3"Q�kM67Ւs�P���ϒ�'v���i�E������I]f[9�������XC��~�%{��Ħ���������\�W�>�g��)\Of��������L���������DX�88`����Z��x��1ay"��hR��I��>�έ���-��()��ǑD@�ߤ)bc�V0�8�i:6ӱ���WOCs:��o��M�����H�9�KĲ���K�$>zC'�m�R�x� ��et�cPR�D؟���Na+K��<�~r��0�CZ��_�S=��]2M��C�(2�EI�����'�%�[]���5V��7J�������sp��Ϯ��m��ZC���FN�tƇ��G�Ã��g���׷��J������ꁫj����aUE[f�(7����Ȕ��(U��}�~�L�a���������x����)�1~��*]v�b6L�C��?8.����&�;ֵ���\6��'��j�y��(�0�Q���B�"_��,}���1�e��O�|����{���� �0-d�9�� �:�Y���DZ�ſ�;�H�\�����0�P���3�s��}�u;�r�whxS�Y�3s֞����	?�
�g1����3�f�,�2b3��9;�����\�(���KG9�\�)/�R�"�&���v�!��N&kϝ<�#S� x�-�cUx��,����|t��qe$͉K&
;y�����7��P�1TY����_��?�c'��O�V�U-�G�lUf�후1f��7�/;DժcY``���RT	c=�kJ77����?8���LV�M�Uʢ9lu�VL��U��*��('v���+��1c���1<�8@��a��t��m�5E��*j�+K3Ư/�����W�%��"�q��hּ^
{�뛜i_{��sU�R�S�g����ǥ�i�J(����� �,/e��V�S�����!�ݨ�o�
��Sc���4��{&�%�%�뫊�j�Y_�7`��0���~�"�.6X`
f�,�]�av���	��<��N�a)de��%�	]
l�U�N�4-U6Y�W�MNY(a{z�a4��OMƳM�e��_z@es��@!��@&P�8C���IWxkjq����_B�߉���D�u�^$�9�ۄp�*���s�h���ܗ�?0rA����ZWZ�H�"��3SQس)xm�+01�&�VDc�#�t��W)KGY�?Ȝ� ����(��0���ݕ�ȫ�u�|�~�"r��j6`K3Ģ(ט�� I�j�n����d��J>�`��n �B�������A��	ԫY���	/�>�E��7�`x`��Q�<U��VC��g��C�Hd4:~�\�Gjs�g^M�� ��5�����"'�[�y+G+�/P��J�!�xE�q�D���6 3%O�F�3�XW��32;���Sqb�&�W_c��<�hXuEJY,<����y�r�!o5pt��44��x�@�����]A���q�D<x�d�-`���ባg�/R�ѵʂ�>���C�ష��`������5��Mp�s�o�!�L'���(-��5X�)���~����S��*��?g��BqW �鋬����+b�;�w
�fL��czP��a�e(�p�4����h/Nf���K޲�w0���^��p��&��(��U�A�r�HF���D�S��	�v�9s��J3��wbP���cE�y�v��>�f��%*�	��"2bN��L�����hЋyٵ�!&8�S�nyg�$l�y�X�2s��_��*�*Ic�;��O5;PW�ď�
x9\���+�_^�E�3�ك�D߯|DKn��etD�:��j��~��3d�eAe���ɂT��J
�5�,��f�t^�7�sd9�ȥy���J٨��&;Bd�/`_�L�5�\6,�!���"��)��y�3)r\�A	(��ȼe9Hi���Ey�-�>D_��Wd�d�P�@�e╡�RIC��{.e�M֬�l�nW޲n�ˇ�����H(9����iooG?�<�_�#�5+%0ʢ�H��:��t�>��I(���//�'"&��TS����������*?.'�V-Hk���x}'5���y�T/k.]����֟;�h�.?R���^�9ӊ��ͱ�#��=pU+nڸN
�x���8���K���P)����E[[vw�¾�!�9݇�@��a�;�)���f�[,ڮw�z��
`U�Q��-�y��RE���̓�u����&pv?~����GQ][+�b��Ə~�#|㕽��l�06��g>�lٶ�͎O��G��K�����68�,���,ʐ�7"�H�)�סZ'��Hj^ۥ���V͙wfu��ަ
����B�q �PY]�O�٧����'�R��/��ؼ}�T��
1eˮ�x��
���p*PK���wf�)â9r�:::f�s8�L��D�Uu.*�#.2)���ҥ:�������e[��~���}����m؄M7�(eYg�#�͠���ݲ'��&C}���[,�� ��t%�K��`)��w�L;lW&_&��/$/�yn����aF3f3���5d��;;.Q+DGWW��=s��L+��1d����rŋ[0�0�b_	��)
-�z�p��5���bb��9߹�z���D
(3,�~������|��\�@�bL����R�*�%�xAx�	��}���r�̮�S���^8;,E�̂2����|ny�|(��]��(�Y�
����}��$:M������*:�8ݾ�-���a���Lb�G�Q9|���=s(���NI���G҈ݶ�c!Q3�4^�u./){x[3�Ul������q���9���2Q���Uu�g�9��p�����0���C��Ɍ�]���0Sjp,���r�j��H�pr�gNJ����]�]�MF�ۿ��fHYfCAY�u쟿�u|�k_C$���0JUB!��@���Y<���bt|�d��֥��v���B��ٚƛ;�LDG1���$t�E�/�]-XᔭmRN6�Ɛ�ʮ,���-.Zz�պx�i�D�P8.�)�����'�A��q�cޟ/����l���cH�"�C�_�iQ\s�vD�)�ȡONO#�����p��Ĥ�v5����O"�JK�v��6��Dcc#��uT�r~&6�&<K'K��|�Օr���XJɤ`��2�At���|�R�ᩞ��E X�yK�l�[��ZޟX,�JD.N0U� g�Lv򲉒efŽ��Ic����N��鸑��\1���7�����d\��l�_Y�x۶�KE�\Wᒍ@}���p���ۏ��fX[6H�SA���և�SIL��M� �]qU:~v�t+K��$Ō�ON�Z����i:j��睷�q;� :#'Vs��c�Ke���#�d.��ppi?.��1���
`�|L�4��?0S��vz�v�7�R���.r����?C3��&�sr�!��^u�L?.E�C���y"�b1OYj� M�ʾev$�5�%?1��q8���&�����3s��'F�?Ra��:�/�I5_)��G䊆<�,ȩ�OFxH�:k���YE�a$T�X��&d+?�`�Of1_�a���ʏW�$�� |\7���|H������h
Vs�o��B� ���H�^�ұ����z̳�2���j�*�l��A��O��X\�X��YԸR#�Ҙ���S)�x(fy�ym8
)8su���I��Ǣ\N#�b�p�5�>r~H�tr(��8~�"�t�s���#�%A�0�	25�|��'Ϝ�����Y�d�5$���z���35��p�!6̈́#L��S�BOdq�d�
u���ӲAǫ���IL�I}����ǩ˿�t!�T��l*�*��v؛:68[��31���	?A�}�D��s�B��B�{�i�m'�������B:����)\�!�N���#)U��G�@s}O��|.�Օ~1s�x�n��Nj���e�,2��}>��}7R��<�f�U�^����H}I%��x�bw ��I?��*%$ϤS訬㯠h����J&Q$f��6��u���?#�|��[�!�<dl}/�w���b!�a���zq���dR�kJYp���YImy(g!�ǎ�su%�NP8/���-[��_�9��[���If��`�#���Ν;)�Ȣ�p\w�u� SvapP"�M�6!FAƉǱm��9&�5}z|#��c���8z�� �i��_L$O;MG#��b玝b�O�<���fT�z00:�����m�d-_":ݯ�uw�!�������t��:� Y���w/�4����]	"�ljS�}�fю"����mb�y������ۥ�-�=ߴa���		�Ch�J��;�m�v����5�;I�,bf�>�ھMp�RKc��ċ�I�wn�j��֮�܅���ڶM�E��o�qԞ�����͍(^���23$)�?h~X�s�bb�?����#F�,��_.�ʸ��P�V�-E��U�|����/N��Q�C\�����W��)yk�����[�߽�9��h�@4����fJE��YDp�g�]��Sw���n�m�F����a��7!�3d�_揂q���޸~���M�I��)�G�2�_n���"S����,1��d%�³�����1� S���    IEND�B`�PK
     B"BY,��2�� �� /   images/e28c3bbb-5472-4456-9ec9-e60c5bfdece2.png�PNG

   IHDR  �  �   ��ˋ   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���w\������9�=U�nQ8p��{o����,+Ӗ��̲,�Ծ�*��,5-���^�
���կ!p�}��7?��}]OM�����^�
!���?���ۏ~��������n޸B!�B!�%�c ������?~>񏯄��{@,pИ7��Q)@�� U��y��?� {�r	!�B!�B����$��� W�����T0!�#wa)<�@]��?���%�B!�B!,Rp�"� ���%�܅R��f@�?~�G^�!�B!�B!~����V�D�D���0� ���*G!�B!�B� ���g�າqDq'wQTl�&@7�P��&�B!�B!�M^����ce��F
�܁@�-�l!�B!�B!���� l*�FRp�r"o{�RdB!�B!��G�����#��܅!l����+�l!�B!�B!L&��v3�;�le�k"w��r�0�y P�(B!�B!�B���x_
�W8��Rp��Zc����*�B!�B!DIs����j ]�,�BI�]���TP8�B!�B!�����HP8��0Rp�H^˘q���Q�B!�B!��X��z`6pQ�,�BH�]��0苴�B!�B!�BW��6`>�p�0)��``��� �B!�B!�1~��)D(C
�%W�&0P+�E!�B!�B���g`*y��D
�%O5`:0)�!�B!�BQT��&�jq�"�D
�%�'yO�^�"�B!�B!DI��^��"����D�SÁ�@G�@T!�B!�B!�I� c���' �rqDQ���[k����A�B!�B!� \%�`�J�'��,��W� BaNvvv��у�͛���Mzz:W�^����;v�V�tD!�B!��O����M��ӑ�{�"�}�B�G�,BaVժUc���T�R婯�;w��^{��ׯ�9�B!�B��t`� i3S,H����|�S:�B�[PP�W���ã���ׯ�o�6S2!�B!�B'��x?�ta94������@��!������n�:||
�����L���ٲe��	!�B!�:� �&��wY�n�d��u V-��$'''�P��J�����?_*�
'''���@�V����F�!77���d ?~Lbb"< 11�;w�Kbb���\!����ذr�J�4i��}Æ��ѣE�J!�B!�///)W��?�-������������;666��j<<<�j�<z����L����Qo��+!!�[�n��u%�9`pV� B�J�,<�b���ԨQ�:u�P�N*W�L`` �������5KJJ
������Å8{�,�Ν����f�"DI7i�$��� w!�B!��7j׮MHHAAA���־�����������p��9Ξ=�ŋ���6k��o�Ze�}�
w��|U:HQ���%44���p�ׯOݺu�U�JG+�V�%&&���("##��� ""�����	Q,5jԈիW�V���733��M����B!��Druu�q��4mڔ��P�֭K�*U�|eN���\�x��g�r��)�9�ɓ'�{�G`pW� B7Rp�.ϐ�B���AL��Ņ�-[N���	���E�X&��h8�<���G����ܹsG�XBX=///v��E�ҥ㭷�b���&L%�B!����Ϗ֭[ӴiS�5kFݺu��-�/�<y'���<x�8v �<K^�]X8)�[���b�N� �P�reڵkG���i߾�ů^7���hv��Ɏ;���_���T:�VE�R��_Ҷm[��9z�(Æ3Q*!�B!��666����U{iڴ�ů^7�FÙ3g����:u
��Xtd�󀷀\���H���ˁJ1�Z��y��0�nݺ�t$����c~��'6n�Ȏ;HMMU:�oذa̘1��q4M�6%))��PB!�B�0ggg�t�B����С��%�ؿB��űk�.֯_�/���F�Q:��vÀ�JO'w�V�L�A	V�v��>��Ç���t������?�̆ؼy�߅x��U��u�VM2ޛo�ɆL2�B!�B����:t������777�#Y���Dv��͆سg999JG2�5�/�t�_Rp�\=�ow���bŊ<��s�5��+*�*����a��-[��Ç��#�E���gӦM�l�0f���'�B!��Ƙ1c8p ��VW:�w��a�ʕ,[����h��"�S:��')�[������4ײ���u�֌;�޽{��7,��˗��oX�b<P:���6m#F�0�YYY4j�Hv�!�B!,���;�bܸqԯ__�8ņV��ȑ#|��Z��'O�(I_�����C
�ņ�o��Jѕ��//��/��e˖U:N��������Y�p!���J�¬Z�l����Q�L��֤I�رc���B!�BS

bҤI:ggg��k<`�ҥ,^��{��)G�@��A��-�+��U� ��R�
'Nd����f��Ç3w�\v��Y\N�"_>>>�ܹ�R�J��?��&L(���B!��P͛7g�ĉ�����(YYY|���̛7�s��)GWG�^��GP��-�?����@aaa���[����ڲ:�deeq���߿Obb�__			dee���@ff&��� ������
���������J����篯���[��#gϞe޼y�[��8��-��T*�.]J�֭�l�'O�ШQ#k�6(�B!�(f�j5���cʔ)�6&--�[�n���������"--�벲� prr����k�coo����?�.�K��\�r888(�k{�V˞={����匽k�-潢t��L
����R���PfΜI��݋����rrr�r�
gϞ����Cll,qqq��]�*���^�:u��%88����R.^�Ȍ3ظqc��an�=�o��V����/��O?�<B!�B�4*���={2k�,�ԩ�h���tΟ?OTT�/_&66����<[N�R���O`` �*U"00��� �֭K�5���+��u��?2m�4�;�h����J)��஬P��E�'�jժ�̙3�۷�����s����o�q��	����p��ՎJ�VS�R%BBB�W�͚5�Q�F����=KTTӧOg۶m�jFX��ի�e���pزe�'O.�y�B!��ߺt�¬Y�hР���~��	Ǐ���Ü:u���(�_�nq�����U�u�֥aÆ4k֌�u�bkkk�Z��;v0}�tΜ9cֹ��t!�͌03)�+�!��t���������gԨQfk���CDD����ȑ#DDD���c��mj������N˖-i׮f�����W^��ѣf�SSrrrb�֭T�R�,󥤤иqc����2�B!�Bԯ_��?���-[�m�Ǐ��~<ȑ#G8u��~ruu�Q�F4k֌֭[Ӽys����j��]���S�r��m��i�4�7 ۹�L
��hI^�vw�������Ǐg֬Y��}���x<�Ν;ٱc>,�9�`ccChh(ݻw�[�nԯ_��wh�Z6n���ɓ�q�F��%������4Ȭs>�����of�S!�BQ����0m�4^|�E���W���_%33���T���3���t�ޝ�={P�s�����g�����Z�� lU:HI"w��l���o�{�f���E����͛lذ����s������B�
��ߟШQ�"-����1w�\,X �B
�СC����ϻn�:�}�]��+�B!�(x�Wx뭷�|��S�����ٰa111E:���W�d��T�T�H�y�&S�L��+�y�6*�����y�#oe���A��|��|��t�޽��x��k׮e���DDD��"{~�߿?Ç/҃Q�]��رc9p�@��!��ʔ)î]����4��			4k���z
!�B!�_xx8_�5�j�*�9.^���իY�~=׮]+�y�QXXd�С����<?���ƍ�ć`�^� %��ͧ)y��*�O*��1c�0��"y���j9r��~�-�V����:hРcǎeȐ!������V�e���L�4���D��/�1�j5���Gxx�b�����_!�B�������L)O���pqv�����'Yddd����������������pvvfڴi����E�>&33��۷�t�R���'accC�֭;v,�{�.�CW�<y�̙3Y�`��-��� ��R�I��<B�����A�T�fM���k�7on򱓒�X�t)˖-����&�i�ݝ��v���O�\�puq��%�GGG{�ΰ����7�\��'Y ��h���"--���RS3HK��Qr�I)$&���(�&��w�K/�D�ڵM>�ݻwy饗شi����P�?�<��������>��E3!�B��R@B�+Q�Z9*�A�V�t�Vw�'q��m�_���K���-�Ϥ�4�v�ʒ%K�P���Ǿr�
�/fժU<z������Z����_o7|������Y{q̫�8�ak�Woqt���?�992�s ����IFi���e������'<JN#!1�Ĥ�S�0�s��+2z�hƍG�ҥM>����=z4QQQ&�O�.�/
�(֤�^��  ���iĈ|������tܘ�-ZĲe�HKK3�� *�x�S�߇r��������_������\-��S�w�!�����HܝD��{HN=�l޼9S�L�k׮&���a�ƍWl��#88�6��D�����ѪU+Y"�B!����@��`��į�i�ߥ<N��ɫ�?IBb�I�����Ĝ9s�8q���>y�$�~�)k֬)���66j��xQ����})��^��:?(2VN������M"�N"qw��@BbJ�|Vspp`���L�2��-�������5k�%=,K#��ߔR\I��h� e�y��W�XA�.]L:���Ǚ;w.[�n5雽��-˗"�Bi�V.K�j�qq��������~�#�F��z�]�\�#1�I�e���4Ȥ����0|�p>l�1�Ї��۷o/�CltիW/Ν;�t!�Ba�\��ض>����h_$s���r��Uv�p����"�C�aÆ�Y���ի�l���\6o�̼y�L���ўJe�Z�,U+��je�-j�Wff6���}�k1w�v��OL�rI�VӵkW�L�B�f�L6.����9r$�o�6�Fx�"�RI����@U�� t�Ё�����lٲ&����̜9��7��	�J˗�vPE�����6;Kt?��/��ܥ�\�GVV�I�

��7�dȐ!&����hX�`��.���&S]͛7�>}�(�/K�,ᣏ>R:�B!��2*4iX�~=����d�95�\�v�-����)�唤R��8q"������tZ~��g�L�©S�L2����*�S;(�ࠊ���6ɸJ���%�f<�/�����ތ7�
�v����f�� ���?~<k׮5٘F�4n*����{�p��wP��lmm�3g�����ڑ\�x��ӧ���nkkC��iR��Aqws6IFK������8�DEs*�:�S�?@6$$��3gҳgO$�s��a��;wL6��ԩ�/V:�?���о}{�c!�B+�������Y��"�ߏ�����[q	��_ҕ*U�u��Ѷm[���g��M�Ɖ'���ّzu+S�nejT+����
��i\�t�S��9{����-|T�Tt�ޝY�fb��y��^y����L6��́�?����驁���(___֭[G�v�L2^RR�f����?''��7-5A5*�0�*�u+���`�|�"7W˥��9q�*�#�IK�0j�F��h�"�4ib�|<`РA�߿�$�	���e˲s�N<<<����:u�ڵkJ�B!�V�z�r��wwe�egkX�� �E\P4GIS�~}6m�D``�Iƻt����*{��1j''{B�T�a�jԪQ�� `���,"��p��5�_�IN��-�U*Çg�ܹ����$�ɓ'�۷/7n�0�xF:@^Ow�xPH�����Q�~}6o�L@@��cegg��7����o��`���Ҿ4�A�&���t5:Wq���y6�CG�s��-�O�6��NN��s��5z,!�F�V�z�j5j�t��������ϕ�!�B!,\h�ʌ�Ѣz^���)��<b��K��#F��_��d|!S-r�P��iܰ:�vF�*ҟdr��5~�5��w��Ņɓ'3e��?c0!!�A��o�>��2���h�CRp7�	�gJ�=z4�/�����������_����ݯV��R����ԨVu�)����-�<�F\ -ͰU����L�>��_~�$��׬Y��ѣ��0n��6q�D&N��t�|�?ޤ횄B!D�ӬI-Fjm����t�s����݋����/f�رF�����_|��i�x��Ac89�Ӭq-Z�צl/�3gע�r��9N��F�ưU�U�T��O?�K�.F�������_gѢEF�eo��QX��
֫5�P��J�b���L�>��=zĔ)S�������`G�&�h�*o7��$99N����Np�aن���l�26lht��G�ҳgO���K�z����wߙ��ߢҪU+K:A^!�BX���J��ΨՖۦc��l�uT�Ŏ����=�;w6z��W�2v�X~�����pw�e�ڴ}&�ĵ�5V��t>���Q���߿?�/�t��F�Y�l/���Q�L@��(�8���iT N ������+V0d���ڹs'�?�<qqqz����L�֡����t�r�DZ���Q����Ibo�_춵���_�>���Ũ,���t�����B���ɉ;v���aQ�={6˗/W:�B!��0��xmBo�j#�����Б�J�(6ʕ+�Ν;	5j���l.\������������>tnߐ�U,���5���淣�q�)%��}���s��a̘1F�v���0` )))F�c�G@ ��A
�Ƴ#�p�fJ���e�֭4kf\���$ƍ�ƍ����ő6-�ҾU(��Rh7���o�yG7n�_x�Q��W�6z�{BB�z�����F�#J���{���+C''O�d���J�B!���فw'���]�(:���0��ܼ�@�(V�A��ر��e�5�ٳg:t(gϞ��޲e��ܾ!�TG����)�h4��;�#9E��{׮]Y�|9eʔ1*�ɓ'�޽;w��5j#����F@
���*T���z��F���~F��w�GG{:��G�V!8:H��(i�p*��v��w�;;;f͚�o�a������C�\���l޼�jV`���Ҽysi�$�B!�2~tB�TV:�^�<bּ���R�U�Uk׮[�n5j��V���O?e�ԩz��V�׃�ѸAu�<3�8����_���ϧ�n5S�LV�Xato�7nЮ];�]St��:��6%����lÁ���<00����S�Z5���������g���$''�|�J��iXM&��J�ځ������R���7�4��ӕ��u�Snn.���㧟~�u��xyv����- 66���H��%�J�bɒ%F�1'�J�͛7Zy"�B!��zu+ӽS#�c�����KW�|"Ct�ڕ�[����l����4��>�L���vt�А�#:P������Ɔ����2�6� �F<�:�m����ڵk����C����0��ӓ��w�^�߿o�&Px��T k&ߩ����<((����Ǹy�&}���ĉz�W)�����R�q�d�q��3�a�I~>������ެ^�ڨ^4cǎeŊ�!J�>}�0o�<�c����Ì9R�B!�Ba����|s(>�nJG1H�Fì9�q/^���%]���Y�fvvv�q�����Y�JE��5��#ww���x���a�aΞ��뾺u�i�&�V�j��			t�ԉ�'O<�������?�dY�a�=@9%&�]������3�X:    IDATұcG�^���=�.�Ԛ�}[���j���4��l	�Q���J�ފ'Y��=�<y�ڵky��	mڴ1�	�Z��G����p���z/
fcc��ŋ���P:�����Y�z��[>�B!D�ҺE����\ij�GNE^W:��2d�W�6�ؾt�R���Ǐu����/��J�uqp0|na�.N4nP���\��Cff�N�ݿ��+WR�fM������ٙ��믿r��-��0����R"�����a=���N�:���/�.]ڠ��Z-���g�ȑz��7���qݩR�ϠyE�qww�E�Zxz�r�ZM�N�>|�ӧOӹsg�ߨ�R��ر#III;&;E��u�f�����j�\�¥K���"�B!bc�f�Ȏ899(�(e��9~�*ii���0#F�`�ʕ��V6KMMeذa̝;��\�>��ب�ض�Gv���:wRg�~�4oZ��l�7uۭ�����������g�1h����#���z��h"�@i@�Ӄ������ԨQ����S�T)�����`Ĉ|��'hu�?�����ҡ�<Y�`*���
�	�_��;�$&��tߕ+Wزe�;w���۠�;u�ĭ[�8}��A���o���oY�FÞ={��!�B!Ҹau��BՒ�T*T*8w��Q,Z�~�X�j�����7oҦM~������+/� �~u�j�A�gggKpP ի�s���<��龃r��iz��aP_w{{{���Ǐ?�Ƚ{��������JLn����~|�(���U�X�C�`��III��ݛC��|O���1��_���C�l�~���z�{{{�e�Z�liМ���Ç�n�:����3�<���˕�a���T������m�B!�(^&��IP�
J�0���&���^瀕$:t`���88��!**��]��Y�VӡM(=�4��F
��$##���s��5�u�k�.ʗ/oМ<�U�V\�p�����n*1����f�,G�b{�r�8p�������h���u.����2�O^�_)�[!�
�<�ۯ����N�$%%ѡC֮]kМ666�\���ݻt�(���t����R�N�c!�Bxz�P��a�1K���H���JǰHmڴa۶m���G�7o�s���ۍ�&��O�p)�[!GG{�l͸Q�pv���LTTM�4�̙3�Y�T)���K�ʕ��H���r���:��h�A������3����4nܘ˗/�t}9��1�6τ4��������4mTS��3336l}��A���ٱ~�z����_?�J��U�VJ�0��yOB!�(�j�wْ�	2l1_qV�^=�m�f��f _~�%]�v�������2}�`�U�7h>a9�V���	���Y�qqq�j�J��CW�\9��ݫT��6�%&�6Rp׍�'���cÆt����J�HHH�����՘:�eJ{4��<����ڎa[c�C�9�V�믿�ԩS���ё�۷S�zu���K�N��{hi�ի�t!�B����)��jT/~�&c����}�v\]]�����?�mz�j}��3fd'���-,���;S^�K���u�>99�N�:�m�6��R�
�v����٠��4�7�BH�]7�w"�Y}�駴o�ޠ{8@�.]HI)��L�Z��~G��`��exm�Lꋏ�n'�ϝ;�	&�|�������{�n�>$S�F۶m��`2�>�B!�֭Ze�w�-r~��pwS�Pgq���ؽ{��=��Ν�o���ggWG^~���է�m�������a��-����L�ƍ�/,,��+W*qȮ;�'�6Rp/\`��'}�wx����w۶mt�ܙ���B�uvv`���7|Q�T(͛����6��?����Ǔ����\U�Ta���o����ٙ&M�(�dʕ+WlV�!�B������ۢ%k�W�K�����c�ƍ��|�7t�^�߇w�Tl��kV��&���թ�k���<x0�W�6h�~��1g���5R7��[���x�s������_�'nǎ��׏���B���q��	�	�XƐ��
98��$�&�q�^R�ן8q���x�v���Ǌ+��-[�+�X�ƍ�ӧ����V�ٴi�N���B!D�����3��(�HD���ƭJ�P��ŋ4h�A�N�2�����tmP�
��|��
/�����ӕ�U9�&�i^���˶mۨ^�:u���~ӬY3nݺ��ӧ�k�g�@���J
�����6fS�Fv��a���}��ѻwo���K��^�z�SX15�C��R��kq�^��	=zD�N���+$$���$�;fHTa����C�F���aR����֭[J�B!�fP�F���T���|��σ�հa�����w֬Y|��:]۬qcFv�޾�#�xqvv�q��ܸObR���j�Z�n�JPP�k����:v��޽{�s玡q�J^{�]��ZHK��U&�sB777�lق���E���z��EFF��j׬��/���m%�J�;5�o�p�z�-Z���3g4�G}D˖-�WX��� �#�\�rr.�B!DI��P|�8+�v�����W_t�E��>}�N�v���!m����[I�����/��^�ʅ^��h6l�w��{GGG6mڤ�Yzc�z2s�-�L�R���T�:u��:uҩg{�ځ��;;�� �c��89ڳf��By�1cnnn���z�agg�w�}G��{��1q��R���L���S�U�P�f͚Q�fM�T������ڒ��KFF���ܾ}���h._�̑#G�}�*�
///<==IJJ�ѣGJG�Znnnxxx�V�y��!��J˒888���7�h4
%BX{)�7>>>lݺgg� .]��I�&�tm�.���1L�9D�ckkøQ�������b��feeѿ���K�f����B�
�]��N�:���96��OۘkBk!��kt7�S�L�W�^z�w��M�u�S_���xnX{y�*��e�`�Y���BH�<y2*T���z�Q�lY֯_O�֭���1&��R�Մ��ѨQ#prr����+T��8��hHKK�����233���%11����ݻǭ[��~����2����B��w�������C��t�Bݹs��6d�С��Ջ��@�Ƹz�*;w�dժUEҗ1**����?���ݻs��a��Yʖ-K�֭	'<<�J�*��!Ynn.IIIܼy�S�N�o�>~��"+�;99Q�V�"�����5�xM�4�G��hтZ�j�����rrr8�<G����l۶M�]�Jx���<y�?~��Ϗ���+�HaM��(ɚis��-?j��5k���ݻw��/�PM���[��Y�+�?�Z���mqt�c����MOO�gϞ9r����kiծ];�{�=�z�-c��5y�n6礖N�S9�?[�4`�j@������N���)))�hт����Y�1rp�b���Z%����=I��Ȋ���D���^S��m�`[��3V�i��ժ��2�Y��Y������3��}����Jٹ���66�llm�:��Vpqq,����agg[|�g���ʽ��ٷo���z�1s�Lf̘a`B�U�~}�̙C�ʅo�4YYY\�r��/r��Y"""���1jL///�?n���c�ҥ̛7O�V�̙3��X��۷o��H�Rѽ{w�y���L�����Ӽ��{lݺ��{��q�+V|�k�Z�����&���t�ؑ�^{��mۢV뿠 ##����3g�.^,xő�:w�lЖ`C�Z��#F5���-Çg���z�|��k֬��?4w��լY���H�����S
�B]�կƘ���Q$~�����t�z���u>���Ν;G���INN.�:�
FjC�&�yஔ��m��Ԕ�����9��5�k���[[��.�1�����p�!�k�K��[��F�ck�&��R���'Y9����T*ue{{uUGG7�R�..����Zh����C��*W�LDD�K��k���\:t���}��i�h�6r��_d���Ì�v֮]�w�=;;�~���Tl�W���W�]��ć)��^�H�:d�h�c�J�~�:��'z��Ǐ� �i�_����IupRRZ{;�V�.��Ky����)6��B�����5?X���ȠG�=m}��w9p���p�ѰaC�����|�������΅��8�����ݻ9s�ޅ=//������F	�7�|C�V��d�z��y�fN�<ɳ�>˹s�dkP�Z5���+Z�nm�8����1��C��d��N�j�N��	5�8�РA���k�իg��������<��̟?�ٳg���e��qpp`ݺuV����2dd(�^V�22���`V������{z�w���t�Rh�`P�g�]�]��h��%�G�dg�s�p�!4,7r�k�&����쁧���/9ܾ�����������k-_o7��R�R�``��de��[ą�����[�n���/z�@R�լ\����������+�sMh���On�sN�駟�]��0a?��S�����s�ۣV[��S����{�2�d������[3�5�;ǀ4@�_��Ϙa$�T7�<���^������%�$��Y٬���X�޽;ǎ���C���j5�|����:�A�t���|��G���|�r�5j�F�"&&��kײy�f���	ym�#��+
ҹsg���{��܊|�p��	^}�U���"�����ߟ+V�ն�lll�0a�ڵ�[�n\�~��1���>n�8-Z����G���0c�:w�̀�y�	��>���B˕�d=gV�+!��?����ɉ��GGG��KKK�K�.ܺu��k���u�:�F�Z-$$�$'&%�h�&4�k��Wךm��ĉ�e�W��� ?g�X��1wG8��.Uʳ����~�!-�J��&++�c'�x��������Ǻu����\�r|��W���Ϙ��zX$�sRK%�z�5�d�{�����������K�z]P�
�{��U�lOz��~�^�/�6��}����y�n��Y���������%ǧ����֧�����>�x�Y0���l�Vp��+W�0l�0�mۦ�6�J�*�x�b���[����� ��R�J���ۼ��+�\��+V��8;�x������(y����ڵk��������?��R�J1s�L�ͫ�^x��?���v�լY���Z�jŅ�:*�5{�}�]f͚e�q7n̩S�h߾}��=P�w�y�1cƘ}^!D���A2����-�t��?T:��,X���sUƏOddd��u�FǶ��f�Z-��?|����������l0�Ǩ�M��4��/^�g���ܩeJ{���v7�
3R�U<7�YYٜ9[�o�w�}GÆy�����o߾<��s�X���p���ĳΊ`��$o[�Yz!�.]�.����}Ǐ�E�dffx]y�x��U�<����{����YY�i�-ݱW�<�x�>Y�ٳ��{���t����o��}��ŬY�x��w��_�~lڴɐh�~�jժJ�0�Ǐ��'��z��|W|��_�Y���l�,�����p�ȑ#:���j����r��9n޼Ijj*��y佼�pss#  �z�����s�	&����|��YS��}��aÆB�퉉��߿���(HII��ח�e���3���m�kN�ܹCÆ�{��AY]]]INN6[�Ɛ�'NdѢE�^����O?�ĉ'���#;;����B�.]
������<���K/�ĢE�
�s"=܅����P�����Z��Io-#=��Bqо}{~��G����'L�4���5����m���G�i��$�rvr�:��ה�c�I/�l��Q}P�T������y�����G��{���lmm�駟�n]���Jpp07n�0"�^ҁ*@���@
���,@�������;��=���4lؐ������p��W���i]�$�<�s����j��'O^e��
�jQM�}���������XS��V˒�{8s6����j5;v�K�.z���=jժ�Çֹ���Ã'N���q��9�N�ʥK��󚧧''N�P U�9r$���CnԨQz��oNNNL�>=��gΜɓ'���O�?.�]���#QQQT�V���:ĪU�ؼy3III:�_�|y�¨Q��Y�f��feeѢE�;���g-��� Ξ=[`˞��Hf͚�֭[<s�L�2L�<�����������i�Ơ������~�o��U�V�۷��̝;�E���w���&L��w������ܼy����BwG��o��ܹs�N
�B}ؚ�ᵕ�aR��xo�wJ�(r���DEEQ�J��;r��[�.�<���8��Uu�j�V܃�ɏ���)�p��3��AU�w�v!�m�2^�K����'d�?a��x�Xp��ҥKs��Iʗ/���{��ѻ^c�E��s/�Jf��|�[��n�ɺu�Ǝ;��'77�N�:ڷ�����/��B9�u�1ڭ�⒒�X�l�r�
�Ng�"Gwm`�d��J`�ƶ��V񽗕�Â�6{3��뼽�9s�N�A�nٲeV����ߟC�,�ˑ�edd0c�6n����N�<�WkТE�W�
����,�a����Y�M�2�9s�?(..��^z�-[�<�Z�楗^�>ȷ�	p��)����.[K�}ǎt��-��.\�o���Y���l޼�J�*�{͘1cX�l�^Y!o��vh�ZBCCIMM�{̂���_���ruu������w8�<�z���5���{��|��Y��aÆ�4�!lmmY�`/���N�K�]�����3���1L��ٰ��/$Y�p�N���.>>�����+x�n��y]�����@�FCll�������X�ǟ0��w�+�/`-����?d�ǛHK/�]~ӦM9t�P��5�m�С�]�֘��� ���5�%��?zEn.f�1���ιs��.L~��G����^�R�?�!��p�$�n'��'$O��=�+�Ŝ&�ԫ
*�7������X��`JJ:�/��G�o:hѢ��F�]\Z�����[e�Μ9Sl�ǚ5k�9s�?
}[�l�N�?4�O��鄄��-�4aa6�Ppwvv&..OOϧ�~��ڵk��![��[�.�����7��#F�`ժUz�k�&M����o��f�>
���GDD���O}����T�Z��V~��t�ҧ>P�~����fΜɴi��}����K�.:������{��~�����޽;;w��kL]xyy��w�ѡC��B.Ύ�o��V׭"_}����┎Q��������iϞ=] ����[���;��w�B���Z���윬a�~���y�i<���P�T��Ytq��m>�b{�h�O�Ό3�;!!�Z�j���#�e	0�\�Y"���Rt���5��ٳ�.�GFF���oz]׎�����QrdT���W��������O���p�N𵘻�,�~������uƶ�����̛7O��U*K�,���xK��h8p�@�� C�e��x�~��y�^dd���?���7�b��Ǐ�ر�Ɋ� QQQt�Ё���W�躺�ڼ��K���~�z�Z���޽{t��-߂z����ٳ����w`�ɓ'�˔���
\�w��m�u�w��Z���7��1�f�2y�V�Z�W�]!����A��X�c�L���\�~G�E��Ύ�˗�UlX�dI��v�ZŘ����s���Wn��h�ВVlX���=����ҩ��~��?LT:OajT+O�M�����׻u���/}�����?��9'�4Rp����h�Phh(�ƍ�람��^�ʪZ5*Эc#c��'O25���^R�n����w����m�}��Ή�k=��M��7�ʁ~�Ӣ��M�������ժU+t�����믥��nݺ�p�¿����[o�{����3fzފ!N�>��ٳ�}�A��z����+}��y�k������kF��?�O?�4����x���?�5��ÇϷ�F�a���$$$<~lll�~�իg�Ë�qqqa����۷O�,Ba�#��{n��:z�r��3a��w�^�x�ɓ'z]�nM�Y]�����Q��衳n��ٗ�O+�Gi_�ؽ��֔:y���G�i7�WX���hX��ݐ��M��Ç��T:w    IDATe˖��Ӈ=0�\�Y��^pw &�k�O>�D�'�S�N��ٳ^S�ǝ��vB����$Z-\�z;2���r?�:~���7X-�^����ז:{>vqFF��X�L�`�6*�ྜ�F���a�S�N�\9�{�y��٧�//��t��W���ѣ���G�Q:��0���O����,V�\Yd�Ν;�����:u*���жm�|wA�^��۷M���?�w��3�<��X5j�ȷݘ���lذ��~���9֬YCt��\=z�����ۗ�/���x�ka�	!�>Ξ�%�E���Iv���\_�v������zݓ���СCIOO/��!U�����,AVv��t�����f�,Y��l���J���o��J��*u=��~K��:rp[�����֭[z�O �c��<����P��C��昨��z`����Y�xq���ب�l'����Wd��f���>r�⭡��m�f��P��~�t�K/ߨu�V|��y�3�+��|���˗y�����ť�U���> .�x�?������ڵ+���DFF*�$�޽���%~a��ʔ)��׮\�Bbb�} ���,����͛��Jhܸq���{ }A�޽ˉ'�����o�탞&�]Z��S�N�������o[��h4�|��ھ}{��� ��V�Z�믿�q��BW�/_���>�̠y��i�Z-?�S�=�T~�8OrJ�gsY���{/��?�����������#��R�u�A��KwC�,�3T9�oƌ5)smn{:*�_B�e~388�1�َ���`w�ʕ���z�ݠAF�iL<}���5��)�w�9&rtt��CLVV�����h
~��޹�K��\��{�ƽ�_����Y�Œ?\�`���g���eee[�#W{{[F��Ph?�����]T6l͚53&�"RSS�:uj�Z�m�J��ￏ���v�*�9rssIHH ;;�H����;wzp�(Y
*�� ������Z�Z��|~s��ד��k�]/]ʿ]������ԫW�?]���A����4���>����ӫW/��[�t)(�RNN/��2�G����[!�(̱�W�gx�-�=y���p���U��޻��^�Z�1�JųC���doL�"���ў�xc��KP�%˶G)��Z|�b�&G�'��_���?˗+�C��O�Q�w�ƍ#55U��gϞ��������`g��,II.�wj�c�I�&��=�g�.���jU��Զ�ɊƓ'Y����ߚ�hS�%���dižX�{���7���?LV:˿U,_��]�_qyxǍW���S�T,X�����CDD+V�P:��pssc����ٳ�����Hz��A�&Mhٲe��z��͕�A�?
z��g%��������y�k���V�>��������Ç�=��P������ߎ����S�ek�/^�w��!�0�W��Ӝ-[�,��B#���w�qQ\���?�K�H�WT�J�X�1v��K�`I��5Q����5��b��Q� "�{����_�ӄ��awgv��~��?�ݹǰ;�g�=G�®��v�ͱ����e/�b�V�\	��U*���K�%Q{v@���W5-=����]V�?�Ihh(��iҤCE+���WLܷ��zw*�S{_�4��:'!!s���u]777L�>]�����_���	�;��	bGGG|����^���C,\��u���>�U�궧���%���ak�q?:����W�/X���WW���(��H�u�����x���v�͛7�r�JL�4��u[�n�>}��رc�SPK�.E�-дiS�C��ڵC�p��5�i���:�o��ȑ#�������q����ٳ��a|�9sϟ?W;O"�����k׆��;ao�~����<���!))���L�ĶK�q�ư���ӄ���"8p ������@zz:��ӑ�����H�R^<�ٮ]�P�zuxxx���U�V�����Ҵ��N>�}M�W�^�q�ʕ+Z]K�R�ѣG�\k޼�V�*++�O?�����{����S;~9���5.Fw��Ν;�K�.�^�y�f��kVwE�-5	M'�^�>����^�-<W�X��-�C��(����w7���tH"F|��K�!/���Я���O>����X&L�ʕ+Y{Ci�D ��XH�Tք{m ���4y�d޻�&N����S�ށp�b�IhZ����ii�[��Ď�XL�t�@����Zݸa��Օr�D"�gC;c��(--�% ���b�С�Z�{���'N�0�eee		����acc#v8za���X�~�V��O#���B�[������o*�
�֭+wL*��Y�fD˖-�����$�Mjj*bccq�����_�s���DxYYYHMM-�A���F��5k��4��Ç����b�����3333��$`KHgffr�F�j����T��	wƱ������߬Q�F���FA��eSϟ?�I�&M�B�a8�{��rGu/���>),,��g�T��|��~���3X��d�Id2�)�T��(q��'*mml]X�����БϞ�DխSUoJI��ZaH��ش��V�B����~�?����IW+++L�6!!��En	��!��s��h�wwrr	x�����j�ԫ�v�M4	M�T* �A©E�7���lׁ5O~s/����R��B�8١OO��2yyy��7����_�~��&���D̚5K�0􆍍:v순�+#-_��1!��ݼ��Oi��5k��åK���~L�0�[��P�x{��s�Θ4iv�څ7n`�ƍ2d\]��?y��ի�c���C�z���r)--e-�R��挥N�J%��.��6L�z��E�_�� 2�6������Ç~��� J�B'�+�q�i���ZJ��w�AF�qo��ٳ'ڵk��5s��Ez:{M��]�Y���b(-+Sݹ?�������_�4��}�U�JG�hV�Mj�ιz�*�����cǎ����&��������	w�%w�ԩ�������}��SS>�Yo:c�
܍��iՆ�$������5�abPvN>��u��j��nݺ7o�04w�\H��y{:y�$:$vz�y��05լGJRR8�8������_X�d�?��A�X�b"""0v�X^�6����@�Ν1�|DEE����=z4�U����Hű}ΫT��s��U�V5G׮]O'���r>yp����fffh۶-�M��M�6��ѣ8{�,��ñc�̞=~��֚Z��x*.�~���q�ӳbupo߾��Ç�������B4�&=��?���2�Ca�R�\��	b��s|w�?z�k׮e�Sս
zv՛����+���O�~K�/b�b�Vm<9�NL�l�\�79��;��i�ԩSy� ���P{�C����.5e�-����L�;������_�zͪU�����9uo7W�7d�B.�����l��-aSŎ��ؼ��ń�o|22���ۍT*�gC:�&ǕJ%&O��뺍5!C4O4���óg��CoXYYi��;v�������Ǐ5Z���Ν���l���`�ܹ8q�z����e��.[3}�t\�p'N����~�av��Q�2իWǥK��k�.�l�u?�����:w���p����[�"++�/_ƢE���_�o߾�ҥz���>����éS����=z�w]�c{hP�J�����|����h߾=�g��+;G1N/�`ݖ0���_�]��B��b��s}�����֔)SX�_H$���;��D?J�fe�>y��j���ab�RY��6�~l�Ȓ�R�H�Wq�A�^�Y�$''㧟~�u�ѣG�F�ƬZ� `��ʘp�R�E���[^I�����R]��Э�~��,-+SݍM�i���b�R٬��$)=�ћ��(�S�������?p��	^ם6m��c�������:�1Xٔ�����W;�ŋZ[s߾}C�N��aÆ�ŉooo�ԩS������???������B��㏬s�R)��k׮���ۘ>}:5j$P�����ۣcǎ����s��Ėp���ƹs�p��M�5�������۷/Ξ=�˗/W�97۱y]��b;	�����ZK�,��˗5�B����X��(�����R�®�q�B�(�<m�4^�/_��S�N��iռ����>MN�3s��<{�q[����*��[�w�{�ط��D/��wl�/�G˖-Cjj*�k���a�ĉ��ƕ �X}!~AX^ ��z+++�;��k�-[��!׀�m��	kY�\u'���[�7�Ke�fMX«̌���t��a+XY��Ι9s&�i>>>�ڵ��������j��._��X�]���ZY��ÇX�x1�O���7��SԨQcƌ��Ç���P
�� 6l@X��F���X�p!bcc����[�����Xeann��x[����뜮eoo�Z�ʯ�ٽ{wܽ{AAA��om۶�͛71i�$��Ǵ}
�����ތ�ԣ�bL^$���G���^\���X�����g; �h�mڴ��u=���Lѯw�&aiMFf^��T�-���;��j����c$�Շ~zR��>f�UPPP�ŋ��_|''Az��Y#R��C�<1r�H8;;s������+W��iP��Mkk���
�=H޼#b�رTvk׆�N{��$=#W��26��݃��zLL�=��|K�蛽{�����b�a�.^��i^^��Ϟrrr�`�l߾�G�6���nnn>|8v�܉k׮aɒ%

��9�C0�9�R��Ç�n�Y�^=�7��ׯ�5k�P^�g�f=u0o�<�����e�oi���o���X�l�l�ί���a��A��}���'�*�h�B�՛�l,��.]��z->x��~ޏGO��	@S��n�?���uN�.��`o�IXZ��[P�����[�DP�R�m�u�D���!�P^�a}/���7P]�~=�������1f�MC���[eK���R��~�-��������e�.�H0���ۺ�T*�W̋�6l_%v,䭕O$�ſj��T;�����#�~���.�nݺ1�73f����y��&�
v�؁+V��_?JwU������6�ƍX�jz�����h.++]�vը�E�F���W_�����֮]������]�ђw}��ǘ>}:���s�p��1���߫Q�Fa�����n݂B�(w,00�uG:_#G�dgk�J!���L�=/��_� �U�`���b��sX��r�ߋ%�Z�j�o߾�^��?��Wq�E�����/��=Kܰ5�ر��6n?}�^l�X���ߥ�4�o[���l...ƢE�x]388X���	��>�L	�� ��z�޽{�aC�'$��Ұz�j�9-ꫭ�$����7m_*v�}�w�{��ir��"q�8�dR��يuNll,<��!!!��%���\���@.����IOO���B������?~<��I����
={��/����ׯc���4h�N�#Vv����ܹ3-Z��Ϻ��7Ə����#%%�n�9sФI-DK��%~v��Ÿ;//_}��kru��]����gϞ�_�>������v��a�ر8r���;Æ����9�����+W��;&�J1c���U�����:��c�,.?�| ;��Ǜ4�=,O~A1~?u��F�G��KHH�r�'O�ĵk�X�������O��BY�\��IҐu;��R?�i���M1�_�����l�Z�o�ؼy3^�|���nnn2d���q� ����2%��y} �_�֬Y����q�T�����9�Z%�_�9�R580$�v���WLܗb?m�/O����ŋ���/Ԑ!C>	z�����/b�apbcc9ϵ����gݺu�V�A����cǎX�p!����w�^�9�w�B�L.�cƌ���ǹs�z�f͚a�ܹ�����k�0j�(^�D��6l���0���J�¨Q����S^��������ԩ���0w�\�>}O�>Err2=z���(lܸ@�5�x�b��V�6m�0l���޽{s��T�6�M�Pb�J%�\}�9�`��pܽ�B;���ǧ`�����agn��X��΂����g�}��5?��븋�=ڴ���R���/�n�qD�@�u����0��H��;�á��R����m�����`�SeK��T�Z�ХK�󋋋�~�z�9mZ4��+{�]{��楃[3��^YIl�snkL��7��I$P����ݻ�p��k���cذa��&�M�6!**J�0ʣG�8ϥ���d2�l��f�¥K�p��Q�?u��;4�p��}t��-Z��Ν;��_�]-[��֭[��u^)��ԫW�������K���~�s���Xk�+
L�:mڴ�ܛ"++ӧOG�6mX�J�R�]�fffj��s�N�2��;w�Ԩ�̬Y�85<����B�R���ϱf�)|7{+��>�?�=DzsI���/��ϱ��%��q��8�KW�L���!C��������7o�-�׻GK�d��b�ؿn��E���jÉ���S�����5�6f��q�Fdgs?eӲeK�J$V��2�%�^��q�=��AԿ�ر�����2�uo���*,3;�$;#�ehh����z붆��,���1�6���]Y�,[���5ǎ�IHzA�Tbʔ)HKK;����+�s�V���H��D"���&O����DDD`	�Q��ء��7obĈpwwǐ!C�c��~�Zkׯ_�><�#G����Ek�5f�������YOvDFFV��J�F��r���O?�ī����ݻ�V�Z!..�qN�����矫�V^^�.e�����+W��s�μb�H$X�x1�Ν�i~II	��B�1�/(����}o$f�ۉo�߀�?����ر7�����G��k�l�vKV���1y�����c���#�_C/|�%���?�̞�vwsDˀ����������x��4�4x�Җi�9��*гK �̘w����aӦM�����I-� @���TY��$����Dm��w�T*��;Z4�g';#���2��I\r���ô�! �g^�:5K�[*y�H���ل���*���֭[k�������w�U(�R�I�׭[W��Tu����	�Ç���T�DC���8p��?%|���0u�TDFFj%�د_?ܾ}�uw5y[�'**
^^^�s�\���?��Bu�
�lق���#>>��k�����~�P�{��5���"�9'N��@uٲex��㸣�#"""�v�Z�����^@@ .^���S����r���%�	!())CbRn�}�+����p��\��ŭ;��<>�b��w���ѦM����;�=��R�W f���S�S\�J"3K6�y�ڭ��T�����>h�~2q�ʕ(-�^v��O?������q�_�E�TY�=u���~OOO��#""���C�9];���ރ[��8{F� oK��)x��{I�x7~?��pu�gW�TX�j�k�3FӰ����y�zYYY�晛��~}qw�#???,Y��N���o��k�s*�
w���O?��.]����	ݻwǢE�]ᆫ^^^��?дiS-Gl:w�.�Օ��Օ+Wгg�
� ����_|��� Ԯ]����]�6ڵk��k�V4��ܹs��Aj���ѲeK��),,ħ�~�������ǏG||<N�8���ǣk׮hҤ	��Ga��鈎�����Ѿ}��\�~`l|]\L	$B!����ڵkYǲ��B�f�}���x�4iȺu��}�!zc��3>x�R�@];��>,JNN�ѣG9_�������!�"b�	w; �VЈ#x�Ww��Q�j�����.�LJOZ��45I5P;�EF�>LZ'��R�A�t���cm�o�������_~�����a�=�; 6lH��u�N�:ؽ{7�7����)((��3g0c����=z���ŋy�#���������IG���",,vv�'���O�����刏�GTT�V땯Y�99���6=�z�*�����YZZ�W�^X�v-Μ9���ܼy'O��Ѻu�r�)<x�/f,�C	wB!abb�O>�^u���۷og������;u)�a���/- ����§>�Ky,���Nv���:�oY��+� s�G#Pl��    IDAT�] ��r[[[���}}jj*N�8�:G����%���t�ɰ���u|B*s�5l�k+����\<x���lll��j#4�)
����&M�MII	nܸ�C�a���8y�$�߿�X.@���m׮��b oYZZb�ҥ�`C������ӧ�Y�f�Y�&&L��K�.qz}�Z��z�jGi8�O����ܜq�.������{�2������k�.�3F�e�~��7|��P*���233��&!���!((�W�cǎ�͛7���f�h�{�I]z�*=�ū姢@�"� �Cn^�h]��uf��?����u�ԉSYAI t��"b�	w����ӧ���۶mCY�g����V�Fh��a⊭[�1w�"##3�{qq�(���LѶ{Ma�OZ2�f���ɘ9s��apr��yt��C�����1k�,����o߾���ǠA��r�J^��samm�i^���.)��������RIHH��U�бcG4m��V�����kj���̰}�v,\�����ɓ'ѭ[7���
��.\��8�����Z�7oF�^�8��b�T*�`�8����J��'RRR4^�BH������Z4`�$�Kr�\����/44�|�͛#S?O�!���k��fu�҉*�
۶m�|=�L�~�t�
0�2�!�� ���J�-[X�l=�t"�eګM;#&��:Ѷ���<z�(a�X�l��^�������9_�W�^��������سg��a�***Bpp0����W(�}�6V�Z�=z���<ȫ1[[[�s<==����*{"WL1118p z����t�y�'N02���䄳gϪ-��a���ۗWi3}q��e�1'''N��w��������p�����]�v�5k�?;�mmm�-7�mK!��ajj��}�r����H�9����~���#;���- �U���/}��\��۶a/o۶�W�(�6;v ^='3��{ ^�\���ݻw�<��?�d�j"��u������2^�f�O�ŉά�zzL��LQj��8ۣ~�f»w��|=+++���KӰ�����#��`������"��ccc1c�t���6m�\��<ի�?�3`� ƄѾ�5k�B�w��i�k׎�!���S)cV�n]DGG����o*�
�f�¸q�P(�N{RSSYOJV�R��5���1p�@�h��w��� B�P��ŋ0` |}}���7^�F���wB!|u�֍׿q�w�f-�V��ս���Ѧ���B�ԓ{1zb^geXRZ*Ji��`n�\M;%%E��w�o�:/�������g):�z�޽{����C�����ֆ��8�!=}�u�ٛ�,NtF"��Eb�X-�l�E]Y�C���Q7`� MC�+%%%��R͚5y�������%K��[�n8y�d�֮W�븅�\�k������-yߣG����3����W��mڴAtt4�}���#G�Ă�L�T*ktM�ߺu�~�)\\\ХKL�67nġC�p��l߾�-������N�:�ȑ#�&4�N%$$T8FB!�S���y�W�{sw{|���7n��7э�;#�<|�tT��-��Т��g>=��R)�%�y�V,ƞp��|�8*�J��W?h͞�ԕ��"y���x
d��l�y�i\�(����օ�s�6..7or�ӭ[7������?�y��F�,,,4:N�������3��aQyZ�n�:>l�0��2ת#���ghl1~�x̙3�V����q��%<x� �-4��'O"::�q�y��F#����#22��Όsrss��Ga�ΝF�;l����5�~QQ"##�d��;�0j�(̘1�Fjj*�5������J�B�E"��G�Ղ=z����q33�����x�OH}�yי_EY��\*�43;_����VM>��~�U��O�S:�ۊ������2�]�v�<?**
��Ɍ�v�VhXO�p=~��}˖��R��ee��˅?>oj*��:�s�<i���3ʝ��'��\����Z��F�8�<>��CDEq/SX�n]ԩS�{�jժ�ꫯ4����֬�2pvv�ڵk1w�\|��78p ڷoooo�h�B�x�vni��5�&M���Ywu'%%�]�v8w�閣�#�XFF���0c��~�޽
׊'�R9�����������>�j���LӰxS*UHNJc>�H�ƍ'
�ǥ�c�Z5���T~�z ����ٳg9_�s�����(F��6ʿ��S@5].ТE899q��nw{�_H��wK��)(�P�+��DP[v�������b��ܿ.�8߲2={��4$�4{�l�������U�Vi��mvv6F��k�iyIu333,_�����C�y��1�?.v�b�� ��έ�P�}���X�lk�۷o�U�V�w�閉�	�����@/J�YXX�U��Kr޽{W�h!�:>����d�}?Օgq)�v�h<; H�<k���&-G}C-�H��^����D�v�4K ���1cN���XߤߩS�XǛ���[ҕ��_mݾ�X�ŉ���
>-+�ޙZ[��{��&HHH`M��_�E~~>���y����6lؠqo�B�y��a��͜����C����;99a�ƍ��&�����0~�x�m2�-������вeKA�a++�IW]Z�d	&N��:����h߾=^�z��X���жm[���cǎ��ٳ�믿b߾}�ݿ��N�:�H�ߠ�����WAAA���)w���U	!�u��^����8nnf�&��{�R�BnNᗂ/L��Ox�L����O�:��L��ʽ�b�	�KX:���!�8ngg�:��?���SP�]h7Y���(��|��l�W����\W*��ϧ6.G3����M�r����/<<<t�D�����`�̝;W�P�#00�w��W_}�q-�ŋ���Ym#�D����cРAHOOG�V�`mm�����O�<��W����+���B.����666���G�5РAx{{C&�i���JHH�_|���D�C�����裏�>|���D�����!���P|����sV�\�ɓ'�hȐ!X�����������z�۷g�S��](.����{�\.GDD���!�b���vzWxx8븯O-��	��iܫ'w���?���l�y6t���\��u^��]ս\���7i�厧����͛�7
����&M�f��	�^׋͘�:-�lgg��� ������|j�RN�y|��C�N��vZ�3Y�*����q��ה=�~��iL�:�ӵ$	:t�}��i+<��g��h��z�;������ѣG�7nht�ٳg����j�R;���&qqq�x�"._��{��!''��kѳgO�7�ah"##1e�����޸r�
c�}ذa�3g�`�n�~<$�M�:?���J�BHH~�U�^dl'�t�s�S�N�c���k��� ���������pqq�����vr���}��)w,::��!�R�v���*��%�.���\n_v�Q�H���ԝ.��c�^�ϧΜ��q<<<�s½aÆ�Z�*RRR�^yt�S,�ZR�@c].кuk^;����x����T���M|a"���#/?�-�VՆ�<aj���ҕ+Wx%A?��(����6mn���ZnnnسgfΜ�Q����"�\�R���/??�w�F�޽ѭ[7,\��/_��>���,�ݻݺu�4MC
�.]�q��Q��_�zN���a�����ajj�aÆ1�cَ�#Gb��Ō�
��F�4��'ܫW��kW�:����ׯ_�c
�B�=�aÆ���/ѻwo�n�ժU������K��5b�������V� �Ryr�\RR��/2�K�4���V�Jx�&m����_��Jba>)/�P���O��u=>��
����k½ s].�g�Raa!._��8n"��a}Om���Ӹ���7G2w�#F+5-�9c�#��&�_�ywpYYΟ?��zƞp/..Ƙ1c���s�C)�T*ŨQ�p����Ӈ���:���())�jl���شi:v���P<|�P+�-..Ɣ)S��6vRR������jf\Y<{�����1c�`�С:�#88�������O��<!`ݺu�㥥�<x0v��!`To����6e���ϵ�Vpp0�������W���֭[�����	��>LLL0mڴr����m�6�� �R��I�]�|�����j���Z��T��*}����m�x��y|��;��֩
ss�I7n�@FF��	�{� ���"B3ք�����v�k]̺u����La񒕙*��D/l�sn}fV�v��4���:~��%����񁽽�=}Ovv6F����$�Ca����˗��ѣ�ٳ'�Z�
����s6O�<A�~��d�dg�_�N999�>N'�'N�w����/�#�X�|9�D"������'��l��m���d߲e������%����x�F�Tb���8r����;w�d1b�ׯ��~~~		ag�#���ׯ3ֵ=zt�c�۸q�P�v�rǶmۦ��=!��gjj��͛s����d5�Gu!?�Ha�d.��7���W*���d"��a=/�q�B���@�)�n ����2��s�#�m�6�
�O~������0�&zA"��Eb��]��9ڤ��.��CC���+<Xow���I�&X�jΝ;ǫֹ��k�G><x��C��ѣGZ�^y���P����Pu��� �}�&N�H%d88v�k�l333�޽�V��J��w���aaa���7o�`���Z]Sl���cMXO�:�0��ڳg�ry�cfffX�f�F͗mmm��~Ɵ{tt4�/No޼��s���ڵ+k}xu�5k��~��ܱ��B,[����&�R95k�VVV��ͽ�P����חW�
|��;���WbR���%ԕ��{�����9� J�ͺ�Ѹqc^;k��Q��RfCW�^eP�J���d���"�]ak�ܤ�Ν;(((�|=j����T:���Mg�E�j�0e�\�x�BHH�����<4�6m�ʺr����:�=iff��Ԕ�x�!�w���郣G���A	f=�&�H��7������ꫯˀpU�vm�޽���;lmm煆��C�z��!88�q�ĉX�t�������ذa�x�.]�f͚
��ruuEdd$4hP�xII	���K��ۺu+���������;ƦM�",,����?�|$&
�>�B����E.�������榨���8�+9Y�s_�蕔��]B�Y�NU�q>	w�'M*H�y\1po�lXt������<W�T��ի�㦦&�^�Eaq�P(QPV�|�T
;�]����Y�˥�PkJ$@��Uq'&���I����W�գ�Fff&��իWD�z�T
���EEE(--�J�����V׻w����z�w9::b����ߞ+�R��7bŊ�;s	�;w� 88�5�
 ���X�f�ϟ�����㈊�Bnn��5\]]ѵkW8�z�R�C����j��w�ތI^mz��~���>b���g|ȥR�p���3F�� Ο?�gϞ�Ι9s&���ww�r�ǎWWW�=YYY��m۶-�mۆ�u�2Ι;w.�����;�<yR���#,,���Crr2��:�ׯ���]�㱱����BH��ɽ�ۼU��;�Ra����f��>|����T&��ee��LM+���<ܝ`me����7ݺu��Ō�'���Ϗ�����m-w�i"f�	w �Ŋ��I�k<x����fuW�hpĸ"_����񅠋����V��e��k֭͜p�>i�p��1�SG�������cڴi5j����fiiɸ�QSl;~5!�JѫW/L�6Mk�o�Ajj*�L����h�C1h7nD�ƍ1a��s1v�X�;
�O�>���ϑ�����(�JH�R899���4@�Z�8��O?�J�R���{&O���k��z�j�	�5j������H$�7o�.C������&�srr��������;�?��c|��X�|9�n݊����̑�d����1d��]�.\��?����RZZ�o��gΜ)w�e˖�{�.-Z�M�6��pH&�!((��=�������D�~�PZZ�+FB!��}O]e�:�� �K�)��_����/f�L��X���`5�$�vM7�<H(w����n�⼡L�܋�� �� c½�NMZ�gW�[�X�Ÿ�N�:%��D/��.P�T�+rĽ���f?�ħYc�ڵacc�ډ��(
,X� ׮]âE����(vHz�^�z6l��٣��YZZ�W�^5j�V��s��a���w�v!!!())�w�}��52�6DÆ��ӧO���t�\O_�=Z���b8|�0,X�Y�f1�quu��ŋ�p�Bܻw�=Bzz:lmm���N�bbbЯ_�
�P9{�,�l���(���	K�.ŢE�p��<�YYY���D�5ЬY���
����R0 O�<�!�bbb�F�q���m��:�ؿ��B^~1����hed��Wǃ�-�S�*c�x��ѣ�;�6�K	w=�};X5mʽbMLL�x��&�U*��X�J�E��ڷ�⣆�<�U�j��^.0�� W(��w��kI�R4n�׮]�Vx�ܹs�w�~��t��]�p�Bhh(|}}�z��
�
vpp@�v�бcG��F��� ����h�"�=� o�T*|���x��	V�X��&��DFFb���x�����
�gϞb�P!�gφ��	�M��:O*����~~~�׸v�z����슆�q������{�f�cjj���@�=S���1`� \�p���B��4h�����=R"j�p�FX�ed��;tQ}GsR)�eʕJ��;�T�͎u����+�դIH�R���-GM]^\hƘp��ˋ����͍��Z�����M;ޤ��=t񎠋���&�VU�*�Z��Dw7$��(w<..������M�6��	w�m�㯿�;v�̙3y��0F����C�~��?��Ϟ=Cbb"������hccxxx�jժ�_�>|||P�f�
544�?FHH�>}*v(Fk��͸t�֭[�ZbC[�����?b�ҥ���Wh֬��aT�������c�^�Z�a�lق��`^M��#��1x�`�ر�Rto�7�1>|��kB�|�lt�����Tq����f��z���=�I��Ν�kVu���p�jM/5�F>	wkkkԮ][m�E���Ņf�	w��D�s�	`[X���c��t%55���aR)��� X� �<��J����hժ�ky{{k34�t��E\�|�1���xy鴍�Ahܸ17n,v�S�Tؽ{7/^�����1zO�>E�.]ЩS'̙3:t��C���"l۶���Cjj�V��O�V�*xc3m۾};����\��z���z�?Ɣ)Sp��I-D�VQQ�Q�Fa�ʕ��(,,��t�R��B���{O�>Eqq��!���I!񒛛��������s��ù�P�Y[Y����9�oҸ��?}������u�ݨv�7�����giZZRRRǽ<� �f�ܼ�0aW$��Yᴻ���WM����ϓ�ʾ��o
��FPPƎ��/�W�]ff&Ǝ��s�R�K`.\@�N�P�vm̜9���5���刊���_|���F�l`4�)���лwo�j�
;w�D^^�׫T*\�xÇG�&M��l׶m�P�fM̘1��w��$&&bΜ9�[�.,X@�B!Z��{����BWP�T����	�(�{%��&[�%??���%@��1�p��;�f͚��>~��u\觬* /+���=�:T4����j^.B��Y���ϧ���de�P(���HT�R;vD�N����ww�4qDEE���Ǜ7o�E'�����ϋ/�p�B,\�h޼9�6m�5j�f͚�Z�*���`ccSSS�T*dgg#//qqqx��)�ݻ�?��Cg͡k�����
���?�g�����q��u�=���h׮�7o�*U����	U�T��矒��'O���͛����s����E������?ڶm�V�Z���NNN���F^^233���Kܸq����믿���̙31s�L�� �RAZͽ����mo�r
�o�h|v�FT&�{�
�Z�L�5�<�����ٓ'OP�NN� �ϣ�-    IDATbT�)�1�^]���D�ŋ������J��-�{$*N�E�A��ʋ���­=�Tug���SV������~�����4����ׯWWW����S'���eee��˃��+кuk88��Lii)�={�7o���������Z�IYY�/_�͛7C�R�yGqq1���E��*3�\�7n�ƍb���b$�b��|�KHH`ww6����C������[�kh���S�k��.o�.r/ L��z!![���N߸|��{�:;	[�==#'I�����/� X�������5�����=������Wvv6�_��ޟ����y���С:t�����G��m�6�9s��
�1~��g��m����1q�Dܿ_�P!�B�0333xxxp��>�"X~ ��[HO�I�����<�|�ZϹ
�{_��R N ��t��%�u^�K�OY���p��/~ ��`�)�g Lj=�T
Gdd�;�g�;��sI	w~�5k�!C��{����z)))X�`"""��y}��Q4-Z��t���b���|SEm9|�0�͛���B�C!�B!D#իW��{>[�����fZ����RE���QPXr�p	w5}����3�$�nl�
��H$�j �{�{Ҥm�E�W]�9�.���	Z��Ɵ��Ϋ�����6B2z�={�DXX<�~��	�l߳gz��ӧO��9��t���&L���/|}}1y�d^O�Mnn.&L��iӦQ��B!�>��
^�|�8�,�FG�R3�tQb0
�/	����d2��/������?eiuH؆:D	w���ajj�y~rr2㘵�,,�}�Z*��tAb0:����4[��I+���ߜ��枬38|�0V�Z�����faa!&L��~�j�s�9�رaaaP((**±c�лwo>|X!��7o�w��;B!�B��J�*�禦�����䳓��r�K�o��-��`(�RA���]]�IR����^�&�cl	w���qv�w���4�1��*}�\��R�~W�E�A��/�&��=�g ==���~6+sssL�6��탯�`'א���pNK�R4i�D�S�N��ϊ��0m�4�^��w��H�P��_Űa�x=�"�B!����p���{�K�Q�r˯�J�C�.�.,*)������^222XO��� ��I�[w�>	��$G�T";�������6B�,'���СC
A%���� /�ֳV���p������РAA�}��F���iy@@ \]]�΋��c[�bLLL0n�8�����L�2���ءB!��|�ߩ��(t�%��䍠���SPdei.�.\��KYYrssaoo��Z�Ý;c�����Q�yceeeA�`�o[[{���/�^�TJ�%�̙L�Q�����|-J��W�f�p�����/_��'�|��h�ȑ#9͓���˗/�ٳgy�m�J%��݋޽{S��B!�5>���}o:�RR\�\P� �łV���d�{`���$w�-���.Ґ6o��j���V\\F5��2�R�_�%ܩ�Lŵm��v��Aě7o0b��y�oS���7�u��i��%��S�Tbʔ)���͝;w0`� ̙3��B!��ǧ���܋���	w����#R��e
��6s/����ꐱ%�uڅ�ښ����L�Ϗ�r�VZ&�tAbp�rA1P�� +��C_>�Mc׶m[�_���悮[ZZ�q��!11���R)BCC!�H8ͯQ���9����T
ZO�^�x�ɓ'c����w���B!�"�u��}o:������ 18eerA��>|r/|>�$l"C��-���Vqq1븙�������ψ�JI%�L����MY��}�޿��ܓ5ҤI�[��?�?~���C�E@@ ��u���4�ƍطo�x����D�Tm{��!���ѽ{w;v�WB!�B�6s/j�wj�R��{51<�
�-�Z`�&��'�bf��}� %���N�|n������&2M��E.�SI�J�P	Z��D�g@�g�]������;6nܨ��.�={{����:oooL�>��kZ�n�y�+����7�����#))	,����y�2\.Ǚ3g0z�h����N�b�B!�B���������u\&6�%/SR�T�J!��p75aO�������[�]�?���M�+�"A$�G��r9u	w>7�ʾ�����W������k����~��:{{{�Y���n�6m�p�����u����?�6m�ɓ'�����ԩSq��U�K֔�����˘5k��W_�ҥK���B!�Tj����{��)�<A$G�6?'3aO����(@��hvS
[�D�t���pW{��)�B�䞽$�R�R)h��T�C'J�s7q�D�������x7I�����P�zu��yyy���w���4Ϟ=7n���y��.̘1ݻw�ԩSq��888�U�Vhժ|||P�zu�&2r�			x��)?~�7n��ݻ(*�g��B!��K����Ri����T*usl���mv4��%��\��M����u\&�SV �~��ᱴ,4��)�����V�����_��vvv6v����5������_Ѽy�
������s½��{������+�޻p��	,Z�{��EDD"""�����'�ncc������ '��VB!�V�j�wj��BA$G�T	�QW�Z�r/F��1��2:���9�/�H�]L�h�Q�T���&Zg&�S 5���[V������,���J�N�8���8,--�a�t��Y�u���ëV�޽{�����ļy�0o�<���^aa!^�|��/_��ÇHLL�d;!�B!<h3�"t�FI�D�ݕİH�RA�#J%��@�r/F��4�����H@.6A(�J�J&��B!�r=���!$�'�|>��dԨQ�S��h뇇�s���䄝;w�}�������A�q�����7nh��}��'غu�(�j	!�B1V��q��{�����X	� 18&R��_ )�"J������ڄ�B؛�D*5�cD7T*�p/���F0v�XQcx��1�y���8~�8�������SSS��O�<�����u��	ѭ�B!��JA��a7;JM��p'�$�=B	wqPmv��)�L
kA$�T"Ӭ�$O
5����믿����h�T*�?���0a��ݻnnnZ]����}���QQQZ]�]m۶�ʕ+E+�C!�B�1�nuas/R��A����J$�&��<t�y�2�^*��<h�)��ǚLL�]��DZ]����p�f�c���aÆ��D"A�ƍǂ��p��	L�0��Nt>���k8::r����K$%%�$ �ڵ+���+�]�B!��� 7;�ʼ]�S����is�{e˽h��<s�km;���X�7���IA$G*��r��"�π������)���%L~��GԮ]�������Ç�رcذa�������a֬Y��?y�D�� �~�-u�!�B!Ǝ��;u��ν�$ROA$����Y�����?O�{��0$999��:9�o(/(����33S�jO� 3�z�^��π�3�����5�`��ڢ��b� hذ!Μ9����d288z���Μ9����s���u�L&âE�УG��v!�B!��f�%�@���ML�U]�SS�c�ZB�q�w2228�U���8�niaFu�+s��B���>7���tM�1�R{�FhNNN�$���`�ԬYS���|����鉐���C!�B�����N��F�7;��VtAbp,-��@�̈́;��heG	w���mll`aa�8.�M���J�2tD��r��|�π��
�L7�����qpp����akk�:O�R	�ȑ#Q�V-A�"�B!����~�~����++s*)CX��X����͎U�p��W�͎���;|�zloZ��5��X��h#�ĠXY��	�^A!=e����u��;�T�n]�ڵ�u�}������d��oY�B!�c�������^��,��M�J����.�Z�����������UYr/�@	w���\\\ǲ��!�fK �D"��R�p+Cco+�S�̬<�qJ���G}$vz�I�&صkW��u�i�F�Xz���^CYB!�B7�L�ge뾬��i�#a4�_ۦff¶��d��ɻ @ff���T�p硰�������,-�#/������Դ���ѷoG�*���>eM��e��d���~��k����A�y{{�رc1b�?e�$	&M���U��_$��0l�0��#�B!�X���q�����wz&�F/m����ؑ�%�r����R_V&G^s�F����R�*�fGm��;O/_��<W]��o��V�-]�S�R�D�5�3��033�|���Dm���5j$XICgkk�ٳg#::���ǅ0f����ׯ��y�B!� ))��|��azF��� @"��N)R.+K�@!�S����{,55%%%Z��r��;O/^��<W]m��.��Y�tAb0,MM;	�^i�������J��	��={������E������%��ݺuemB!�BիW�P\̽�)��ǲ2�X���tAb0lm,��\O�	>����xMéT(���7��%�]]m�I����pŭ�vw;�SVu��w�~��W�'Cս{w�Cй�\a�B�%�B!���wS���^��l]�g�jB�����:�'�B	w~(�����%�[����R:|@z�J���پ���%�b��y���3i�4hP)p޼yS���]�vTV�B!��9����(hR����w�bǽv�$��79�p��m��;O|�`6�L&cW�t�Sӡ�/J��g�Twv��rMu��F�q�Vex�ZYvI_�zU�����-ZP�B!�B���{��f��!t�����䓁�h�;y�D��B�����:�'�B	w~(��S\\繖���[��9��7Y����3G{� A$zOf�/%a���aФI����4T=z�;�+))��;w�C'ڶm+v�B!���ϟs�۴iS��$6;Z��>|Q�����R�^3�pwww�����U�܋6Q���X(�J���n�
��S��g^NuT*�]%z��޺��k&�b~�jii����������FHz�^�z��ŵk��Ag|||��B!��r��}�s===����8.FuG[��5Exqw��}g�dd梸��q��ח���=��m�p穰�Ϟ=�<_]�%1)MӐx����}6��ǂ.J��GU��B�WXX��,�Nٍ�{��T���Ez�JST슽`AG�QlXб�gg}콏��G,��D����Ny��՟Rn��g�Y���S������OC���*S����Ldd$���Z�Hn\]]!�]$�B!��dqqq��˽##S�3hu�ck�Е-�I��3�kGSc}��o+����a���HOO�6�
%�%�$�'jkӛ�Ti�aLWW�O��4fDW/#���:)<���L>�KJJ���+D��~�r2�j'����`kk��0!�B�1޽{��L�>~O�s��ď҆Ĉ���ڛ�1r��(--��S��<�R�Lv��/(�.&	wQ��%���> Զ1�$�I�R�3Й'�9�|z�M�6b�������I��rrrbT^��z��)��������$19��B!�"����D�/v46ԛ*�I�R��6�k�v@t����]�bcc�燣�ٍj�dk����������bD%>sC�Qû����(;[��Sԇ~����ɨ�cǎ ���I����St�B!��(Lr/��#�� ��,�SY�;�k3k+SCy���!��֦��hР���z�:P�]111������7Ii҆Ę���|�OJ����a&��Z򜳌�ER��_hԨ���=|�Pa)���Laa!BCC ���
���XZZ*:B!�Bj�������������%���zz�ԓ��M��D�h�i/���^I)�(�r�o׮�s�T=�R(�.����}�V���۷z�ūw҆Ę��ez��c35��M�s&&���\�]�v�L�y�,�RJ���puuUt�.((����ϟ��R�YXX(:B!�Bj�[�n1j/l�cy9�^������l�OJ��]ms�o]."�رcG�����œ'O��C	w	EEE��V�֦'�R��1#vR�>�PÆ�0tt�h*�y�%�Ϥ�LAA�J��V�gggc���߾NOOGVV�#�>�����B!���իWHM����ŎOD<�V'���{Ց��D)����573Ԗ����Lr/QQQ�
Y-O�F	w	1y����&tu����̖�b+sC���L���6��Z�Zr��$�C���C��ܹ����	�͛7�y������^�����B!���Ν;b��<�T�	wu�k�����D)�,����HJ\�ZWWW�!��c�ӄ|A	w	1��SSSCϞ=��QěVG{�:c�u	Q�v���37�o�>���ؘ�)٪��_�vm4n�X�aT��w��СC|�=z��h��M�!�Ba��s_�&M`cc#�~���ΑEX��s�B%}<cFt���h-�ɤ2��y
��y�w��ZZ��ʥ|�%�%���8��^����'�Y,�M6�}b�PF��nia�+�y?KO�g>z���()ɤ�SMӻwoF��4yyyX�`�����EDD�? 9���Pt�B!��8L�,K�N��'IRFĜ���fJ���OL����n�Ϩ�Q�|���p8����6��a�PYY"""���%V{OOO���U�`���*)�@KK�I���l��zwu�,"I����2�C�>�}-����R�+..ƍ7�Ii1���i�\.f͚����Wy�ѣG��ʂ����#�^jj�~���tuuѼys8;;����p8(,,ć���k��Ƣ��PѡB!D�DGG#;;FFFb��ݻ7ޏ�}�.r?�v��~@I�ĸa}̝��t���e\.�Ⓞ����{���(HՏ��R�p��	w333�j�
��ݫ�>�S���D�iY_�!����f�� �E���s���u�(PM
K���[��Y,���ׯ�lR���M�4Qt�f�ʕ���x����ܹs���cT�O�w,(R�N����
�BBB0g��D*000���F�	www���JKKq��?~G�Avv��"%�B��*++CXX�"V��={��f<�+��Gd���P���m�M'��9s�+Te��m��W����W]=y��¢��]\\���$�x/^�EX?$Zr'�.0j?p�@���?L�&��Է�4fDw�f��B�Z�lPļ�^�Lȩ����Bk�U��g�&Q�r2�v��K�V�СC�	�?T��ߩ������ɩ������f��p�B$%%a�֭�С�X%�455ѹsgl۶���X�l����1!�B�������v�*�>��C�#��^��-���@*n����m�m=FD^qРA��S��Ku������K�ۏ1Bh����d��"4F454X�&��>1�+ߟ{N��cn���E}�>��x�����J��d�ƍX�f�Xm_�~-p7PME%eȏ�������'Ui(,Y���ьV�B!D�\�x�тQϗ�Z�heal���k�B&'r���>�SKK������a�{IMME\\��a��( %&o{���ТE��9��޴6p�m;j�Gg�LN�]@@�����x�N��-�����g�Xbo���$<�\�)KKK4o�\�a����ҥK�u�VF�6lP�fB�tuuq��5t��A`���R$%%��ӧx��	RRRPZ*x�A�ƍq��J�B!?�w��!>>^��C�������o�>���Y�Ƙ��Ւ3�h)drR�&��j�ҠvwE��$Q�"����Y�fb�w����y.O�p�ҹs��1b���7n?�&����agkrX!��j�>)j�����"掺�\�a� о}{��ى=ӟ�����ʪ"++�Ǐ����?Z�߿�۷oWCT��J���i�&4m�YBB.\777�������5B�ƍaoo}}}�l���Wq    IDAT�'>|���������B�	!��ژ<���C�}�u�,�b���@�S�ڧ��I�31�;������A7���ϴ��*�^�2 R���@zz���&��̛�T���!��sr��=atϙ
��T���[�֯3Qs�x��;�_"1������	I��飐2o�"::^^^�u��c,_�\�aG5�p'��E�7n���kעq��X�z5�����.--Ń�t�R���`�>�g��͛c����;!�B���@Qϙ7�>�+xaXurmP{�رu29�6��z��s�qV�ܟ3r�V ��^���~��(�.���2�:uJ���ҥ��67D$(�S�����N�+y�U�t���/���RW��/^��UOSS#G�{�>H��Uf���BKN����X�fF����4��z�����d�bQ��3f���X�~=�ϟ��������Ä	�wo����А:VB!��<�=³g�J6l������-Dܓ$D�\-mM5K#c�f�� __m�z�;��w��S��_Z�l	777��EQQ�,B�aQ�]��i�4i���w����T1�:��45���ɉ̍�c��sm�t���(�u�sss��;~����45Y�^������"2s��U����v��˕ɘ6l@RR�L�R$*)CT�ł��W�k�>}��ŋ%���a�̙x��m�떖��ݻ��qB!�f��������o�_^��9Y;O��@a�J�H?enj������rD��2JT�2U�, /������*k�
2d����	�_XX�["~X��k}���?��� �L��hԠ��E�a���Ã�7B�L�Ȭҍ*����O�Ab���5j�L����d��]TT�Y�f����t\y��D�թS�����/���X�1���c���]�v�xLB!��l�^���E
>�fJ�T\�Y���i�� �LLݽwc{�Շ�~�
�9�תUK�y�������˗e���2P^^��'O��^KK�G���J�C��+�4`55\�������B!�P�cE��+����GBW�;99	=Ȧ���dܽ{W�)SSS�j�J�a0���#L�6C�Ž{��m���x�Z���ƗJ�Ufjj�w����R�[UɾF�I5���6�ԩ�֭[�C�pvv���|����A���ѩS'������R�sXXX�iӦ�ڵ+Z�h;;;����|��,--Ѹqct��͚5���m�n[�vmt��	M�4�C�򃉏�Ǔ'������;�4i"�>�\	$��$b���a�gpCa�͞=����M0�����WE|{{{���H��N�>-���[�����@̘1C���&M¦M��X����G�ߠESŜ�ab��ii�@�"ODi�����mSE�_\\��"N}�8q"�2���Z��&�ٳg�)'��pp���۷>�ۼ���GÆ1x�`��)K�pW;v쨐`�{�.֭[�h�iӦUX�]PP�w਎��o���;S����f��粵�������������������R����+�~�EEE���@FF�D�;&&&���E߾}ѩS'�$-��Ãp��9"%%E챵���Κ���Eaa!�/	��ӧc���_�>_���D���`��݌��~�b���ၟ�����kS^^���X\�zǏGLL�y�ץK����[�nU�WXX���p�?AAA((�⪲=z������<����? @�Ν�v�Z�nݺ�\�O��ڵk���&�B�'00���^~~~B^�{��u��A�����޲������/�VH D:���������[���$����[�c߾}҄D�?U� ���lLtt4�U�}���ŋޯ�h�����"4���j#}��,Fy�iҤ��Z�4���R���x_GG)))U���Jyy9���d^�DY�޽��jy�r�����ٳgq��E��>�:ijjb����ر�B��ǏѩS'E��r<==��=t�|||�mΔ�ԩS���'O��СC��o�>���~�:;;����O�:۷o�p���]�vō�C��������޽{��N�!���BGG999`��oGaa!����ܓ5MMM̜9����ثz����y�f,_�yyy"�����322BNN����f�����{����9s�^Q������۷�=���BHH.\��/_���r�ֶm����.v���T���_عs�Xg�L�<;w�����s�Я_?xzz�̙3��֮��˅���LvVBQn���x��=�����]XX;;;dddl�S�Vط��Bd���Ë�K����k
�06i��V͝�)rmզ��x�L�b�6m�0����K���(r�c�n��\�����ٳ�Q��s�
��:�#��|'MHRk��4s��^���������l/)�ܖ7q�D�����Z���l���B�v����r���`����ԩF���Ǐ+,� ����:u*�����h�;��Ν;q���
���԰w�^ԪUKd��s��%ۓ����!Jaa!�ܹSᚎ����_����t.q��ŋX�z5�-����X�`�_���_�v-v��%V� �l6�N��3gΈ�@h۶-n޼�(�|�,8p �����;w.���%����
۶mCpp�ĥm���,0� ׯ_�d;!�� 222p�������`���Bۄ߈CA��Jhhjj�Ե>?e
���)����ؤ�}�"�S����𝙋-b4�?�������2t���VC}գG4o�\h�3���_��luV��6�����Sh D$,S}�]+c�� ��c��
�����_~��ј���a)��mۊ�8����;vĈ#��~���+:�o���0i�$<~�Xѡ0¤|!_�x<L�0��g������о-Z�����+\+++��?����,�Ǻ{�n�k:t��'O0g�FIoi�ƍ�֍qLvv6N�:����c�ʕ8p� �����5k��oߖ(�>s�L�E��ň����˗q��}�//===1o�<��#88��eFQQ�]���b͚5X�r%��݋�ϟ�a``�'N@___���U�Va�ڵU�f������v�Z�ر���(++�k7h� ����H����E��?p� �q	!��\L;���/B_����5Ŗ&31��6�1�@Jnܸ>����4�����;�wrrB��������~��!�A����|?~�Q�ٳ�Wky������]�kd��i[�2v�����ʈ�̚�������"c()��J�����Fݺ�M����s��I�����"p�\ܺu���;ڶm��I�����1nܸU��V�I���U�"}���hӦM�}tttp��a��ҥKq�֭j��ȑ#|�܁/+�׭[���4���a��hڴi��L�X,�q������`ƌ���Đ!C0w�\���o������#z��ɗ������Ç���dɒo�;!!>>>011A�6m���֭[���~~~U��X�p��D��ŋakk[�ڶm�`ii��ݻc̘1X�`~��7L�8����ӧ_yKKK���~��;w�m۶�_�>Ǝ����cڴi�������o�.�[�O�֭�k�.��U֩S'���O߾~���oߎ�K����HMME~~>N�<�h\B!5۵kא�� v{KKK�9Rh���X��I�T�-r�^UhD���a�����(t�\�x"bu�ܹs���y����2�e�F�/������(�M�w����kKc#5�f�mUN���Z���N�W���J�#���%��b1�Ҵs�Np8iCSZNNNr������͛X�x1ڶm��c��رc��̔{,���Ά���]�e)�N�q��Y�D���:���[�������ťµ���o�OV.��#F,����	�Z�
�=����q���7N���~~~8�b%������c�֭(--���իWѪU+DFFV�޵kW̚5�Q_lBBBмys:tEE�m,**={����WSV__�{��rl6��1c�T���ӧ�ey��Exxx�`Z����c�ƍ|���ߏ�;
����'�����ۛ��{���5j��9+344���W�\	WWW�����?����/лwo���=&!������a�֭��̟?_h򱤔�K�ds��4\���?ы�~"79�8���6����'�.�������e�iB"�P�T����p���/$544��m��6���64�99X9�~z)�%��I��f4oZ�WE��r�
qY�����E�b�YXX�m۶I�R�d{�$���p��u���pww���/�?^-�%䥨�S�N����H�p'Қ;w.�!��7��ŋ+\0` _����t����uh�4RRRйsgܿ_d[kkk�3���x��5RRR�1c�H\~��f��_�p������Ë/D�/((���޼yS��ܹs�|�!L\\F�)2��ի
+⿪� ԩS��������ŋ|R_x̝;��0�+W�`���|�׫��ӧ�]������ڳg~��7�~III��� ������F�\]]E�r����҆&5�F�'������ ͚���k���'4����x�J�y����+�ҵ��Ѹ~������P½�[��Q�1cƠA�B���BI��W��ԯ�q�~�):�Ÿ�{�n��q��v��p��W�r��p\�t)�1��߯�U�-����H,Z�m۶����q��	dggWۜ���r�l�2̜9�o�2��DZ=z4ߎ�E����K51KKK��+���رc���G�ę���:`ѢE�>k�ԩ�oeBN�>�!C�0��2d���+\۴i����#??��%���5��������vA�*�bgW��9��� �:d����`�������X�v-�N�Ze�|�����1~�xF;9��ك˗/W����
///���p8"�, ���)((`\�}�ҥ`���s8e��64��������/��}�m�#�fꄟ6t���8��r�8}Sh�*KR
�f�i�"U�@5�t�bcc�n���.r�{Vv�������}���Q�L�4�sx���A�
_:�����>�f���hڴ��c���W��]Մ���t<����p,\�m۶ń	�RI���?ĳg¿�V�Y����K<jjjbǎ`�Xسg_Bvݺu�x�<�Dii)V�Z[[[�7QQ�\���0p��o�aA��+1bD�����%�{��I�CM�8UTT�S�N��>--o߾�p����*�a�l��<�^LL�5k���c���عsg�/c:u�SS�
�N�<�w��������1����D�BQ}�7oX.�*����رc���y��W�����7uu54kd�~��^~���G�?�kO37�ъ���#5]�.�%K�0Zݞ���ӧOK���Մi�p�ȑ||Uv�j2���'����gMpE�q��&��Ӥ��1E�����S7��xc�ٌW������+ŗR�n�/_F||�Tc����ڵk�?>���1iҤ*F�.11C�������J�YY�r%_	�.]� 44����p�޽{����^���ؿ?:t� �7G�e�s�q�Ƹz�*�/_.���b�C�����H������ƍ�U[���XF� ��*a���|����5OOO����s��2�MӱcG�kǎ�h�˗/����ҥ������!�������������Î����r�?O��lV�&uwMׇ�s"�L�w�Ic����8WPX�󗢅�qttd\�}Æ(++�&4RJ�W�Ç�� FMMMd���)ÿ"���SC�:=�����=?�q�g�h�_KS9��w�_�\0y��o%�U���).���ӧ�%PD)))AXX�Νwww���������U|�AE*))��e�0u�T�Z�O	w"+\.>>>|?�Kt���`�ȑJs��Ǐ��~�5
���hժ�Ν�s�Ή|9����ŋ]�^�^=XXXT�&͎��O�V���ʊ�\� �k틣�ߧ�D@yyy���;w���H���"((���011a�WU-�w�Dc�x<DGW|8�W��
zA<P�v�B����-��"_��ۋ<���ψ�%ݢ(Ya�����a��q}�}!�j�~��ڏR�G��3�PPX,�͚5k�=�����{�J�%ܫ	�����ͨO���Eִ|���O�W7�����;��y>����G0mR���ݜֳ�l����/(Ɖ3�_#  �ѸgΜ����&z��������k��
q�ҥoI�ɓ'#$$yyʱ�E�\�z����K�(
%܉,%&&b�̙B�L�<�ыy*//GLL֯_�~�����mڴ���˅��������d���'�߿/��F�����F����.��"^�gƺu�� 377����=���tܺu�/F�-}U.M���.ՙ#U��V~A"����B!D:/_�d��}��Ű���������~������Ѣi�es�Vt,????�9�F7r��Iѱ|�"�=��	_LұcG<�Ѹ+W�Daa�4�(�^�8�/^0�q�F�ۛ�G����V���hoYO��M�8�OmEǢ�x<����Ь��luu���=~���
�l�2����=&��c��W����߿?V�X���Xdee!==���G`` ƌ��-[���!!!��W�_���Ǐ1z�hlٲ�Ѫ��@��Yۿ?���~���p��q9G$9.����h���pss����_�^e�իWCOO��zU5�---ѲeK���]��WAu�+������Lxyy�|��������c��刉���w�~�z�h�B��W�gffJse����^��B	`TC__˗/ڦ��G���22�a� ��Cf���������1����Qn��s�V�����2�aUS�V�`���Ç�&�@5�r��믿��[�.�������)����U����Ĵ�����{�
��_?�_�Mp�o�[ѱ|�ɳܽ/�����+�L��h�'N0:tX���� 00C�A�֭Ѿ}{x{{cŊ���R��5	��ŦM���ヴ�4��A+�Iu8q�D��k�����pt������;����Ç��#n2\��!�|/_����֮]+��z̞=111�u�Z�n-�m�d���SU�;300�/�`&�"JBB��������o! �=IB�C�:W̵~�6O����,^�;"6�1�;Z�'ձ5��A��^��O����7i�$�lْѸ�����/�$���{5;v�_PQ�.]Z�ʪ�]�����҄&s��:�n��L��w��cQ�|zvq�2Nqr�rRt,�+,*����B۰X,l۶b���r�l�2i�#�Ͻ{����k׮)d~J����������6m��ެY�УG��D�Z�d6ֺu��w����w��c���b������ƨQ�p��Y�շ}���s��=�Kܰ�l�b�����XxRB!������ѡ�jjjزe�Յ/?z"9����*/6֦���F�&��fV?����kQ�Fv��Lt��^'~ĕ�GBۘ���ܱQYRRR��g١�{5�r�X�h�>عs��6<t����a��Vg5i�8{�/�͚5�H���d�~^[[5�nfj �셌<��,��&L��nݺ1700��*Bĕ���ɓ'c���~�eK�ّ$ѫ�+��'{�쁕�U��X,���/ա������͛7���K��塰�NN�{G��ʽI�&|�*Y����%��:$��_�TTT��G����055E�=�z�j������}OMM���O�/g*�q144�*ƪ�S�PB!������۷3�����ӧm�_P���Ä��P}��n�'gL�=lHh�<ݹ3�n٬�JmmM��s,..�ރWP^^.�݆����c �g�%����ٳ�x�"�>}���r���rrt4L�ЪM��6M���R'����Xj��S�l��д�����r���[w�"�Q��6VVVX�z5�q���d	�N�������1l�0$&&�m^J��.&�x�����ĉ1p��
�>}�T�k[[[�رC�y�Q�vmt������j��i�Ff�{�>|�p��	U������Y5EII	��°p�B4k����?~<���QRR�מ�fW��u忒�    IDAT?OKKK�+ ��������G��#�B��l�2�߉DY�b���O�� ,R�ʞ���pk���ǂ�M�_O���4����4�a�5�g�V׎������|��ݻ7~��gF�޾}G��&4"J��ɜ9s�_޶m�ȷT�'���xiB�6&FzZ-���5�X@�0���i
���J��cQWѱT%�S6���!���͛'����O���J!�<y���c��2��:*�����d<�4	�z��aÆ����]�v����p}���3f��s�#!��l�Νe:G��U�"�� �f͚�4����Ǐطo�;;;lݺ��M����J�|���׺��hР��qT>�����޽�x<B!�*��ٌq���`Ϟ="Ȝ>�w2�	����6���l�bڤ�kh��h�ڳ�m��x���@�����^�K�qf����m��h\��Y�f	�Id�2 r���3�ڵ�Q333���?}�o�%�Z�������G-����):e�˔���7<����R]]m�<q������PR"��ѐ!C0l�0Fc'$$`���҄Gc�������1cƌj?d�V���ʫ�������\]]%���f����|s.X� �_�Ƅ	���nٲ�'��(�Cܽ�����/�񵴴�V�%'�a���k��=z���e���;z��hkkK4Fu��Ѐ���.]���/==3f�@hh(߽�Ʒn��k#�SSS���U����c�ۣ	!�I�ٳ�?f�������B�p8\����"�,áSKK�Yc�yK�|?mR?��������&���ХN?�������L�g���U��r<x� �ݻ'ih�J��Q@@@�5F�=z4������p�ر����tac#=��M���c���i~�:*:e0Loִ�]����ձP��GND�|�okk��� ̛7����p�\��P�]uU���N�:���m�V�E/^��m�V���s����X�bE��

���0Ϟ=Ó'O*\366F@@�L�����+�SU� nܨ�����8���p��a\�pϞ=CQQ>|� SSS�c�ZTT


���3�<y���+�1Μ9�w��¢��7o��k3a��s_~���w���	!��>.��ٳg3�i�&ԭ+|�y��l�=xY�W׶1�vs�so����3f�1Wt<�b����ۼI�Cf&�Ju0���KJ�s�E���'���3;??_���d(�.GX�`�~;w���6�Yy�t����� ulͬ�Ծ1{���3��C5������w���Af�u���W��{�"cq��s�m���p���	����#$$D���Zbb"�͛7W˪K�%ň�z��}��mmm���(vQ��qww���^�Z^^&N�X�oŊ���Xc�S�NX�p�D󊣪��g���ɓ���ʪ�m�jN8p��ڒ%K��3f���ׯ����m�iii��ݺu�K��R����;%���Q�Z�V�Я_?Fsb޼y|׏?�hB!����0>|�Q}}};vL��<qO�����҄W�����R�N'��f��ݹy�-EǤ(���=m���l�99Z5Q�uP<���U|L�P���{��e���?��;�TJ��Y`` �^�ʨ���!:$ru��oq��mi��:\��bgg�2kꀋ��RtL������'��_vjin�F����j1?mO�^$�ǉ���͝;ݻwg4vnn.�L�"ih��TYY6oތ�������2���
I�Ty'����O�.V_///�j��������`���/X� III�q8�7��%O@@ Z�l�xnq�޽���:���Ν;�k�.1�����ᰱ��p��իx��A�}.\����ӴiSlܸQ�y���<Dt���b�Q�Ξ=[�kMMM���b�g�X|;'�����3]�nߵ]�v��{DMM;v��k��M���B��̜9�(�Z��[�P�����I���ɏ��ۭ������铼6�����Y���A����?S���k�:��}�# �w9���%����޽{ae�,��-[�Ha��r���0u�T2�ױcG���o"�]
{�����)�����KO{'��g��`��V�����Z0^��>;�<��k��q����r� 5-;��.W���V�Za����_�h�F��͛7���UeIIQ�]~������$������|�fΜ��C�
���ba	����������\����d*{��!V�ZUᚆ�:��-))����QVV�w���o޼��+ШQ#�㨫��]�v

£G����R�~QQ��-�<�-���=u�T�ݻWd)GGG\�t	��w_?|�PiVd=z�o���ɓ�`��V9���_h׮]�k'N��;���-22��5kkkܼy��&{e���8r�F�Y�:���̙3E�I!�H+##s��e�o���"�H��xص�"��$O�t5�4v�Y�Q^0wƠ��:LeK������������yzCW���5"�y�aB/���_~a����`�ĉ�r���G$��ox:	`���ǂ��E)//���.\� ����f�y���R��S^�C������U�6-j�iZ3���+��,:���R�9��+��'�9#Wh;ܿ�QI �s�:t�@���������K]��͛7�ի��"#_yzz��ŋ�2vNNN�+��l6���ѠA�
�y<N�8����˗��ͅ��ڵk�ɓ'Wh��}�j���all\eૹ���777�������BLL_�{����=�kڴiغu����Ǐ���S���"==<fff���@۶m����x���EPP��8֭[�9s��]OII�ڵk��� _^������ƬY����[�OAA����������w����������{W�\A�=�}/0�=y�d�ܹ�����ױe����WH��S�N�5k<<<*�),,������lll���C��5�w�������r[[[<.���-�x��ͫr弰�o6ĳg��!�B�	e��LKKC�V�D.32�Ţ9�`b�'���))�'����p�o�q6Rt���5ݯ�h=]�_�,]��kD���W�?`����	O��k���%����b��P �):Y������lܾ}���8233ѪU+$&&
m����3����4a*LNnA����/j�i��n��hE��į�3��\�����hk����)��-�E��WWWǥK���)..F�-����[�Ɔo��^xx8&M�$è���;�4Lhh�D��FGGcҤIx��ѷk��VVV����[q=m�4�رC�\�[�FTTT�R4<^^^U�ԗ����c����Ғ]�P��)S� 00P��

z�|aa!���`ddėd����ÇGhh��q�pg�X8y�$$p���l������@�˜��r�=Z`M��ڶm���P��ï������'
�A�b�
,^�X�\�p'�"k����������~�o�F׮]QZZ*����)�mmfIPe������9瘮�ڊ�[CkT����qxKlm����ʨ��ҳ��(((����111���f4����Ѽys_�D@E�5뵏
)++�ȑ#���+���	N�>-rKxqI)6�<��O�҄�0��Z�]�4h`s��?|r~��������x���h��Q��~���>Drs��f�g��d{������b�
��v �?>=<�#::^^^�x�����`%�̹s�����x�Ntt4���'VY9����@�$�kת\�,h���׋5���M�6�w�LƋ��G��N�_��F�B@@����:::����l���#z��-4ٮ(<���8v��6FFF����l��ͅ����d;�eG���;?��d!�͆�����M������#2�N!�T���d���/���k�6l����l�}�����j+KcӦ�����~��B�w3��6�VO�q	�`��3&�;�|��̺�u�7�ZS����ظ#Dd�]CCǏg�l�p8;vlMJ���L^J�Ƭp����O`Va>�:����c���01֗4D���_T��������?#���WWH�v}����#����L���M���kq���{�E<�}-��#p��Q�+<���?xyy���%DٰX,���`��V��[�n�m"�)j��W-Z��ƍѩS'�����~�z�\����pvv�˗/�ݯj����?�n��7��R2�ikk��Ç|��CCC1`� ��a��b���~~~����3��޽�;v�СCR՛tqqA@@ �&V����l�ݻ��rrrD�W�
��8˖-C�&MĚ���G�E@@���:�b��7n�,Y"������سgV�^���T���B�˱c�0b���&N���{��l����~}����������)#7���1�1:pP!3�Q7-�`�������������Q*Pn^!�l>��tыdw�؁)S�0�c��X�f�$�)RTd��
�+�q	w ���1l�0�����O,]�Td;s#��e�^�U����~��}[XX򤼼�����kg��'���j�u���I|��x�.�ji656Эkj��/I)e����pnG?ٶM�6g|�ާO�ФI��	QF���X�z�X�0 X�t)>\�Q��LMMѼy�j���b�mԨ�6m����
������3���`dg��/�:::h߾�й:t��w�gZZ��U�������
 �n�BQQ��222B������z�����&&&��҂���������W�^�����z�*^���	sss����]�6,,,`dd���,|��	���s����?F&����֭�3Abb"��[�h�o_����Ν;b�oڴ)�w�f͚������çO�������ܾ}���_��EI����u���ݻ7�5ksss�������?F\\�_��.����{���puu�p����(((�*fB!����=���=�~^^^�|��ȶ͛8a��b��Ix< 3;/?+;?���4��[Q���EA����Fɫ��>��f��:���jljj`o�WK%��+(,ƺ-���C�ȶ�����ի���ݻ�ăR#@	w�T#�fff���c�= ƍ�����lgce�9�a`�,AZ���_TRPP�]T\�����*��q��X`�r�555���)��PW7l�X�������&��l]]mSC}6[]�~N��x<:���>�{NNN�}�6�j��ѿ�;wN�0	Q���:u*�M�&�К��,_�'N��st�B!���:u���p�3\������;"..Nd��-�1~tOԴ�;%QV�����d�r8�Nyf9���^*�\���f�s ���hkih�󠥦βd������Ljii����2�׫��j/*�RPX��;B��"z���!C���2~�����f͚1�ͨ$"@	w�T#� Э[7\�|���f��p8�ӧ�X���L0� �M�BT[y9����=�+����U�JIQ֮]����K"!J����&M���׷�#���ž}���&�,B!�B�|,Y�˖-c�/%%�ڵÇ��uk�)��@CC5�����+���x���ȶ�ڵCXXߎWQ���1`�����1�pWJ56� s���ڵk����A���#����>��������P����Ūٮ���+W��m۶��	G�^�PVV3�!D�KKK ��I�B!�()555�����ˋq���Xt��YYY"�6�g��~^��bv�QM�Yyذ=D���6Ddd$����#n�i%J�+��p��Ǐc����}��ݺuC||�ȶ���9�?jۘJ"Q�%�ع���x+�m�Z�p��y�:��x��-Z�jEFB!�BQ8###DGG�^�z��޻w=z��;4�*�um�?�/tT�O"���,l���L��3u������acc�x�+W��O�>5�n��"@	w�T��zzz�s�5jĸozz:�t���E���Ҁ�XO�5r� JR���`ˮsHy�Id[�:uJ� ݺuí[�$	�B!�B�9777ܾ}�����FEE�W�^b�maf�_���*?�׉�m�y��lkkk�7n��ё�<���hٲ%22DĪ�"�"	w�?�����������ڢT���.]�$֩�%%l��<"o�^OT���X�>X�d;��Ƒ#G$J���i�(�N!�B!D�<~�'N��cܷ}��8y�$��D�\O��������$a�,�Q�o;#V����aaa%����1`� UH��U;�a WE!���ܾ}�F�b|����!����#33Sh[x�4	��24p�K�6<��?M��g��_$����&�=��C�J4����?�Y�F���B!�BHu����˅������Cǎq��I���
m��!��+XZ���D�pI���/E�hp$�\�/t���q��U��2Ogr�\x{{#22R�P�Q��B(ᮤ�������!C�0N�b���|�2���D�Ox��^�[C:�CE�x���:zee��y��������߿�D�8qӦM�h� !�B!�"ׯ_���Z�jŸ���:w'O���Dh[.�bPXX��u��FUQqI)�]F���b�wpp@DD4h �|3g����%ꫤ�@	w��2	w �@�ڵ+�zzz���FDD޿/�}Ff�?x��N�06�c<Q^�ť�'��oĉ�^OO����ٳ�D�ݻw����B!�BQ�˗/�m۶�[�.�vvv�իN�:���B�����2�=�\�i���IM��x���X�]\\!VY説]����D}�XT$�j��j�����X,�ݻ�ƍ��NN�k׮��^CC#uB��%��(��t�9p	�s�joee�s�Ρe˖����Kt���?���2�ж!��1��VD?x�{1/!�B!�(���!nܸ777����ǣo߾HII����&��D='k��#��N�>���X�۷o������I4_pp0F����r��+��ȡ��p����q��a�1B��eee�>}:v��%v�F.v�s�H4'Q,����(�qE���F������]}��-:w�$��+��:�G�f��Z��xg/�St�B!��0�������D�?~��~��!&&F��,��`�PWW�hN�X�ť8r"w������q��!ԪUK�9�\��~���,cTCE@E��]p�\����ܹs�g��عs'6m�$v=�'�S���cx�4Y�9��df�c���8v���vܼyS�d{zz:z�ꥲ�vB!�B!�-==={�Dbb�D�����~���՞��!,2�6#�S�Ds�y�����g�l�9s&N�8!q�=**
�R�d�J��5Dyy9Μ9������Q�����W�.\����2��KJ9�~��y��_�l��}���u�)v���iYb��8q"�9]]]����Ȁ���>}*Q�������F�x��/D��@!�B!�,77�ϟ�СC���ϸ���&����lܽ{W�>�9�u���4�`g!�BI���e8u6
������X�>���ؾ};/^,���{�ЫW/���KԿ�H���p��5HQQ���(�����q��-888�՞�"o�㏿�A�k��%��SF.6�A��k(,�M���v�څ={�@SSS�y��������_B!�B!�&KHH@Ϟ=���.Quuulڴ	���xezKJ88v�:Vm<����K��˄��k�1\	��r�X}lmm???�獍�E�>}���'�D�(�^����W�^�z���c4o�111����ONnv^�����S ��D�ʸ\\����G���[����?33���bק#�B!�Bj��O��s��x���c�=QQQ�[���}�$�b���8{�8ѕ	�|��aߡ�X��4���/�өS'DGG�]�v���ݻ#3�^��$�V#DeK�|��� 88͛7����DcԪU#G�Dyy9n޼	O�7sR3y+��fH    IDAT��r8�[��
���[l��?D?x��d�=z�ʕ+hР��s��]�vEll��c�4TR�B!�B~		A���all,�VVV=z4�<y�W�^�է���˄��}�9��j���TeF1��rD܈Î�����&v?��9s��СC044�x���Hxzz";����))C	�������puuEÆ%CMM�ի��Ñ�%^�o.�/�����06҅���D�ɼ��������{��/�����,Y�={�@OO���w�aRU��?w�Wv�K�MĀ,�"�(c��;���O�hQ1F�1KDX�b	 RE�^ؕ��¶)���a�6�S�����<��-�|fYfv���s��vv�F��;v4��PD�    ����͛7O\p�ڴiӤ6�x�С����k��v�Ϋ������}�>uJOS�䦭����q����gZ�n����i�Fs���w�!���T-Z�K.�DG�6�Y&�D�=(5���$9�N}���ܹ���v:u�k��V{����͛�>���R�~������G�����K���z{���ytn�޽�h�"]q�^-��e��=ZYYYMn#TQp   �槴�T|��F�����7��0t��kҤIZ�|�v�t~A��Y�Y�{sԡ]+%'�7/<�&s�A�>�+-�b�����(�q&L���U�N��ϟ�)S���ҽ5��H�(��fUp�$�4�`��\.�s�9M.����i����֭��.]��
�_T�Kʵ�Lm���R[%�uZ�o�Am���Z��j�>�K��>���?ұ�n��6���{�ܹ�W9���k]p�M^8&�Qp   ����ѣz�w4h� ��ٳ��i�F7�p���˵f��>�>R�e+6���|uJOSbBl�s���Y�4g�R}��
��{tnRR��{�9=��3JH��N�?��Ϻ��[�p4�9��D�=(5���qK�.�֭[5a�EFF6�������ב#G<�����T��n׶�������S�M���?��?Y���_��s�����ѣ��ϟ��o�]QQQ^ey��7u�W4�[�j��    �WUU��Ν�V�Z���E�ۉ���رcu�%������=:���k�:R���d���iJ[������W�g�G�w�E�?���ƌ�U��tꮻ���?�х�0�%
�A���%i��������'*>��%&&��K/�СC�|�r{ve/��Dk�ߩ���!)�C��z s�A���2�����/W._h���t���k����ѣ�WYL�ԣ�>��ӧ��tβpD�    �7�4�p�Bj�ر^X۵k�n�Aiii��oܞ��x���l�fmݱWII�j�:��U��p:�f�N���/��Pn�gu/���
�����SO)%%ū<����<y��̙�U;a KaRp���K���V�ի�>���&/�z���"���/��ы��bu��uֈ~j߶i+{���eZ�v��Y�E��5��1c��/��O��KKKu�M7i�ܹ^��\:Rc��n�`�ɢ5�d��c    @ȸ�K��[o�E��ݹs��O�����?Mn�]��yf_�yFo%%�y�)�-��[�b�V�5����H�|��z��Ԫ��k�ڵK�]v�6l��u[a`��s����Tbb�^{�5M�2�'��ܹS=���ϟ�U;=���Yg�ӐA�(&ƻiNB�i�ڑ�_�Wm��?f�no��=z�����ɓ}�-33S�]v�6n����w    ��z��>�@�I{_}���O���g�Ȉ�M#��>=;�f�ҟg���a�n}�r�vd�7���{�z��4p�@�d���t��W����'텁%���(���0�w�}z��ǽ���D�-�}�ݧ͛7{�NTT���ꬡ�{h��n����I�P����V�ݮu?d��Ȼ9�SRR������Vt�o��,е�^���"��.(�    N����W_}US�N�I{v�]����裏*/��w�KRB|����O��}:�fk����NmݱW��gj��ݪ���SO=U�f�ҤI�|���r��G�c�=&���6��QpJ��0z�h͙3G���f�i�˥w�yG�>��v���u{1�Q�߷����~}�(�Ex-�QU������ik�~ܸG���^�������K��{�Z���4=�C������O4�:�E�    P��ӧ��'���`���͞=[�g�Va��y��Er���}:�wώa7𱸤L����M[��qs��EvI�ҥ�~�a]w�u>Ț���믿ޫ���QpJ�둖���^{M�\r���t�\z�������N�v��Y���ԿOg���Q�tk����zp�\�i_�v�گ�[Ҏ]�p�f����xM�6M<���.�HRVV����-_��gm�
�    �����_��Ϧ����_z�%=��>�="¦�;�_���٣��tj�����^Yi��Cڞy���Ӿ#^Ms�6m�hƌ����Fulʠ뮻N����Y�af�(�%
�0C��z��~�i�����ݪ�*���z�g|>��f�C�T�ڽ�N��^���ԶMJP�UPX�}�;�2wTV�aUV5m��������n��߮�m����7�|Sw�y�JJJ|�n���    hL||��}�Y�r�->m7//O/���^|�E>|اmGEE�k�6:�{u��V;�)�U�O����e�Hn����ծ=��������t,�{�֌3t�5����^YY�|P�g�fF��-��D��}����o��!C���]�4�x�b=������/}���"##ԡ]+��OU��������V�JKMVB��^Od�;��W���������?��}�t���/}J�`�>}����z�^$������7��ܹs}�n���    p�%�\�W_}U�[��i��׿��g�}V۶m�i�'���Vz�T�wHU��?�^~��DG�fz����U*7�X�y���/ցC�w W��nw��OI5j���>]|��>�y�f]}����|�n�Z"
�A����"##u�}��GQ\\���߸q�^y�����>�k�]�1�j�2Q		�JL�UbB������bb�~>.J6-��$9�Uٝ��*=Z��e*--WIi��J�T\\���q��iڴi~y������뮻�ҡC�|�v���    �DZZ��}�Y]s�5>o��ri�����?��O>�Dv�o�oHRR�Z$'(1!VI�qJL�UBB�����Ȩc���9�.UT�VYi?���J�?�]J�V���
������y�ݕ���_��W�6m�N?�t��_UU�'�xBO<�*++}�~�Z"
�A�����w﮿���3f�_گ��Ԃ��+�諯��֙t��QW]u�~�ߨK�.~��������;�������pF�    �g�}�����SO�K��?���׿jӦM~�#\�~����u�W*11�/}�\�RӦM��͛��~["
�A��{��o�Q�f�R˖-����ݻ5w�\͛7�[i~֮];]~��2e�222�67�����/�����w*..�Kᎂ;    ����c���;�Td��d1MS�W�ּy�4�|�۷�/������kʔ)�2e�z���~�����C饗^������QpJܽ����G}T7�|��^��۱c��͛�?�P�ׯoV#�;v����kʔ)5j�"""��߲e�t�=�h���~�'�Qp    x����={��f8��riŊ�7o�>��eee���`3h� M�8QS�LQ�~��ڗ���믿��z���63KD�=(Qp��޽{�g��E]��rrr�d�}��Z�`A��+�3�<S�Ǐט1c4d������۷O=�����5��B�    �+cƌ�_�����7 ��޽[_~��>��S}�����H������ѣGk���7n�:u��~W�^�{�G�V�
Han�(�%
�>4q�D=���ݻw��t:������jŊZ�|������}!))IÆSFF�222t�g�m^��i֬Y�={�����o���    ���h�u�]���~�V�Z�߲�2�^�Z˗/׊+�bŊ��~�}��1b�F��#FhȐ!~���D�v�҃>�y����f`�(�%
�>�+��R����u�)�X�!;;[k֬�ƍ�q�FmذA{��	�Q۩��4h��hȐ!8p�ߧ��Kii���y=���*((x�ᎂ;    ����5}�tM�>]-Z�x�.�K�6m���_]wٸqc�L�ҵk�����5t�PKkT�ӟ��o��pX�!�-��D��O"##u�u���V�.]�����RmݺUYYYڳgO�����������<�,P����֭[+==]]�vU�n�ԭ[7u��U={�T���}�l�SVV��^zI�f�RNN��q�w    �?�j�J��{��뮀�)_�#G�h����5��������ȑ#***��0������4u�ܹ��r�ӻwoK.B�l���z����ꫯ�����8�j�(�%
�~����Z3f�������˫.������tV�"UVV���*���H�������(���V��GEEY�TPP��_~Y�?�|��{�(�    !--Mw�q�n��6�n���8������˫����Ree����$��622R			��M����8���U�_��]S�ܹS�>���x㍰��>-��D�=�F���3g��/��p�����_~Y/���O�&�=�    ���S�j�̙[\Ǭ[�N�?���̙#��iu��b�¤�n�: B����5a�:To��F�L��i�Z�t��N��=z詧���    @����[o��hҤIZ�x�O��E�*++���jĈ:t��z�-��h
������_���j߾�n��}���VG
z�W4p�@�s�9�7o/�     4#.�K��.��u��Y<�������6�mۦx@�:uҕW^��+WZ	!.��aJ� 1t�P�p����˃z��`TYY��?�\o���,X ��nu$�)e     �#22R]t����:�7NqqqVG
)���������kŊV��1K&S�Pp�_�l6�1B�'O�ԩSնm[�#%�өU�Vi����3g�rss�����Sp7��Z�QLl����������i�K�    BW\\�ƌ�ɓ'뗿����㭎�
��'�h�������UUUeu$ԴD܃� �ѣGk	���u�)�X�R���/��g�i����Ϸ:�X��C����s��c���ʊR�ڶ\��o��
�    Z�h�	&��/��矯��T�#Y*;;[�-ҧ�~�ŋSdnKD�=(Qp!={�ԅ^�q��iԨQa��ri���Z�h�-Z�U�V��pXnj��ޣ�(u�>$��<�g�J�ٹ��}�    �DDD�3�иq�t����OWDD�ձ����B�|�-Z��j�֭VG�����{P���"##իW/eddh�ȑ:��չsg�cy���L�ׯ׺u�|�r}�����˳:����{j�nt�Dy�Ժ�UTp��
�    �5x�����ȑ#���bu,�k͚5���o�|�r-_�\V�B�,��D�=����C��v��h����ڵ��sc�%//O6l�ƍ�q�F������Y�4��Wp<�2�J��C9�2�qݧ��Sp   ��'22R�i������k���8p�Z�nmu�:eeeiӦMڸq�6lؠ���k���Vǂ�,Q��#� �'33S����?~����d���W��r��u릮]��k׮�֭�:uꤨ�(��9t���٣={�(++���[�lс�G�90�Ҫ��!��"��    ���ph���Z�~}���ڵS߾}��.'��}��~�p8�o߾u�={�h׮]ڲe������/�k�R����j�*�Z����-Z�P�֭���Z�������$IRBB����e��]}�QAA��cs}���(//�֗��̓DȈ����:/���qVG     �C��СCu��l5j.'�^��}�LII�a���������nWii�$����V�%''G���{��?�N�pCQQ�������iu4�7�Q#B.0     ��\.���(''��(@вY        �p@�        ��       �Pp       �(�       ��       �
�        �@�� ���Q��~k�S�.jӶ�����j'��>9��r؝�/,�Q:����#Gj�ڵ�����/)1NqqǞg��銬j�K���P~^�v�Δ���*s}���Un^�_�      �C�a�]���͍��ݴ��գ�(�'�����݆��V蓶��N�Q�${�:::zݗ��\{v�Ҿ��L��;�;�j��>m      hw0CC��9眣�O?]mڴQrr��=���effj���Z�|����<j�u���ܹs����B�ڵ��1Ç�E]�nݺ�S�NJHHБ#G�o�>-^�X�-�ѣG}�\���.�ԫ�9�������8��w��Zk��/��� 1��ztoou���'밾Y������5W�ku������:t���    �B��������u����o߾;s�L�g��s�=��R���<y�^|������&M�$I9r�fϞ��C��{��7߬�G���g�լY����%&��g�sD�ݷ:t���}:���Q�g=O���X#hDGE]�}����˚����� �t��A>��&M����t���h�ҥzꩧ�|�r��A/>>^3f��UW]��={��ph�ڵz饗����4}{g.  <�hju��UK�.�믿�h�����=��cڹs�F��U�����.]�`�����=���Z�n�:t��U��Y�n��0(��C��[   ��1B�6m��߮��c�%%%i���Z�l�fΜiqB ����k�ڵz��Իwo�l6EGG+##Cs��ѻﾫ�H�, G��	F�����kĈ����1�ڵӗ_~�����I��{ｚ5k�l6���z��ŋ+**�I�6w)��� ks���Z��\  4E�6m��G�e˖u�7CO>��&N��d@h��lz��L7u�T��`* @����^�zi�JI��`����o����?_-Z�PLL����4d�=�䓵�r���ћo��s��l����멧��~l�����ok�ԩ<x���飱c��駟VAA������[o�գ>qLtt���Ztt��   B��w֭߭[7zܟ��� �Bτ	4|��F��1c�RSS� ʸ�z��w���\c�޽{5i�$}���5�WTTh���Z�~�^x�͝;W��;��t��A�2t�ҥ��+W���W_�ݻw�8f۶m��/�����?԰a�j��[�׿�խ�pf�����4M�Y���h�4n�86L�;wVUUU�k??� ���?ޭ����.]�(;;�ω��r���u\ll��;�<͛7�ω  ����~��_��N�����:묳��u�������hѢ�m�V>����N���]�V�w�����=�����8q��o߮-ZTo�ׯ��w�^�P�3�K�<��1<r˵gZ^����������9��O�����;�s�=���o-H ���9��ѱcG
��I:v��c �w̘1��c�4u�M7���ѣGu��W���Q �����c��ȑ#n�c���������>|X����������C�@��v�(�U����*j���ڷkW���Ҫ���=:'))IQQ��z����#t�/���ң����<:�dg�>Wɭ�v���r���X��v)?�'�r @s��B�,������ 4�w
7�v�i�ӧO�m˖-�=j';;[/���z��mqqq���+��sϹ��ҥK�e������ok�۵k��� .RZ��ߐ���u[GW�`�G��o�^��R��:{�F�.��{x����HG��    �X4�Mcǎ����^kR[���LӬ����v���K�z�_VVV�m���� �.!)U�~1�'�v�WZ����x�x     �0��MC���mɒ%Mj맟~Rff�N=���m�F��a�
�uY�~�G����Q@s�iK���kN�z�,\]kێ��=�    IDAT$	�S��RDD��1�Vi�պ�)�9�iu     �F��M'/�r���ݻ���}��w5
�Z�RJJ�


=7''ǣ��=Zk���ٲ}��l��o>))I={��(Q�|�h��,��^Nu��kۡw    @H��ꦴ�������U{�QڪU+�
�u�XoH]�����4q�-x�A�	)VG  �`�u��.~���G��Ѳ
��ߦu��w��ڗ�U�m׻�y6h}����؃W������i����~����g꜑��ǳ/}�쟎��  �A��M-[��񸨨ȫ�
kmKMMծ]�=���E�� SR����+5 �l��#�	l�� �$&&Jqq�������m6���!:�w�_6#���'**���#�� @p�������j<����t:�:�娤LI�$9~�f��*���V�      �	
�n*,,T|||����d��KI�}�|]s�n�/i�$�I�]�r~��.�O�s      ��\�)??��㓧��T�V���5�ШÒ~T�b��vK���8      @sE��M���{���D���k<���������)��M:6_�;2%��/      МQpwӪU�j<���������Vtt�Tc[ff�\�Ɔ('9 ��MI�~�      4s���o���ֶ)S�h�ʕ�5q��Z��-[��lh��pN��S4+111;v��:�,u��A�g϶:�G���+++KK�,�W_}%��nu$     ���w7-_�\���5�]{�jѢ�G����o����E�y��Te�΁�Ѝ7ިݻwk������5q�D�cyl�ԩ�9s�.\��;w��+��:     @ؠ�����5��j�J��_<j禛n��g�]c�O?���>���h��r�
��x,**Jo���^}�Uu����8>ӥK͙3G���"""��     �(�{���WEE�	����:��p��K.�D�?�|�����t:}�Mr��i�^z饰	>m�4͚5��      !������u�=�������^}���u�V�y���z������+66�ƾŋ���_�K^4�%�>�⢋.�M7�du��1c�F�eu     ����������Ç��믯�}�ĉ�0a�V�\��k�����JNNV�~�t����Z$U�6mڤ�S��4� �G�I��YR��ǧ����y��#�����i�رV�      Yܛ��o��Ç5s���m6�222����h_}��&O����B�Ds�WR���F���4D���oƺu�aÆY#`�;�<���)77��(      !�)e���r�Х�^��۷{tnNN�n��v�;V~J�f�&i����[����I�o�@�8��#��f�СC��     ��>�H�~���N��I�&i̘1JII�u\ee����͛7Os��QYY��}dffj���5����x�����V۶m�9CR/I�$��؈w���jo#
�MԺuk�#\s|�      �B��K�Cs��ќ9s���t�k�N-[�TUU�:��;w�n�7��ŋk���^e,((Д)S�j!"ZR��!'��Es|�      �B�݇��������
� �Ys�d�֭VG      Y�� �X�n�rrr��0�����"     ��Pp�zTUU�o���1���\.��1      Bw h����geffZ��6nܨ^x��      !��; 4���T�&M��Ç���7{��ե�^���J��      �4
� Ј͛7+##C�V��:��-Y�Dڵk��Q      Bw pî]������/�\�~��������d���5a��=Z{��:     @X��:@��p�/ԭK[�c@�W�~��?Y͘����￯��_�����v��Y��3-Z�Pqq��1     �ȩ�tи1�[�����VX#hQpoD��mԿo�c@�w[ڿ��Pdd���i�:�Ǌ��C��N�    �R������h�#5���Tv4��a�n�PUe��1       �0�pӡ���2���1�ҡ��d���1   p�q��)%%������>կ}^>y�*+k���p84�|��4h������j�1��Z���Z�����j�o߾:s�/���ik�_�*E��͓��lr;�z�Ґ!C��w��J�ܱ�m����v����n�+V(;;ۯ} P
�۪��*�U��Q�JEy��v��:   Nr��w�G�����W����J����n��V��pG��E�u����ֽ���T��5@:�T}���*+k�]�z��}��3�N�ٙ1cw �%�Rp�i����=���(a��8G�W�/����(      ��ᎰUV^������ݍ�^P�Χ�{��Jn�*�-«�$����2�.S�U�-���D��r�����c�����Y���/�L��ꧬ�ړ��V_��_X��6     ��PpG�:t�@�_���!%--M��������e�2��      ��A�@���\�#���HEEռ�!..Ƣ4M_;�����      @x�� n�t�p�9gp�m.Ӧ��[�5�sOL���Ek���5�     /,�
       �Pp       ��R      >3p�@]s�5JLLԞ={TXXhu$��á��"mذA;w�:�4�"��zK���W'I	?��|h��RIG%헴��m���6yM��������[    ���fӒ%Kt�YgYa�4M���;�6m���˭�?����;O3F?^�Kʕ�ƩI?IRIg���4�E��?-2���; 4Qd�M?���1<����:   �0��Rl�������J.�K�^{��q�C��I�\#]w�Ԯ]��N�Tߟ��Tl��X�[��2�>�N��      ����j	V�@���ս{w�c�K�!]r��j��i�4sf�b�?%K�F��6���5M�B��      �ddd�0�c ��!C�X^�<Y��G�㏥a�,��Gқ�v��n�Wᝂ;      ��r����0VZZju4���J�.͛'`u��IzY�w���n<��p���S�V�m�c�϶����)�T�c+���]�V��xRX�G��9s�222cu�������(..N�ij׮]����j�*��   @���͵:�TAA���������(pSt��?H��{��Al��妩J��0T�F�.���t��s%��E���wIʒ�ZRW�EC�6l����%%�r-4W}��Պ+4e����{V�     ?3MSw�q��=ju��sgi�\i�p���͐t��1��+C^�ȴ���_ҵ��J���l�����0g��x�����?W�  ���W_U~~��1����ϫ���}���>J�8o�[�N7�|���4�{��2M���oܸ1�yau���}��wn[VV&����1v�]�C������r;���Pyy����Saaa��3N�������|mݺU999�ԩ�*��t�Z�LS����z�\���?m`gu���v/�L��?�-|�t t���4u�a��4��{���%�,�Y�r��P�JJ+<>�t^��L��9���C���s��)JKKk䮪��l.:Oߴ��r��p8�j��t�����󊋋�������/^��o			:��s������(   A���8�
�QQQ^�_YY�����F�mު���~�##�+�����yIMM�:�0|�p�^�ڲ�;t�X�?��w��a�V�c���c}^p��n��g%[h�#�y�ToIw��T�w�=A�M�����}�y��֭;��V����#�C�۷���tlm 
�      �1��'�����$>u����_�<I�k���h�-�95�b;���H      ����aWl?n��OLS���菂{/I_Hz]R?�R� p[II��     ~�S�����n���~5F�\��l�_�I���Q�y>l       $fΔ���q��=9�Ws��JzS��>j/l�q�r���SOY��U�V�6m��      B]���u���NP7��v��q�`_�J����@=\.�x�K3��ٓ�;     ��J4q��2���'MS�C�6v��S����(�      @ز�\}�犏��:�"%�k�Jk�@o
��X�=Ջ6�_��       ̜>l�ڶ?du+u��Bc5��>Z�<IqM< B����U�]N��    �2���6-R
5`�z�c����qД���>�ӤH &Lӥ�B�c���$��      e��DN�c��MS�������C�g���B�Kʬ�  �޿��n;���     @���c��;�:F0�!���vzRp��4Wj|b�p�����p6��������v����|�c4��������      ��������Y��tO
�%�M��q8�P,Xiu A������0x)�ۧ�~,��:�e��14��    ���'��ݲ��&�oYBX������f�����	1_-�A�NMנ�ݬ� UV�j݊�Jk�]im�+&6Q����TEy�r�V�,y�v~���,�+�{    +1��A����f�<q�;�dI��'Sh0M��K��Ԏ����:� d��r�RΡ]VGAʏ���X�q�VG�
��Z    ����yj�>x����Kz�č�L)�'I��(������z|�Ճ\ �djώUV���U�ڗ���1    ����w��B�5'oh��>X�m��z�\�
�� �ܷE{�|ou�����u��n��:
    4K6�K���au�Pp�i*������<���ti�g�=<�!� ,vnY���>QQ�A�BN�]��m՚o�Qa�~��    @�վ�~�ǳ���tl��j��>H��~���oإ���>��( �&8>׾a�)2"���1.�qj��߰e���x�G�z꩚5k�z��U�1�ij�ܹzꩧTYYY�q'3Cx�J��l�օڹ����    �����N���1��~�AC����ZLS����u���u<s�@p2].�]^x�Y	���:x$ǣs�Qƨ�u��몫�ҙg����49�N�ٳG�/��/���7z��f�I6�������|   ����p_�����J�5M�C.���{�4��f�N]6a�RZ$X ��8�N͝;Ws�ε:
     EGW)��gĚ�TI%� �?6�1w{�\.�֬so� ��       ���m�0�#�Cg�C}��$d�X���       ��F���*L��R��Z]�a�z.Kh:p(_���6~ �,f      Z�Z!U����}| ������1=�� \�)��[Ҏs݂M����E�    4G�po���u��`���m�>]4vh��0�; �ֻ_�w��:��r��u��V�     �[#c�J�#������xIg6K�ڵ��v����n     ���l6�����ryt �4v/oT�= 9�L�i*�0Tqr�8CR��B���������#����(??_�����0%$$(;;; �    �.??_���@��X�2*�* 9�P�T���ߊ$������� �p8���gu     �f��\k�dI9'߇ӫ�#Q��G^D��       B�a4V�G=l��9w:Rhu       �	�=����X�]p?ł !-'��;      ��`���T%R�{K�����F0�T     �d�ɴ@0�WE[!9%�K5�6I��	a���       <��D����z�'�T{�;�r�d�;��       ^+*L�:B(�~�'��,���VG        �0�x�Yp/� HX���!�9�      �
�MRg���$Wೄ�����"��       ^�=����h��?�Xp7u����4�j/�      ����8�Z#��H����ȓvHJ
h�cu     ��c���B��fSTT���{lC����EDD4z܉\.�����^�4M��s8r��7GII	?/v`_�Z��Y#T,5U/�yr�}��΁��ڤ��:|��7���EF����/�6������)��V��U_�6�������Ng��Y�ͩ.���r85�;޿����LӬզi�2���
L�TDD�


�    �/���(!!A2������Of�٪?�:�N�\�?���9Z�bccUYY)����>7WUUIjx-@��%��^���N�G�����F�	v�������:F��o'��������\�.���e	}m�6���!��m�V�a�������.7�e��ݺ*ZW_�&::��M=ڴa0    @����+???�}�j�*�}���/�?�ewVUe��c¿>�%���N�PW�h�&��͆��Paa��1�n�    ��C���o6�����;{�w��VG	v�5�=q����l`���ޞ�7,     �	~�F�[c��VG�:y�ɗ�VJ���J�n��lZ�b��YY����G���
�      �Q��ֻ��v�:����F�3������-p���I��{��5��
D�P�r�������g��v��i�����ʪ>�S�N��_Y     $��	|O}+'�H{��o���t:T���Z�zu���~�{魷�H�7�����	��+
�n5j��x�u��Mұ���{OӦMSQQ����/�p�?~V>�t�>�|���v���    �V�l�{�p����x��⋺��k����M7ݤ�J��yGz��G+����^�kG]�O$=��8a�{����ϔ��P��0M�<Y-Z��\`a:�q�pw�����Q    ��1`������k���+���ƶ:裏>�Yg��5k���f͒^yŢ����Pn];�<���M�����?�(��h�ر5jT���7H    @ ���/���2C����Ul?.::Z�<�������~}�҅�C���og}�c��,�eذa^�gxq     h~�	������b]��n�Er���*d�0�;�x}�IbR�F���7�?!!��{	     <������5V�<y�ڵ�k��3Q���0�nC�Wp�'i��� &�a    �����48̘!m�nu
KH����Z��O��Q A�W     �)�	�����PZ*M�"��[����C{;0��}[%-�4�W� o����;  �^{�ڷoouIRUU�.��R�ڸ���5y�d%j��_���S�L�u�]�4���/����&�饗ꦛ�0�g϶:�����	�c�鷿���W���s����9����$=,�bIQ^Gtx�  @}���ԥK�cH�*++�*KRbbb@���y����ʫ�qqqA��"I6[C7��9aJ��^xA��C��n���$��݃{�$�y��       p��-9p#�̘!͛gu��X#i�a���	�\�����M��/�     �.��z�.�t��_X�į6Ig:��I��K$ݦc������=e�<    @ �94<P
N��҄	a;�}��sC�����f��2      !L)�We�t���/[�ħ>ձb{nSN�d��%�lJ'�/p5     x�4̀�X�͍�)��7�}�Iv��i�bJ�-�R�PYS���.�JI����
���)�     �S�B�3�HҞ=V'i�"[u�'����KnY��J*��S ���Ƨ�r�    @m|� Ik�JC�J����I<�A����h�)��l�t��
_ �@����ڵk�ݟ���-[�0    �����kÆ�����Tfff !�0�=���K���t�R��ZI�N��P��m�RK$]&騯� �����������VEE�k�N�Sw�q��    ���NUUU���p8t���4MR5�Ͼ@�X�D2D�9S�ɱ:M%�����0��aȧ/Nެ�Pҹ���ۅ��$��r�J�}��Z�l��N�\.�֮]�.�@�~����     �-[�L�s��/_^��kժU3f�/^lu���~�`ȟ��Ji�sq    IDAT�,�S'�[�}��u]�u����0�a���Dzy�ZIgK�TRw�� g��Kǚ5kt��g+66V6�MeeM^t    p��+Wꬳ�R\\�$�����D�PO�w*+�W^��|S?^��i�8):��]�tl��Iz�0T���-�K�VI�I���)>h�/�pWTT����h�c��_�ӑ�"�c    �ZrR�&�nu�����e~�z<*+���?���*]~�4f�t����h�(uS"i���t�Ⱦ�G��w��p�+$}+i����xQ����)�0�:��a�ټ���s6�2��h�����[ê�����X�_?Ye�]%���qGZj�%���o  �����h$�UjD�=**ʭ5�����k�٪��u\DD��PDD����Z���h���r��?����<�{qTT�5���ﷱc�z�i��p��v�s�k���5����G��w?BW^�������з��K:SRoI�~��$��Nɔ�_�I��Z#i�a��*?�U�]:������$]�öEDD�e˖�n�^�4e�"#���6M���l���|C9���x�'���\�:��'�ur'������j��0���x���`G�1'g��ԦM��c�c����_�󨪪�>�4����A�W&O�3�;����~������7�DD���#�Z���/~�m;��   �%�S�����)�~�����LSq�%%I2$�Tb:ؔ��e���LI�؈��%���4C;w�:   �l�X�BYYYՏ�um�Iq~�sӖl9���TUUy��Ν;��7KէgG��jH^A�~�����w�[����4�qÀm\S�@0=�8���	-��&y6�ݰ�6,aY�&YB
ReY ��`j�6`0�6Sܻg<}���!����H�#i���҅5����<4sn=�~
/�͟?����Q���CRe�fmＷ���@�x��wy衇z<6n�pF�(��oo�[DsK���/.�|���	Z�V`y�YrQ����w�.�_�Z¹$I�$IEt饗n�����i&�9��s��ױ���$c�}��̘�8�^xZI���o���.x����oL�	�����*�^�ǯo�k��<���<�p��S?�Q>~���ћ+��v�~gII�$)�,�t nN�R�9%U����-������x|c�X,��� ����g�K$�s� ����  ���W<bĻ��v�"��Vf�\I�$I�$U�R�7�~���+p:���4��
p�1��ӟ���c�X,k�Z6���,�K�$I곭���aЖ�{uH�<�,�ڀ^��p^<�y�b��@��u\~�����yY���o� k�l�)�پn'�tR���K��Up��[�%��#�?� � �_�7���{)��"�`�*tm.�U��$I��ɸ'3f�=����O�T�9���-�K*�(
�Z@����?�v&���I�@;d��u�k�E�`>е��Xp�T�,�K�$I껐0��?�M-���.�w�	�]��$I�$IR.B�Xp�TN��HRq����-e$I�$���6��.I�f�]R�$�ɨ#T,�$I�T�x<�����T6�3��.I�$�0�p�$s��T�8�!��{���c�`���@������H��9{�_�����7a�]R�Xp�̻?%I�$2�Yp�*�^�Q�g�V�
�§�G���g!(��wIe�J���P�\�.I�$��3������kc�S�/�m���">�����Cx3p=oi�^����q�{f����$I�T�,�gb�]� w�W�I�����̅�?^�	-�K*�.I�$I%a�]�\�
�x��6�8x��~�T�Xp�T6�{�bI�$I��Lfܥ���<q��L�Y���C���z��0���c���`ZH�@�Lzڅ�� �L_R����K�$I*����4U*� 8����@-�#�!����bi�=L�?	|�t�}�<�X	�f|F�N�_)��,}��{fA�/��$I�
a�=W�K�4��ɨ��j p1�)O�`^�����(����SxӞ�������!��V�`y��K*�����#T��%�$I�T.��6W��'>�/0�D��~�~��-d��,�!��� �C�_��o1&������9s�)�� U���Ψ#T,עH�$I*�-e2��.��i��Ti�}���[!���AJZp!�gH/:��t�l���HO~��e"�W��^���$I�$I�N�!�9j]�A��{��>��KVp�8�ҋ��/�<�ڋt�����"�"�W�����$I�
���#H�.#�k���g�0���E_m�X�
��b�]{ �^��-��h�H�JZ�Lv�Je�$6��aHgg[RI�$I�Yv��Ȗ2R��\u�R�"�|#�O*j�=Lٯ�s�R�4�1�_�[#�"�k׮���O�z^�9�L&�=�7j�|�S7>��l���g���Y�RI����Ɓ$I���Lv���'�k��w'�Ȩ�뻅K�X�`!���477w�n��T*EGGmm�/X����l�d�)�'����t�k�k��!\�%�~BQ
�!4 ?"ݰ�jl�|�@K�q���������K>����hZ�{��$I��J���3y��Q����n}�g��uIy9��o����!�C.'�\'Lo=�UVl������Q�$I�$I�G��ڣ� )/����+ݯ!�;�*����O .d�J�70��檒$I�$I*����mn$U��b�ب�D��¬���\pa*�$0��cT�����AQ�T�~sC�$I�$U�d2uI9�.pt�!��;pe���Tp�@��6}��J6��uI�$I�$I*� ��R��/v�j�u�턼�터+p/0���*�P�o���ύ8�$I�$U���z���=_�9ZZK�Zb�F����K:GӺ֢�U��-m%������,��,��*�0� �r�3j����?A���*��0xU�pm$p?p�,�,����k���	{3~�}�>���^���/}��h��O��~P��}��;iom*����--Y�:���L��;K����d2UUy3Y������y���^�IU��sQ��$�_~�����a�z#�cqrU�]�[Iw&���
I)�Lr��G��,_�u����Ƞ!��rV?����j�ah(�j�XP���$Ie����J7�p����dzp!��C���y��p�8�x�����eQ���d2�#��uI�$I�LKk��*���.QG�ԫÁC�Q��g �w?�Ӳ�>N���/]|,��$I�$I�TVF���a����C�&�skU�uI�$I�&s��ϹR��C��k*U��H��V��v�`.E��������uI�$I�fժU9��r��&����I�or��L (e�ZpF��Zpaw��J��\�uIY�?$IR���O�tފ+�={v��H�'��� �|��&�\�.U����_�:F5�,��6�@��b'��?�:�$I�$m�g?��d2�yW]uUN�I�͟��'�-[���{ｗ�s�!Q�b�]*�\*>�t�����Xpa��R'�6_�o5I�$I���_��s��h5m�4����2���GSS_��imm�xμy���׿^�T����b/Pev��O��x��B��:�=v�uI�$�落���N�|�2��{�)��UW]�{�ǕW^�.���㍍�\}�����?���3Re{�G�:u*?���9��C7~����[o��s�=7�U�ʟ+ܥ���㖅�p$�!d(��08�����W��:�$I�z4t�u
�k�u���y����f���b��vcٲe̜9������IU�^`�ԩ��NL�<���VfΜ�F������93['rmb0	x2�p?��bn�` ���CH�*^"��+_�
�����c�=0�z�Eimm�����{�k����ӧGI���0y��y�嗣�"U����3���cHRd�}::�NQu�������e�NgD@�TѶ�n;��><������6�l�ĉ9�Ӹ�������q*I�$IR���F�	�����ހ�&�5N�$�͋:�$��b1��Ϊ-�w]t���7��"I�$I*�9s�NP�&m�CO�xN(c��6���� I�@'�t�f�mՊ���4(��$I�����'�W�G�1HU���QG�$U��}�sQG(��Çs�a�EC�$I�T�0{=���e
R[v����z��� T�8Uj����룎"I� &L�:B���QG�*�ʵ��u���f+�.�$I�Bcc�	�R=� h�i�A����A���?�uIRY�vm�J���nR��;�M�)���68��SH�jQ�����/�^�75�)H�
lQpw��|��wI�f{�1�;c]*��'��:�T1���E��<�~;��$I*�u�NP��+��p��әꅻH�����X�zu�1���of��Qǐ$I�$�HB*u��U�z��"R�fώ:�$�¬\��/~��u�]44�F���^z�o��Q�P�:t ;�8����C3[ͼ,g�6�n���S��@��Q�a�I��������/!���ؘ�L��������fms�Ɨ$I�A ��ʽ��`˂���no����l=�$I����C�'?�	�vX��<X�n7�p_|1�M�a���O�|��b���w!�܃�<O,qw�cT�X���o]��ld�g����cێ��{�S�������w�J�$e3t��>j�-��F���`� IRq���q��=�I�&�Ht��[�y�Whmm�:�$I�$�L��ŋ�NQuR@lRp! E��jeٶ�ݶ���c��٩QǨ(�>�2+V�:9*K�,aɒ%Qǐ�� N{}����2�Ѧ:�:{>v�_$ո�Cr��okVK��=��J��v0wn�)��rB�|��`��&�ʦ�#����:���b�GQ�[ҫы/�+[�=ƍG�,\��,sJ�V__����Y�zuMn�[k����A�FC=h�ٌǂ�`y��HRj�Z���/{� U��w�'��:E��ػp������IÆ��+�dٲe����,X��ŋs�e�1x�?bT���sO���?���ļy�X�j/��_����&I�$I%1qb�	���ش�n�־d'I��رc�1c��o�ƈ#6~|���\t�E<��S�}\���ԧx�����g?K�&w����r�-����0�$I�$�ƤIQ'�J=�p_�p<_�44D�B�"u�M71������{on��2&�
��;p�-��������:��|�+eL%I�T{��#H�f���6�ac� Raz��˵�1th�	�~���� ���x<N"� ��H$���g�ȞWR��u�b�s�ud�Ң�n@�s� F"�}�����T禚���8��ó����|�}�ݗ_|�����s�9��g��_��~�;7I�$I�T3ƍ�]wy�-��Q0}ÓD��k����a�z=�iaP�v�ml��V��X=p�@����x<N]]]1�E�i�2�{��c��1���G}�wU�\��'L��n���ܹsK�H�$�w��bԘݳ�O��u/m���!��H�YW���q!ҹ�{�l�2 b��������z��0��e���������/Yϗ��K��[�_+��mx����60��y��.��z�o��&L����nu��S�o΍=��sǍ�ל�4�䌷7>yNöy#�1rѸv)kW-��|鲦���GAl�������w����_���}��D����ZZZX�z����ڂ�$I�ڈ�vb�IS������S�9^�u�R�;,���[p��#�>��U�T߫s�ܶWRT�[s��,��� 9rd^s._������(�Ŗo��������T���90��W�^�c�=���MWaI�$E%L���P����NR�q�%Io����s�'�_q��Xp���]=����$I�*AX��xJ˂������:F5x��ny����j�Ԇ=��:�TU,��,ȡ7�$I�$e����Ă��W7F�l�E����4�,O�����AEC�*�3���$I�*��Yp���a`~�!*Y3��?��+N k���JT�:��o���$I�$Iѱ�{Fܥ�J�u�J�kVu�`O�8��!LMh?�Ш#HU��=\�"I�$� ){�gd�]*����CT�v�=�����f�mGu��Xp���2�$I�
��=#�R!ځ�D�]A��D����vi�T��@��{GC�:�{Xp�$I�����.����CT���d:��+N !pS)Ղ?D@RM��.I�K����֨�[���࿋$&t�{&^oI�� �u�Jr!�2Ld�����q���H�#�ͨ�HU��=��"I���٪�������S����^�]ֶ��)[I�5)/*2���QG�j������Q��L෽���=5�	�W�D���ݨCHUʂ{�\q!I�$��+�3���T,g��7Pm�
A���2�p��LQ#ՈE@�b�{f�]R�n]+��~�����
FgnO�+ V�����Ǩ��x��!B��e�wY�z5��_��5k�K6�$U�(2��.�2�K��@��s�[���� ��_������G��I*&�����.�_�S�y�=>��θ}��0mM�肇�
-�f�����kK��}��tI�e�p�̂�TL'�N�Q)�[ �].'f{��>�����o%��\��3�,�$I�
�����w��.�/���4�O����+N Ӂ�*������!U9�=s��$I��B�R^keb�]*�p:0-� ��:�Zr��\^q�V�9R�X
\u�Xp�wI�$Iq�{F�x��5-�Xp
5�|�}�8V��IY����k�Zq�&�R����wI�$I�TU���G�fS!x?�O̸i��CG_�w�Zppk�!�q�e���а�y2���󺺺r:/�L2b�p�x�A�I��$��Y�J��}�T��0�}5IWW�o8H�$I*��n���5J�9�J�p]!�M������6:::��蠭��T*Eccc��Z[[����z.�Lf�wƌ9��7k�c�I�x�	���`y_>9���z�>ԗ��ի��Q��jȣ�>Z�9ƏǱ[�y$I�$�R�k\�3������h���=�D�����g޼���!� ��Iw`������j>=ۻ�y׈ ��SI�+�/�N��Օ$I�$I*�T*Ek�ZZ[�VM�]R-I�N ݡ���@��B��G� H/�>h+d�j�
̉:�$I�$I�$U�{������A�b�W� �ǀϓ~ۢ&%�Ӂ'�"�OB�.I�$I��w��H7KYq�^� ����b�w� �{�� ��bXE:I�{g�A$I�$I�$�j���@F��H��"����\AG1�S� �?� ��'Zͤ���uI�$I�$I�z��s�I/&_e�҅�=!�2K1I��O��%��}Dq"Ec)�๨�H*XPݻaK�Ty�8A���a°B[�I�$�?ˁK���g �k�7�?(U�}S�x&�}I/�h�������EQ�T�0���ψ:FEY��fnF�T�Fm�50�����*Fo�"�����&>���������S���\P�8�o�+t��o���PNH�)x�Lf�4�3_HR945�z��M2Y�[J��*����I���SB�ke
x	x�����.������\L�j�)$�O�]j��ԏ�R!y��U$��l7rk>ul�W���#f��u���+x� V_����[K��o�0l���S���._c�]R䚛ۼV�f��:����~�������
�`ҕ���?��	�Mz�\�Y�1V�(tVE)���%!���2����o�DD�$I�$I���5I����ca��
�Bz�w�X�����R��A χp�mҍy�*��XCz	�� oZ�$I�AA-�N�x8ߡ�a����� ӽ�a�hn,o I�$U� �X��E/�������I޿lS��r�H��~%�NA�$I�MA��~J�1ԃd����u�k6��    IDAT�$I��WI{��2H�r� \H��NY�����b�$I�$I�$�4ʲ�i ���+�Q�Z`u��[Iz5���n��n�#I�$I�$IR����L&�����az����#�?� ��8�`�Oa����Y؟]�$I�$I�T^e-�o*H�ğ[��@��I���X`(��g�If���뀅�\`v K�{����-$I�$I�$IJ���ޓ ��~<qI�$I�$I��R��$I�$I�$�:�$I�$I�D�QG������2�$I�$I���)���M���?�^Z�Lz��E��{}�	��#e�]�$I�$I�Tv�G'���2^�G�?	���S�ǂ�$I�$I�$�,�� _�cc�zl�����A3���X^�9zewI5'��#H�$I�$i;� ˀۀOS����W�pS{�zB�$I�$I�����x�04��//�pW�j"�$I�$I���\��Pe��	���¨bOP�=��80�tߞ�������Z���.���w H�?�$I�$I�$�''?#�P�B���:����(u��a�8��;v#��?��� 3���� Y���$I�a�����S�Q$�˘Hh�F@W�����I���$IR�j ~|'� �ۆtk��B8-�%�A�=Hz���Iڇ�~~��nt�p2LV���m��$IR�	;�|}��mǒ�����AC�#aK�������7�$I��f��䨃�͑��N�B*c��@,n>Ka���!}��m��5�E��$I�$I��b;x��-�o0
�k�T� eX�N�|��su�5������ �?���
��O[�ͦ��33�`՚uQǐ��-[���<�\���k�U���c�� 6���%aW�9r�A/8F��]@X�8a��t-�C��,[�[��_����:�#��V�llU�D"�I'��q�����96̚5�o��ٳgGG<��ç�u���ڜeQG�T�/��b6E-T�m�p~_(�p?ҽ�n�|J�n�G�sH�+�A�	��u��2���%En�5�}�����v0���_�(L{sa�?jwؾ�5�W�A����imZ�¹�>P/^}c5w��^I�P��y�������U������'������_�~�°囹��J7s޺?��
�Ϥ�el�R.��!H��R��E8�R1��M�$���U�Y$I�$IŰ�6�����d�}�x<��_��_uI�8��-�opv���IE�z�� �IoD[�d� �u���K�UR��N�$������0aB�1�⢋.b�v�:�$���625\l��������5	�^�]�1�a�63WP��H�$I�zu�i�E�l���9��S��!I��n�,��V���p|�'��� � >V�XQH��z p
����AQǓԳD"A<����A�
���C�Ų�1W�04�9�X��[f\��:;���O�$�?6lcƌ�:FYM�4)���~hp3P��KE�a� �g;���{8�P[l<	�q�v}��೟����X��n���X��J$<��ω�r��TIo��:�>�-y+��$IU���#�e���uU���_W%�Y�{u��1≺�������ϋ��8��,Y�����DN�n�������������01��������/��=H۷���f`:��+g�jӸq��m���2W��s��g�$I%�����/�\��v���FAh��Nf�aQ���n{��aBss3�_���I�*�CD�@қ����I}���Ǩ�b�c��]�"դT*uI�$ՠk��&�e�t�Rn����c�YP�T*�I�)��޽�Ї���62#�����������̂-u$I���u�]ǽ��u�������3Ϥ��9�(�D�{TI�D�j�����CT���0�1h���[��DO($Uu���*� RM���Y,�k�$I��H�R�|����'?�ٞ�s���c���:�*���d�/LRn�!��e*pZ��y�p���G����FD��{�/��$�
%�q���#�6������1nܸ�_}��\{�5���W���T*Egg'����X��0�q��8�����˗s���S? �f��0{����FY�Rn,�K*�K�e9w�uI����@>���|�x���)�7�_ED�	�{�oǒ$�
��0�l�-[����,`�m������&���ʔ�<��z��b�˗/��vc��e����i����RFR��u�ʴp2pk�9�ÏЯ���x���g�a��9�1�/��r�A�����ǩA� �(�k�:S���C�*Ez��[�H}�︺��p[ ����Pp��@}irU��z�#���*�T,�g�(����(N�䔒ϳ�v��y��S�!��������
���?肂��=Jl�͙�6�m�ߥ�9z�_`�����T\�׳jo-%Ee���CT�=�ÁG6�`.+���.A�*����k��,_ԥ�Yp���I�nȐ��1i���3b`C��x�������Pw�u	��x�n��K��1��9%[�*�W������Y�N��{��Y8��ty������CHU͂{/\�"I�$� ��홋���9=� ��o��l+��V�<�f+�"���"U-��$ͺ!�&��X*st��Gg���1�w�/�$�({��̂����̙L�:Du|�M6O����,y���U�+�ED�J�3���]��&E�*��D*���aY�T"ܥ��|0���X6)���[���R3i Ή:�T�,�g�/��$I�$������#T��6}���n|�a��7I�����i�����%I�$�뭞��I�S{;�瞋:E5�>�]7<ɴ����-3�u�*��$I�$���[=��.���硵5�������~F��T1�DR_$�ɨ#T,{�J�$I*��$��G��}h�z�45�8��a��a,X�����!U{�g�Yp�$I�c��8���O���ʵ	Z]y���Ç3v�XF���������z�B����aΜ�T����C����*`ڴ�	)/��腷9J��2v�=�q��>�>S��S�r�Yg}�j��~�q�y�l�'����������zKRQXp�^�G�1HU{��QG���̙3����������ǒ�$����R��5j;N��ᛌ�A*�y�:;[!�_P���e='�J�ޞ��$�줫�m���Yϗ$I��L°|w!�RI�����%�S�[�vt�/����I�R�aȺu�_sutt��޾��a�����ԝ�ٳI���w�NP�&l�C��{� -o����3H&!�:�T=^z�%^z饒�1n�Xv�V�9$I�$�Ҽ�����V�%;۳��
�$��W����Gyk�;tuu���iR��]u�j4 �� :��
�"Q5jl���p�Q'�$I�$I�]5�5���Jss��jں�w��GC���w��'�$լ�u%I�$I�$�|,���Pز���NT/��!�	�$I�ԯ<�q��1j�(�����Y�p!K�,��Ͷw�$���!�B_�-�"R�f����;�K�$�'kC���std߿[E��?'�p�<�'O��T*Ō3��뮻��m��$IR��z�&ز�[A��ܹQ'�$IR5jY�~��|����G?��h�sc�|0|0W\q=��{n�7��$I��С���	�{���j+WF�@Җl�$I�Jk����{�<���9�{����3gr��2x��"'�$I�!C�NP�B�6[��_�<55E�@Rwa�ࣳ��QQ֬��iI�KC�4B�{<�������2'R�k.�������2�)��ɓ��{�q�+��}�)S�p�	'��;�PR�jni�Z����d�$u7r$��V�)�ͪ R�yK��@<�<ի�::����9I�����:�$)B��x��n��$�����P����2���;��o���+�'O�����9��cm1#հ�u�^�t3n\u��K����3�D���lܜgӖ2���G��E�@�$IR���^�v�m%k�2j�(��F�U��%I�r2qb�	��Ƃ��+�;"R�N I�T��yo)���_J>�A{63u��+"b��H�M��4�]��a��T����4�_�׬���Z�f<��;k�����{�/+��G���w��СC���g;�w�qGu����fG�$��}�c�}����6��x�:�$IR�kjj��W�|�1Ca���xV�[�<�M�d���Yw�+������J:G!~����N;�e�C=����+�(�|��fei�@y��ż�꼒�]��y�~��p�a{SWW�n��dg�ǔ$U�}��:A5ڸA�&� 	a+0(�@Uk�|�B�$��;u
��^{��駟^�9�?�|~��߲r�ʲ��a��A�����[�}�i����O��{�Q���ٛo�ɴi���(˜-�ޅ�a?�]L�&;�D����H��� 6nБ�vp-��2lX�	$I�$�����Ų�XDÆ��/���nY����$�����:g}}}Y�&?����� I�ɏ~���\�`����w�1e�S��tW�$U�T*Uйa�ti枾=���Ǝ����ێe�m��5F.֮^��6>_�t�^)~;���m�>�w��|��A��~Ϣ����ʢ�_��<�L1���>O{�~�}l���I$�_Y���tv~����rUSΟ���������N&�9�+���3�O|�}�ܦ�&V�X��ѣ؇>�g�y&�����������$I}�:�p�ӟ��Q-��I������e�~�! ��[�dI��.^�8�9�;rO>`���;�v;�~P^c���y�1o�S�?�B'��_�\��n�f��ö���_*�<�M+���Ivtt��/�<�xl����G��!E��G;hmY������~���ŋ>|x����I�����{u��iӸ�K�>}:a�H$8������O�ͣ'���Ù:u*�=�X��%I�
���'h�Ӥ��ݹ��9�Ay��.��{��r>wڴi%L"O�߫�����7�,qIQ:��:�ꫯ���g��ؗ��������r�!�{�%�_�$�­�澨CT��xy�t/�G��>=���'�x�G}4�yw�}7�f��z�T	���*��w饗�їT���{�ϝ>}:�sN�ׅ��6N;�4-Z����O��J�$ӍQ�[|��ܟroZ��%p�!Q���]QG�wN;�4�x㍌�_|�E��կ�1�T����/|�{����?����}�BI*�x<ΨQ�r>��?�q�= �����krs�ر9�+I�TL��o�ZS:�-v+�VpV�m	�2�<�����:�$Eo���L�2�+���e˖m���E����K�:u*+W��0�����������q����7fÐ��SO=���>;ℒJm��#��|�O<��y�?�x�cZp�$IQ��'����A�It�4һ�z�b=���:��n\����&.��.��ƍG*�*��R��x�N>�d���?~<+W�̩Ռ��0dH~�=777�t޺u벟�ޠA���bYW�K�$��/��Q�<I��=��R�o��R;?�-��z`�=z.�خ��������-�K��ҥK�:�w��]v�%�1�-[f�]�$E��:���� ���@O+� �K����~{�$I�ʣ�ֵD�B�jk�:��innf���9�ꩧ��+�d=���|���`U�$�~|�1� ���A��=܃�� �V�L��Fb��:����]����f�R1���{|�C���s�9��o��׍ď>�hN>���$I�R�B�mQ�?`~��=���c��Ԑ?E@�$IR�=���9�;d��M�Ɣ)Sz<~�	'p���8 ��%I�r�aޟ���ŏR��$�^�=���W!|8���j�_�9Q����+�%IR��u�]|�;����������Os�}�1m�4�/_����9���9���;C���|#K�$��Y����Q�N'pf �6C�Pp�?�����9�ٗw�$I�$U�'�x�+V0bĈ�?'�q���s���4���>�C�$���.T|8��K/
��l'ej)� O1P�xx2��z�
wI�T,]]]\y啑�}�e�E2�$IR&�WG"���?6�^
� \Rp������$I�j��W_]��K�x�	�ﾲ�)I����:Dy�����Y��R����S
�U�<uIYA���u��2s�<�66GC�����������7�\��:;;��w�[���!��>V��^zu>s�Z\���ͩ��J}]�K�"�;o�Μ[��jŠ�8���QǨ(��Yu��)�v�9�Q`�b�l�O��U.?�����k���|/��r��?��e>�ނ��%I*�-��)S8��K>�w���{�S,�x���p��[��ق{/��֗e�,��i�����U5���:��>h>I���ng)�U�1�u�c��2@��� ��R'U{�K��R8��s�6mZI���/ɯ���!I�Tˀ���R���x=�O̡��π���v��K�T-��x�$IR�����O�;�(���^{-�sNIƖ$I*�%��\�y�G�>���cc� �����2Q�z�r�/�����NF�$�Dss3��r
�w�_~9�X�k�2�������&7�pCV����g��c�>�Ǐ��1{2kV���룝vډc�=�]&~����/@Y��,��΢�+I�~kH�#��R�Y��Q�� V�u�<vR	VC�%қ�6�u����D�]O���B*��Fauur8-�0������$IRA�0�G?�O>�$W^y%�rH�Ǻ뮻����={vV��#'��.}�]&�GZ�Yg�U���ٮ��ʹ�[�����wIRFm�i����A�����(�d!�uy�4�����s�M8x>� RM�0ag�y&���m�TWWGCC���/9�޸�,�SWWǐ!C�t�}��-Ǐ��c�W��uA��j�Ā������/��5v�$I5쩧���C��O���&�vuuuY?����iӦ������z�I%�A#��~��b���_���������K���#c��� [��&4��|^,���隣�1���
�G�}Xn��8K��C��E���~S� �)����B[�H�6lg�qF�1*�7�H�T���N��N��f>��O2e�Ə��ѣ1bK�.eѢE,X����iӦ���ulI5h�]`�}��&
��Se�g���ܥ2y���C`h�qz���8���@�q�zp-�[�^f_c%���]�$I�$)7�W�榛n⦛n�:�$��\�@�T<���H/g�8(|盢z�� ^)���=�g���Ո.��H;H*���Eml$I�$)��2��.E�=��������{8$��KQl���XnN��&Z�O7DDR?��C�$I�T!,�K��͹y�xO.']�/��/�}�ڟ)�dEXN�@��(�7��I�+IѰ��$I��¸�=�Rex��	8�-0�4S-nN ��� ^*�T��c���N��^�1��F��-Q��oq�̯�$I��Bx��Y"Q����H�� ��_��H���LF�8�Z`��ǳ�#�^̼�(�M�
|�H޷/�إ�p6pO�9��%�LF�b�p�$I�T ����#H#��[�_�� �'�  �m��!�C�j&�|�0��e�۫���	�߀�����Q�N�W�o^XW���a'm΂{f���N�$I�j�w���������~����?�gy��p%%�ԃJ|�H�R*��:B�����::Zh^W����ѴK%�hj\^�q[��}�\�4�������B_S$I�>ࢿL,�Kp�pi���U��O�p.�e`�����j���O���Z�,��Ƃ{_-|�e��r�1��y�*�{⦨cՋ��:�$IRͳ���+��o    IDATwI�R���������(�2����C���x�_��.U[�d�1�$I�
a�=3�ʥ�[4����G88���Ǿ���pw 7�.��.8���s��$IR��x��YU��O3f�e�s��>n��5k_����ڙ�R__�K�ή����R���I"Q���~+�W�`���C���``"��������.� M�w:m$�d}07�ߠ�ة\I�����+�%IR-iY������+/��3/��{}�j�|�r�}�YN8fW�x5��bej� �߫����f���I5ʖ2���.I�$��l)��+�%��o�I*+W�K�$IR�Xp����ŷ�$�UWWW�*�-e$IR5��Jq۟�(�|��/)�\���{�&�(Oaq���e�G��ទ�[��ł������:B��@I�T�R�=�RY笯�Gy&�ը#H�T�8�#�=>'cH��0�tǖf`�>����s6�6�Y�ț��^b�O�6����^��.I�$� � $U�	�߁� }��<�����|YYp�TV��/�����1k��0Y�vm�7�:;;inN��~�#��{ަ"�tue/���$�d��R�.R���vuu��{�wv�gC�$I�2��E�d�T�:0���>A{���H���m��U�V�L�~M�v�ھ��jP��VLX�(Dp���y@0�#p���%g�]RY�R)�>����S_�8�$I����+�c֌;��~6�e�O�H�h)��"��o߮���$��Y@*�ڸkC�=CےJ*D=��������J9�wI5�v�$I�����f����=� k�6�bŊ�cH�}#�����!�f)&�߂$I�$I�$I��8x�0��T�
�0d00
ؚ��j�]h�-�$�]�2[E,�QWW��9�x�Db�\�y�{^<���1�ϑ$I�$նrUM���6^oz�H$6{A�����v}��H$A��EN���ݯ�7�p^,#�y�l*�"C���[��R��	��q���2^�A������sK�M�^anqަcl�L&7��d��uvvn��?~<�����o$��pppW������ٻ��}�㟙���P��A�����""(Q��rD�r��Q��稨�ׂ^�X ł�"�E�tI(�'$@�df��ȁ�ԙ=�g&�����g�>��L��^�0T_R?I=$���RR���k��I�)i���-[*r�Wnp��.B�U�cg�ץ�)IEo&gޜJ{����t�=�0��<?CIǕ�r�u%�)���̛NYu


��7X�~}?~���ar�\�9����~)0��     g$&&����%.���������q����?�F��KzO�_U4��#>/��l�.�t��
�-�lʦ�oH#I�%ݽs��}��d���GҊ݂M\\�RRR��T���}:✋P     ���'���J�&�I�<i�gs������G�RI�~��T�[Kw�)-_.��-=��԰�ٽ�*��>~�    �3�������R�5�4��f��4����iS�Ǥ��]��ciڴ�� �㫂��u�bg�3N��VF   �j9���e�V�c��BǅӴ�+Z�<M/�;x� nj,�YI#�Ñ�%	�Ǝ�ƌ)*�O�*8`e"��7,T�ǟ//q~�3"##e�ۙS   �Ϝ<��w?Zbu�8��Znnn��%%%�"�� ��>"�5I	�fT�d�ᆡ0��I�%��F�ۥ��oiǎ��f�íNTMe-��mݻwײe�t��i�:uJk֬�W\aY    &={�����u��)�>}Z+W�T߾}��� @�>f�4]�=�=��b�a���&��))�̶�]4����RǎV���r�|ާ����p%�{��e˖��.SHH��v��u���NC��z&    f�]v��.]�޽{���u�%�h���0`���|������"�IU�L�z�n��&�]$�Z%M�buT/�����/���"##/��Y�f��B     ��_~Y�%L'�ٳg[z�3 ��.�]I}*z��s���I�?I�{ږ"#��3�=�[o�ʙZ�	�(l׬YSݺu+��F��m۶ڲe�S  �����YX��Y_�(""L6���Y�t���Y���W�J}�y��j޼�v����T��?CX(Bҧ�:I:\���C�J��I;�`�h�iS骫��t�Ӡ4��+
�			�  ����C�ҳ����/�Y�~���ͳ���(�\ Y�b�>�d�O����3Wq�/����#�I$�y��킻a���E�ڻۆ���C��gi� i�~s��� �Ί�L�  ���V�:�Lo7�^O]zY�>��S��d:t�}�ݧN�*$��߷�oZ���|�� ��J���t��g�:ȭ��a����ko�����m[i�R�W/�p�7��xA��  ���&�v���[��T�^c
��S����wn��km��������O<���eRJ;�җ�C�%}� ,��Ѵ����R|��I �c�;      P!Q�f�u@��^��(�;z* �o/͛'EDX���jfp��wF�     �KZڃ�f���`�Ԋ����^x��8w     PY�?C���$�8ڳ�w��hI�L
0��Wi��S�^\��r�|�'��    ���������t�4��*�h�a���7�LH^yEZ�Fڵ��$���$}2�}��j���_��J����Ճ��㕶���T��e�󑤓�r,�    P�<���׋)��n�K�#��B��8i��o_�z��(�F��S�9y��ɳ:�i�Be�8euS��  @`��������VlD`E��� ��7�>}�Z���j>+���    ��������O�=G�w�P��i^�`��o�F�STm��    �ʢ� ��0�hI��(o��#�jy-N��SG�:����S�<����^NT����    �%>�>jB�*���~�z%	x	����Ԃ�a(Q�m�Nh�S��/����e/�W��<^\���     s�Y�||O͵jժ2��}�$(>���F��+)ƻYO\�t��E�gJ��������a����rY&`d     �5l6��l٢�?����

4o�<�
h����Ă�a(F�$��	@S�H��Ҷm�4d�����}�0}��5j��	�W3����R�     xP2ϙ�孷ު����+6�����6l�������ZJJ>�Eh)]/��AK�� &}�����?�e˖�֭�����a����Z1h9�N�#ް   ���Vkߟ���������jР��m��K�j�ܹz�[nz�G��m���AY|�F ���������#���/VFF�V�^��������>�J/���]��t�]Ք����:t CI�"�T����N#B�"bP��}  ���B9��������S�N��n�s8��ʒ� O�!Lŉ���4�����<aa���[�b���.I�ұ���ҟ)����ڞ��w�P}U�Q�����{)''���V�߫��6�(U�+,4���.X��     ��nWXXX�ǅ��(4�±�����}�7���Bxxx�����}��~_hh(Ӝ�$:*Bn�_����J����^�(i����B|�%0��.5j�G۶\du�*Ū�{xxx���e>n�l6[����v�����5��q6�����v�bcc��+���r)$���ùw���'��n�a*,,���Tfff�y    0K^^�J}��r���^��?O�l6�l���g��V����r8�~;ӟar8�g��ʝ�#?��)�


=�b�n�2��J؇�kp�����\��WH�S^���r�U�7��7����     ��>}��@�8�q����陿+��B$��y� U���l���1|��7��C�ƴ5      *�\jjn��&�q���$��>O`���S|bF�Q�       ��)��)F��/�w� H@�Y��       ���សW��(S�ta��U	���YD       @�(}JÐ�.���H����jğ(� y       l6),,��Q��҅��	h�p      (�rFGD��(I�9%]Xp�eA���ku       ��rf䈌�M��bHʖ�����}��^����ҧD   ��WX�҂�W�������t:u�СR�INNV˖-�\�t�������-y�W^^�$���*,,�'���?�~  �S-RǎgY#�dJrJ��CQ�� �r��8e���r��     ?�˥o�_��~�9r�������;:t�����ɓ'u�=����.��~���D �`T�V���}e�y�/������EZ |b̨�R�K�Z�o��}��|�{�c���wZ�����_j��V�  xYdd�~��u����(^���zKv�]s�̱:  `�=�LR�>�Tv��˹w�A������ T�����&�nWHw�����d%;� P%���A]l?�̙3��_����VG �:�㭎�J,��� H�3�V�    +M�0��>�n�A�g϶:
���Hկ_�g��8qB999>��GF9��&�O�M����_��m6�r%EY)@Ql*�A�r�\>��r�(��n�  ����M�Zç:t�`u�{���i��գ��#�v�jT��̬l���BI?����ERO��{�8
­� �˥��4�c    Uf`G���� `��olټ�֬�Y����u*��K�Ο�u�o��ӧb��  @v�]�_��͛�#G��09�رC�f�R��� @������ݻ���S�6m*�   �ԺE��ɒs�8��vI�|�%�ef��  X�f�+4����\�.�\�O_��ڵ*uNӦM���K�ڵ;�/�D�4Huj��M�=ZcFߨ�s�j�����˫T�6ó��B��n/<l�P�#ߣ� pǜ9s��3�X�'N�:�O>��� �@U�)|;^�Dv��;�*f��_�_p�!TJ�VG �*�f�fj��b��Hr�8,IK��L�W.�(˨��+}�ܗfT�kzT~~��+<��o��U�I3��w:t��n��\�ܜ,��  PQ/�������+��H���w߭��t��  �Xll�ڵn��[}��B �%i�;ΟRf�����pw�O
������_���u���BBÔT�����	��� �"���5p�@͛7��(^s��	�;V���Q  ��%I�tk�� ��7��G����y�^T�a�t�p]�c @�R�~k5l�������p��:T���#��r��  ����L�1B;vԠA�ԨQ#���X�#�C'O����۵`��<y���  0A��MT-:R�9|�+�S����,Vp��t�0�MR[_�
d�k*/7�� P�4mq��P	a�QJn�I);WYUXXX�bbb���[�5 ��7j�ƍV�  �OUl�{XX�.����Z�������%]0���S�H�O����W`�^��� �'*:NQ�X;#��'6�:����=�����ߔ�����eggk�Νz��Ըqc�#   ~nudH�^�%ܿ�n��q`_C�# @�mu�!"���P��x�ڽ{��z�)u��Yaaa�$�ݮ-Z���ӎ;�����u    �2T���e��Y�͗���Ο�]�I:.��7�ܜh:�Bp �K�?7福����~�>��O�tvŦ����{��sϕ��.<<\O?���7o�[o�UFV�
U���
�t�!����   ���N�1�W��z[�'�
$=Rڃ|J���0},�.o�
t�����U�   �w���j�\��>��GK�b��r�0`����W�"����e�=����[/)A�T��d.�K�}��@�����
] �W�EGj��=����D��I�Vڃ�U���N��{{�
Ǡ>   �լY�d�W~@�?��O%%%y! ��n�몫��o����(##Cڿ���}]��g�� �4n\��}I[5m��̒�Kz��J�Db�i��_��(9����̸  �/�-Z�unLL�&L�`r" (]�����o�髯��_��5n��la=44T���3f�>��SmٲEÇ�81 ����l{��
��Z��%�6I�eT����	"���nu   �c����?h� �� @�l6��N��E��cǎ:�e˖�7o�^{�5F� ,U�n�n���V�!��*��P�&����c�t`oC�c �E �Ժuk��oӦ�II �t/����O����W��~���}~� X�O�vj׺J�FWIz�"�z��&�0�OI���*�[���   ~%,<Ru�V\�:
���Q[��Ѯ�/�o@�>����2����7ڼ�{��~t�_�|�n��DZ�}I��M׮��(���S�u$m��rOz� �5q�DM�4ɣ6F��-[���'�4) �*�ti���:���L� �I!�Q��˜t�f�<�з�<�G7H���P�R[  �o�Jj�6�+4,���LUZJJ���:zȔ��s⼯��k)���#|ꨕ���Dn_��)�y� �R�N=�쳦��裏꣏>��ݻMi PyXq�Z�K$�`EO��}l�%幛(X�j����:  ��H��PubZ�����CԢ�ejи��Q ���Vll�)m���1� ���1�UF��k$m��I��m6��jÚn:�gu   �`��Ժ���*?1�֬uo�GD[�IBBB4z�hS�>|�i|  P�L�l���'V��S�~�l���PZ}m\���   ~�z|=EFW�:FP����VRs�c 0I�^�T�fMSی�����Mm P�0��<�$].�gwN�P��fS��ђ���I ;u*BK�a�<  �1���P�_ x�m�6�� ���$�����m��� �l: �INw;4���;ovVNv5�� �f� {H�Z(�����#))��Ǻ\�
[�^=w�   ����=��z�H�&ݴ��;=�0P�t����.    ��n���nèx�-  ��r�,Ic$�,)���*=t�f�놡$I���s��C�[oIw�nu    @�:t�P��		��iii��,5i�$>����������2x���T4�|�Y�u��ͦ'C�%�gV2cF�    �'�n��v�m��vo;v����oZ��,i����n�RSʜ�f����QM�c҃m     x�_~����Mm3??_�}���m PElT�:���b����3l6�h:)�uO۲��!M� ����I��Q�c��ý�   �_N�S����.�����/u��I���(����~�8qB5j�(�؈�S�Wxxx��s(Ihh����=�����bkG����t-����+2̩�]�v�!6)�׿��P�ݜ�!!��}pS����yC�ׯX{\$����ah���$��<����/�-�Xa~�-���-7]c~��ɐݤ�tV���yk���?Vl��oXf9���t��tZ��f�y�fw�|��!��eb�"�6�M    <���7n�bbb<n���P�>��	� s%%%Y�B&N�hu��Y�fJ���j%DY�#Oү��J�T�	_ulʨt�M�C�$�#i�m��W_I��I���i?�F�zuk�ƫ��;��ԂC    �>�|P�f�򸭧�zJ;v�0!`��;wZA�쩹��6H�'���V�K��j↊=�)i��%**�皞�L��f�q��P�������ͱPF���C�o�ݎ�ҫW/=����ݻ�"##��    e�={�:t��o���6�ϟ�'�x��T�yv�ڥ��t%&&ZA&--M+V�P�v�����RQM��I-$ՓT]R���OI��ϟGTTh��eز�:��&C�l��ǒ�I�M�_�sbE����HG�Z��2d��������    ���'jϞ=z�g*=�믿���[#���n��}���~3�+_^^�ƍ��������%m��P�R��ٔ.���ےQ�43��CZ�Pz�Ii�:+�����z��(��+|��   ��04c�m޼Y��׿Զm�r�ٳg�|�A}��>Hx����E    IDATT�Ν���U�V������Sff�
��� �p8�f�͘1C���q�J�j��f�*ICC�%=$�ZIa���|Ҽy�3�H�6��gxC�.]���lu��Yo   ���7����5�\�뮻N���Sݺu� 9r䈖-[����?gd'ʦM�ԩS'�c �e|2L�f�I�C	���t��^��s�V��w���f�`cu1n{  ��8�N͟?_��ϗ$���)!!A'N��� @ ��6�2$�.�u�PsIWH�'�rI�<l�ȏ?�1w��/�RR<l~i�ƍ*,,dJxŢE���   �*��p�ȑ#V�   ��ji�i��ݒ^3�$5��RR���YOE+�Ʃh%Z�h�ړ�NKJS�
����gʕW�3I�7����5{�lM�2��(2���p      ��&l�ɐ���o-�?����M�����ۘ�ذa�.��r�c       ��E���á�'j�����K�����*''G�����ի��     � @�+55U���V�        I�q        `
�        ���;        &��       �	(�       `
�        ���;        &��       �	(�       `
�        � �� �.u�Q�l6�c@R��SVG      �2Ofk�ֽVǀ��C�VG�k�˱p��#       Uڮ?jן����)e        0w        L@�   �f��    ��Pp  @�9�VGj���   @ ��  �J��`�*o:�~��    �@�   �����c�w[#(e��PƱT�c    pw   �e��%��δ:FPq8��ǆo�#   P�V �@�ի):*B��E/�����Wff�
�N��o�hݯsղm_ծ�R6c9<�q|�vnY�.b    ��; ��n��Ar-�n����nR��ce��J<��2��qRghן�cW������HE ��Q��?~_��,Ul�:
���|G��]Ҿؾ�;���2�5j������P���J����F�{���EE۴巯��W�\.�N�<���S�   �z����%���սkKU��V���v�jլ�Z5���EM$I�Y�Z�n�V�ݡ�C�ފ �r8�ql�)m���uݦߴb��2�{�_�늁n��o�>}��7eӸam��^�ؾ����;t��~   
� p��M�jЕ]վmc�J�^i5�W��+�h�]�{�!}��jm�y��� ��u��i�С�    �b�M �T�fuM�x��2BڙWl?_�uuߤku��CU+1�;� @4w�\��;w��i    TU�pP��l6�����Maa!>�C��j�2Y��w?n�H ��o߮y��iĈ�>w۶m�?�R   �j(���bc�4��jצ�%����꺫/U�V��{����Kr L��fu���ͯ�q�'O֥�^��u�����kܸqr8��(t���
�ȜN��   ��D�@��T'^���%��ZE�[&�{G��W���'�� @�:��>���j������*Tt���ըQ��f͚
��v0]�<���1   1�pP�4iTGS����b��	�z��jܰ��Q����:����ڼy�:u�?�P.W飴��'u��U_}���   v�pP��KJ��W�Zt��Q.S-R��y�����:p0��8~)/��%���Ł$7�jL��q��Q�3F���?t�תK�.�]��233�e�-\�P�����1   !
� ����X�s�0�,�����Z3^�L'2O[��8yJ?�W5k7�:
*�衝VG@���瞳:   �*�!� ����n7P5�W�:J�j�h��
	�%�$��-������2����V�     �'�� �F\s��6N�:F�5iTG�^u��1�R����f����ߥK���_�0��     �L) �5nX[W��hu�JЯ�~���R��:���:qH+�����o��	��v[�a�۰���:��ϯ��{�ͦ�����U�������U*���&��g)��>��5�rs�t��n�    @��� ���6�t���lVG�4�ͦ��W�<��\.F���,Tھ�J۷��������起U꜐��{�z�����X�1�����L�����ҙ^�J�s��?����	     �$
� �Z��m�0���1�֨Am���J+�n�:
L�t:���[������={�A�*((�Ν;�x�b�\���X     0�-�ݦAWt�:����U�vP|B��������g�Y     ��ES�.��N�V��XR�xuj���      (w A��%m��`�K{��:      �A�@P�Q��ڴl`uӴo�Hq��V�      @��@P�xQ��6�c��n��}��Z�j��Q�k�Aق�{�ԽG��p���Y����ʶ:    ���� (�n�luӵnQ�/
�+�l��5ۭ��2���VG     �JbJ A�e��VG0]0^D      &���q�eu�U����j�V�      @)(�:I�kX�k���[      ��� �ԬY��^S+��     @��� �DG�[�k��"��      �RPpt"#���fu      ���;���/ma�!VG      @)��*���/pX�k����     :
� �N~���
��      �RPpt�N�X�k���     :
� �Α�'���5���      w A�ȱ,�\��1L�r�t��I�c      ����P�:��R�U��iu      ���;���}��#�n���{N      ���;���u�>�#�n���VG      @(�J�wP��l�c�&3+[���:      �ju �L			�Y���nիWWTT�$)..N!!!���
W^^�$)++K.�KN�S���JOO�`s8V>5T��eh����yg���b���A�,     p�������jԨ���P�l6ըQC�!�ө��B�\.eeeI���򔕕uA�����[�Uw�5j袋.RӦMդI5n��얜���P���>z��RSS������Գ߶m�����K����uEߎ���f�ӥ����    �* 99Ym۶���Ҹqc%%%y�_�ө���b5�3ۖ-[���ᵾ3٬`��%]gu��e˖�ܹ�:v���۫C�jذ�ձJ����M�6i���ڴi�6nܨ6�����hUޭc���ŭ�������:     �����cǎ�ܹ�ڷo���۫cǎJHH�:Z�8p��y�fmذA۶m�ap7x�X*�r�C���;��޽{�W�^�۷�j׮mu,�8mڴI+V��/����K��رcVǪr���뱩�����z��u�x��Q     ,66V=z�P�޽յkW���GիW�:�GN�:�իW����X�B���Vǂ{����_��@ڶm�A�i����ӧ�"""���U�ahӦMZ�h�-Z�+V0/�����R����1���wk��7���    0�����K4x�`4H�:u
�)W�SPP�+V���lڴ��H������(�����p0@C�ՠA�ԨQ#�#Y��ɓ������j���,�E�az���VbB��Q*�X�I�s��*((�:
      ���kذa2d����vӪ*--M�-�W_}�E�)//��H(�RQp�K��LHH�z�쩑#Gj��ѪU��Ց����ԪU��駟꣏>�ѣG��t�4���M�N�!!VG��ӥ�4O{R[    �Ǣ��u�UW��oրnu$�����%K���w�՗_~���|�#������(���K.�D�Ǐ׈#���hu��RPP�ŋ�w�тXx�D�u���zY�B>��\K�m�:    ����i�С7n�����-33S,�[o���˗[E����_��n��ի�n�_��Wu����8A!33S�|�f͚�͛7['(�x]�����eZ��}��R�c     �Lrr�ƌ�I�&�A�V�	
;w��[o����~���T��w\|�Ś<y����zEEEY'h-_�\���>��32����v�n�e��vjnu���m��|�{�au    ������ku�w�_�~�ق������`�����Z�b��q������(����nW�~�4e�:��8UʡC����k�̙��̴:N@��m3�ԧg;�����mz���r���    �XDD�n��=��Cjݺ��q���~�M/���>��C=��RQp�Kܽ,22R��r���^�j���8�r�\JOOWzz��?���<(;;[����������K����U�Z5���(11Q5k�Tbb�_ρ�����_]/�����Ҭ�pl6i��:����З߮��߭�4    �zu����ɓ5q�D%$$X�Tg�.���*,,TNN���H������IE��FDD(22R���g���+�F���٣�3gjΜ9��ɱ:N�[*
�~�������k	z�ᇕ��lueeei۶mJIIQjj��m߾}:v����M�'&&F5k�Trr�7n\lkٲ�_̗�����^{MӧO��Ç��pZ�L�_�P\\�%��:�����Al�gI�     �P�fM=���4i������z��jǎ��.)))JKKӱc�t��)S�IHHP�Z�ԠA�bu�&M��M�6gKZ���Ú>}�^{�5���Y'X-w�D��d�������裏�q�ƖdHII�ڵk�q�Fm޼Y�7oVjj�%Y��:�}���С��v�:(44��Yrrr4{�l=��:~����dqq�9���wm%_v7i������:u*�7�    �N||���~M�<Y���>���tj���Z�~�ٺ�ƍM�����t��Q]�vU�-,�r��M�6Ms��QAA�%��RQp�K�Mt���kڴi>}+,,����r�J���/���_u��!��o�jժ�{���ݻ�z��^�z)..�g��:uJ�?���}�Ynw��V��k��=մq�W�ٽ��-�U��ֿm    �y"##u���P�5|���ӧ�r�J�X�B����V�Ze�hu_�S��z��y��ҭ[7��������T=��#���e���rKE��/Qp7A�Ν��/�o߾>���ѣZ�l����+-\�P'N��I���N�:�ꫯ�СCեK������'�xBo��&�pVR���yg�k�Pv�9?+�˥-����%�s7s�   @Uv��Wk�̙jڴ�O�۳g�ٺ�����γ,���u饗�ꫯְa�ԨQ#���n�:�s�=Z�b�O�rKE��/Qp�@�:u��O��[o��n�j_[�n�'�|�h�ƍ^���ԭ[WC��ȑ#կ_?�/�r�J�s�=Z�f�W�	Fqq��ޥ�ڷm��M�*,�rSjw�!m�#Ukۥ����     ��N�:i�̙^��r����?�O>�u�����oڵk�aÆiԨQ�ر�W�2C���z�!��1��KE��/Qpw��n�wܡg�yFիW�Z?;w��ܹs��'�h˖-^�'�ԪUK#F�ШQ�Էo_�]�0Cs������7effz��`��k�^R��Ԯ���XEEE(2�薵�|�rr�u"��ԡ#J�wT��N��    ��iӦ��;���g�˥_�Us����pS�zK�֭5j�(�5J�ڵ�Z?���z��G��K/�����
��{��\��V�y��ƒ%Ko���5>����+�4l6���ן�z��S�N5RRR���8t�q��7[�\�������������ت�6x�`c�޽^��?}�t�Y�f�?Wߺv�j���FFF��~6l0�v�j�s��'	F�WQaaa�:u�y�EDD���ƍ����>PVV���&**\	5bU�Z�b�E*&&J1�"��P��ËF#���*4$D9�Es�9�N���QX���<�>���U��e����s		ѠA�t�m�i�С^�rf����뮻t��A��  ��F�������TAA�O?+KTT��W�����8q�E�  A�v�ښ9s�F�mz�.�K�-�o�����J�����Q���hU��VlL�bb�T-��ZTo	-�cDE��p��wH*�v��Щ��N��թӹE5��<�8q�l��bbbt�7���oW�n�Lo��p��g��SO=���<��RK$#�)�WA�ڵ�|`�V�a��o��s�=�%K�������BT�N����T���L�S��8%&ĪZt�W�t8�J�8��S:�qR���Pڡt�O;��l�p6m�TS�Lф	cjۙ���4i�>��CS�P1�k��e�]����+11Qaaa����Ν;�z�jmذ��Ν;k����eggk֬Yވ.I2d�ڷo_lߢE��ܺ�?����5�\�~���{��jѢ��U�V�ӧOkϞ=Z�v�~��'-\�P'O��j��ի몫�ҕW^��;�]�v�8z��6lؠիWk��ڰa���M�:���999z���n�J:t���۷j�*-[����n��6%$$۷p�BmݺՔ\M�6�ȑ#��[�x�֯__l_LL�&M�dJ��a�sE�����k��f͚������w�}W/���v��aj�犎�P�z�J����I	JL�S̈́X�L����f�����SJ�8���'u�p�����*(���޽{���Ӱa�L��g۶m�馛��o���n�Z*
�~��{l6�&M��g�}VQQQ��������{O/����\��6%׫�fM�Y�$5H��:��{}Q�����ց��ڳ��v�9���G�����f����wܡɓ'�nݺ����hҤI~3�v�{��ԩSu�UW�f+�m855U�f��+������2�lҤ�v��}�k�E]�?��Ô����JMMU���s:�jҤ����oz *�N�:z��t�m�)66�R����꣏>�3�<�ݻw���cǎz��u�u�)<<�R�[�N3f��g�}V�~Ͽhy��1ծ]��� Uѭ�ު7�|�ؾ�ӧ롇*�;v�e˖��mݺU]�v5e��!C���_�7y��.�իWϒ�ǌÀ&�Z�j�9s��򗿘��ѣG5{�l���:v옩m����q�:j޴��6NRr�D%�W�w	o2Cǎgi߁��3��L9�}���r��O�-t���[nQtt�i���Gտ��o�3�����(���v��z��7u��W�֦������{L)))��i�I��R�6պE��4��Ȉ�}0����ҁ��ڹ���ضW;�<(�Ü+����7n��qS�����رc���?��&��"##5c��}��e�ϗ���[n������/�W\Ql_E>���+��?�Pl߷�~�!C�����9r�^{�5���{�NAA��q͘1���gn����+��W�o��Vw�qG�.�Qp�gf�]��~�i=��#��w���>(�������5k�,=���ݍ���]�jѬ�&�RH��l����R���]i�c�^��̴��jժ���_�'O6u��O?���o�Y0�� �TARp��= �+������o����B���{z��'M)�GD��C�ƺ�m#�k�Pqq�]E���nW��Zj�\KW�WG9�ڹ��6o۫���(=��m��ҤIz������q�jɒ%z�'��SOq�0YDD�,X��V��ƍ���رc����zܜ9s.(��=Z?�����o��������L�<Y3g����-]ܟ6m�ڷo�[n�E�{w�2D���)��H�����j�*2���� 4u�T}��Z�v��Q ���l����=���
3����L=���9s�N�r��pF���ԩ}Ӣ�-�nNN�D���U�d�j��aCz���\mݾO[��Ӧ?R��[�v�ǎӃ>�Y�f��ք	*}�^I.��rmܸQ�Ǐח_~�q{�_�pb6�M>���|�I��\�p�����y<OXXX�ڴj��;5W�M�/��q�p����[��lױtϮN������}�ݧ�Hs����5v�X�8q� H���ƌs����N|��6nܨ��l%%%�O�>�8q�5jT�X�á�.��>�X    IDATL�V�*����H���]0oj߾}M�{%66V�.v��#GԠA�s �7p�@}��7%N�w��}���ڸq���߯��9�N��ƪ~���ҥ����*կ_�Ķ_z�%M�2�ҙƍ�7�xC����q:�Z�x�~��G�_�^G���ӧ�ڵk�s��4h�\��'O�T�޽�y��rs0�p��#�%i˖-��⋕�����ប�T��N�W�p�����J������ݚ�-66Vo���F�aJ{z����SO)33ӣ��U�T���յss]Ԧ�_M��M��Nmݱ_�7�ֆ�{���~�]*��sƌ�!�.�0���O��c�cqK$#�)����X���[����Mioǎ�����7�x�N�f�ԧg;u��4௦z�0��sH��ܪu���hڙ��dM�6M7�t�)����ۧ#Fhݺu�Tu�^{��ϟ_l��ӧu�M7�/�(񜈈�����ƍWl��m�Ծ}{9���{饗t��w�����;�p�	�g	�3gN�}�>���𾨨(m߾]6,�?--M�'Oւ���믿^/��B���]y����+���k���~�z�ө7�|SO>�d��yhԨ�fΜ�k��������Ou�֭����y��.IӦM��?�v���ݱk�.5o޼ؾ5j���ԲeK͛7O�ڵ3��ŋkʔ)����훪w϶j�"Yv{���*��(��[R��ʭھ�G�����C3g��%�\bJ��~�I7�x��=jJ{A`����^5.mU1mڴ�ڵkM)��8qBw�u�.��"���1�"����z��c�����n��|�]*��E�zӕ�ד�5��˔\Ͻۮ8��o�Y�_~�6m��q��jٲe%��Pq6�MӦM+���ri�ȑ�ۥ�Ũo���n3lӦM��*�z���9R�L^��1�< �?~���]�v�G��7o^�FL9�N͝;W]�v�Ν;/x|����Ӯ];���{ۏ=��}�j�ĉ�Sy�޽>|�~��>7k�L3gάp. ��P��ݭ��b���Z�v�)���[�j���߿�����:�ymo=��x�6n�ڴjP���n�[��;��Gn���]U=��[m�^�Z�z��m��f�µ�_~�V�Z�Ν;{��� s�W��_U�V�<n뫯�R���5{�lV~�u��u�u}4��4��^J���"^�,:*B���L���P�N��zc\�l��v�{�G��ٞe����￯_|���v���+�T�6m������hѢr�u�\��{.�~�M7�z��������o�b�M�4Q�>}��[�|y�E: �w��q�04f��
<t萆����\_|���֭[���l6���k���)������ٳ�V�XQ�LR�hؒ��7�tN� �w�yǴ�0�L�2E�}�����<j��phƌ�ҥ�~����h޴��}��������b����4�jV��=5��[t��Ajܰ�w��\.���jժ�^�u�jmҤ��/_�k��ƣv�_���q����o�U�5<j����9r����j�>��j^_w�>TO>2V��vTXk�VF�uu��Azl�h���V�������P/���:v�X�[�K3y�d}����R�a����̨̔��
�^zi��4�ܬ�Un�����b�T���⋋�[�z�Gnݺ��א�����sǎ�^�z��p84l�0�ٳ��LR�b�[�l)��n�����G�𾬬,����׺uk=��c%<�ٳgk��c�>â:�>�����{� UEAl��@l���+&j|�K��QQ�Ƃ-�ް�H�R�}?��7��{��Y`~ו��̹�����ܳa��Ӟ={,Z�H�X,&:�;`łX0+.�V�Au���b�c{[,���������A�(,,DXXz�ꅄ���QUUũS�ʃMI�7?�����+�iؑ��ptt��[c̝>߇%o�2`l���#za��1���N��{bb"���)S�H��=((111��&�B={���sJJ
�>}*��~y���XA�o�����k�0@ꇱcǎ��VTTD#�BQQ�V�4�^�8p��@�����1�-h߰a>|(uLUUUu֍0` ������ �������˗�/X�@�!A�;uuu�={ӦM�j���
̙3nnnx��Xc:��Ū%!�0�/�L�����c0���=u��Kk��~�:\]]�e��V��X,lڴ	����2����M��Fdd$ƌ#�<�<y2N�<)�X+#��s����T1u��R�� O��n�������O����رc�]��Ç������޽���I<A�$^^^pqqA۶mѶm[dgg�=�-�Q-�ؗ$��?���(U�uOOO����j;|��@r�>�����򂷷7���UUU ''ϟ?GLL�>}*��L�h	�M���n�'O����������B����W�|VYY���8{�,���k�M���3:w��Kf�!B�~��7<ݻw���d2�{�nt�Ё�w	�����bbbЮ];��y��%F�%�sK���Za� ��p���3����,D����w�ǖ��aƌ8�<"##ahh(qs�́��%F�%��B~��{����?��R����cܸqHO��f :Zj2�:�K_/�MG[��{���+��o����c߽{�.]�`ٲeX�lX,�V����[�n�O�>Ro�"�� 77W�^������]��QRR"tL]bG�-U����Rj�d���0g�L�:U�.��� �^�IIIX�r%�9B��"A�D��������<yyyAAAUUU�[UUTVV"??���(((:f�ȑmG�EQQ��q�eÆ���;wp��-�|���OD���0i�$<{����_����A�fnn��W�
|/��Ǯ]�0g�|��Y������9Y��(l��0w�������F��|�cϟ?��m�bϞ=����8��� ����������CЇ�Qh����q��i���555X�d	���+V���� �����1$�NC-̘<s�����q��Ո��@߾}%Ze����nܸ!���	����N�P�7n�\~�����V[�=D�R����
�V����ǈ��:����^�%K(��������q��=���J/A��>}B|||�6SSS,]�T�/_���7o�������8H��|||�/\� u�ھ};F��͛7����$�NMH|||��e�͛Wk�;AțV�Z��͛R%������燰�0���:Zj�0�/��J��4pr0ǲ��1z��X����b����={�T� z�����K}0/A�po�TUU��_���W�9���ѿ���Obݬt�h�5���߷$[%MȆ��9�/��A]��H}�ʵk�СCܽ{W�k�֭["k�!9�رC���;v����Y���dֹ
���C�
|��Z~޼y8�����V�w��	<@����� Z�cǎ	��X�۷oo���NNN066�����q�ƍF�>AM����q�֭Zm_J��{�;A�GGGܸqVVV�www���P�f�0����"Gr>}X,&ztu�KG�����|>7n���7233%����'�]�==����!	�&FMM�/_F�޽%������С._�Ly���*�N�ä�����"�	�b������F������������֭[%����6.^�www�� �n���p����k��;w����������V[HH�D�|[N���G����������?<,(((��+ЦM(**BCC***�ի���'� ����Ν��"A4g���;
k�1����Ç8t������C}G��������+���5�5	�h������f���~����"���n�7nܐj��}�ХK$''S������ w��Q���*aܨޘ V�;w�����oߖ��:t�իW���+�D�#	�&DYY���t�"����'�C/�۳-~\W�Z��j`���7�7TT8� �r��>}:BCC�nFSS.\@۶m%O��SVVF�=�m�6���<X}��9ƎKy���L����\�aff&KTT�����occS�ü.���?��#^�~�u{eyy9�]����Pt��?~�5���G�zP,A�T����8qb��9BBBp��1����޽{���@׮]��� ��=, �>}*��	�h^޽{�e˖	�ϝ;���!䆭�-�\���WWW�׮���4F����ü�`V ��(K4.�V&X68|zw �Im��ǏѫW/�<��� &&���iB��k������(���S��|>�V��_C]��1r��8�]�h<���	?,����q��탷���+�tuuq�ʕ:o�	���`�ݻw���Bqq1nܸ�)S�l����/���o�U�e���b�1f��d���R׭['��0d���?p��Ç�ѣrssk����C�+n�h)���OL�8Qh�P��Ν;c�ʕ�s�
q��E,]�ݺu������LLLھ�&���6��͛��HiB^��������Ҩ*--Ő!C�J�Z[bق���l+�C��?��lꊅ���@O�Ҙ��*L�>�gϖ�777���@MMM��D�"	�&��b����0`�D�\.ƍ�����}��b�U�G�MkK��I�GCC3�aD�'�lj[��޽�.]� !!A�k�ҥK����h<A�T���������!���b��_0z�h�=��s琕�U�m�ȑb��vU�۷oq�Ν:�ZYY	杛�����S�I���{L�<Y�}ѢE#&��g߾}�ѣ޼yC����*���իW�������Á���'����n�H9� ���xEiii�v���4EE���^�|Y�홙����¹s�(�g2����fRN�������G������q�F�ux�u����'����JЃ$����@dd$���%_XX<x�R6Ǝ셩��*�)̄|a0�^^�h�0hQ���{t��>��fff�t�R��F��/����Cff&-Z$�*Ԫ�*8p�V���9z��Ai���k�	[������7"''�b�����ƽ{�j������U!����Ѿ}{�7�އb�QWWǘ1cp��9���c�ܹ�o�H I$%%a����s�́��'-����^�*�ݗ�/^��ÃrY5]u,�� ��`�Hj��RRR���ޘ4�������ի���H_����&%7���#�V�\)V��+((����_�N����:��@�έ%�!,���t^0:�kE�NNz��+W�Ht=[[[�;w**�`]���������믿�g�:tw��8�TWW?��n߾-�����H��MTO���T.�+�n�~�j����I1��v��!�&iY5�h)�<d�޽;ڴi���ܻw555��000�����'O��}��"��37AĿmڴ���2��탪�*MQ-����?�6m�H4�����ի���)�w�5Œ����2��z�����K�Äb���G��g��_~�E��D� 	w96r�H�X�B��YYY�ٳ'=zD��֖X�`8�,$;��_JE���G�WJ�z���a���8}��D�sww������V�� **
���4h&M��1cƠ{��044Ě5kʰ���#&&��ꔯ/��uذa"W�r8>�V��ӧ��f�رc��߽{'p*U׮]h��2� ����X�j�v�
}}}a�Νx����[���۷ѷo_���-	��`&����������ؐ�2D�a0عs��ϻ�ܺu�{�yV�?�|�t���C��N>+�C-,����m)����G��ݑ��(���̙���p���d�䔗����+сiii����˗/)��������BJ�4W_>��'�CYY�6���J�ĉ]oذaX�n�Dc	�%�v%�X�lz��-P����k׮�:�����%�\�A�AG��
a�d��Ԡ�U��Փ'OĊ����������Laa!N�8���0888���!!!سg��9�����S�N�ٹ�ڤ�>}h���� �>���X�l�@��Y�ȃv�Q�X��Ǐ�h�k������b�}9�
�2���B8�i�p0y�/��*���Txzz����]oÆ2d�Dc��E�r�������p8b�������{�}�L&B�{����NX8{tuD���r�9r$���$������<�� �n߾��#G
���2e
LMM)�%p# ��̷�dRRR����+����I9ƺ|�:^WWW����Gff&�9�I�&���]�vő#G�,����ݻw��]��UY���2�� �����Ǎ7j�})-S�9!+�F��ʕ+%{����߿Ν^���P���pu���ZD��`���5,�?�"����{�F||���b2�8t�\]]%	�h@$�.g���p��I�U�T������iii"�*q1���&Y�2��21���9�`I�|Puu5BBBp��Y���y�fr�AH)&&�N����f�)�a�)u���Zm~~~��֮����!|||j�EFF����{����TV����~�j� d����޽{		A�6mp��}�>�;w�w�}BB�@������$����xH\Z[[c���4EE4w...صk�D��ܹ��� TVV��kb���￉�C�V�~��A����ݻ7���ž���*���O���I&�@H�]�0DFF�uk�-���C�^�(=��T��9�hӚ�>j�45T1o�P8;Y��[UU���@��Ĉ}�/�Ϙ��H&A��mI �֭�Tsp86�ξ!!!`��5FMM���+t��j�S�	���;A4���8���O�>xm�ȑu�y����.��;�z��N�:���%''c�ҥ�������!"�9���ƩS����"�����(++����fBWGC�0�f���gBOW��@FFz����T��cii��G���bI&� H�]�̟?AAAb�+**B�~�(�|��QǼ�05&��[:Gӿ@�@.���� ܽ{W���ȑ#v�M-��۷�Z�j%�>8ۣ�U�ߖ����Azz����]� ��\hjj������R�Gͅ��BBB0{�l�]������ח�ܟ?�ܹs�=<<�쟕�%��CEE���2���TUUq��M�Ν;X�f����_� �Ʒy��:K��ݻ�<h#d��d����b��gϞ���%%%"�:;Y`��(�_*�h^���pv �<\ZZ|}}���#�uz��U�VI"� H�]N���[�C���x��Ⱦ�Z�?+z�"�-���w�|���Id���R4�޽�:^^^���+I�A ())H6KRz,22��Ϟ����������...���Za����B�6iK�|[���kDK�C�a���X�x1BCCѹsg�����=33�z�_�|Y�-  @f�|ѫW/p8(((�k׮X�d	�;&��Aa�e$�W&���\����{\jj*����\d�-g+L�8�R�n�e��P���C`f*��K\\$�b�%K�`РA��H������8x��[?�|>&O��k׮��kj��9�CCC�-SM��CIiyEiYEQy7���WP]S�ǫ�g3��VW���� PS�c�&���,ˀ�f�(*�uTU9��*�l6�Y�(�d20nd/�YLܼ+|�D~~>|}}q��}�W�nΜ9�~�:Μ9#M��dhii�}��������ڵk���+��b2�PTT��&I}�C�aݺu_�f2�9r$���|�3f̘Zc���(��PPP .�[+Nggg�c�BCCC��EIjDsTׁ��믿dv����Z���V�9r����BBB�|�rTTT�,��'
��>}UUU2�A�JNNƒ%K�iӦZ�ӧO�ɓ'i��h.z��Qg�"Q���1h� dee��۩�=&��&���o����*�\�����˭ί��TU�r|~|����d1k �W���Lm��f1YFL&S_����p��Ԕ�4Ԕ��Lf�ν��+��C��l    IDATq���	_����>���b�
��ߏv��Q:ߑh8$�.v��ccc�ǭZ�
������@s���z�K����s��S�>W�����2�V�P��!�¿[�;�(>�C_���J���Zj��t�5$9\E^1��DUu�=��799����Ůy�{�n�k�?~�&\�h���]���ӧ%�����2Q������<�>}���_��&��@]����SJfq�\<}���*�:��fKT����M�+Iv�Ds���#����@,_�\����LMMk����[o��ݻw�����fll�	&`�֭2��������QQQ2�� ��e�֪����̢E�h��hʴ��$Z�XUU�aÆ�ŋ"�vhתY&��|������SYby7��d�mib|u�������A��xU���3�OeN[]uKM����0U%̞:�l��yB��={,����*�5���p��!x{{���F�p	)��;ͦL�"�v���~�OWGs�i6����������s����>���ל�`k���� �n�d����lk���F=-���g07�7��j<�}/��G�0~�x;vL�S����	???�%B^���|Ȑ!��_Ğ���G���C�سgO�����,,,������}���S*'�ŝ;wj%����ѿ�Vݎ1B���͛b�C�Qll,�����ے��ǏK=����@�]X�B>�����v�վf��9sF��0l۶M ����+\�xQ��	��?<&L��/��������+W��12�)۹s�@)E*����,�����-1i\�f�l���O�y�%��y�hk{�c�W(h�kG� H��?_���^:�2+��heg���f{-M�&��WQ�`������S��^2��~C�V�0m�4�����y�����L4���NЄ999���
��&+,,Ld�RKSs���V�>`&'��ӫ�)G���[�G�獧�7�<����,Z�����vn�z�o��C�3͟�J�OJZNJMMM��$3�L�.�V"�FEEaݺub_���3gΔ :�hZRRR���X��[�nhӦ�X�X,̚5K������u�����~���``�С  ���ƍHH��V{��9��o�LP���/�p///�TB� Z���*>|X�}˖-����z��Q��z]����~��OZZZ�������T�,^�����W��Ǔjn� �SRR.\(�޺uk�!����P�=����޽{E�s�3Ô	��s��<����Czއ��R~��-�Z��A��[�}~�~f�ܹ{4�.̲5GR7�<����OuY�b�rRb���7i�s���>uue̙6z�"�Κ5K�@i*V�^]��D�#	w���l:tH����2d��˅�SRRĬ)���DH-�TV��m�Ʉ�t�e�im�~v�6��Kw\������-��-Z��q���2��WI������? X,&�B}ace$�����q��%���n�:�e�h��|>8 ����?�5�j��}�w�J�����o߾Zm`0�վ{�n��v�bcck����cǎk��[�
$�;F�*�h)~��W��zzz�}�6�v�*�-HJ�<����
3f�Xҹsg���������ǚ5k��ܹC��D3�u�VJ+�	B+++lܸQ�qw�����/�������dH��]���u�y�F?�|���]g�_��H���X�)���;Ό[��^bJF��oS�((*)�;.Ihk�a���P�h���#F���a�l6���eeei�$$D�4�7o:t� ���ѣG�Z�X��)���DW���Crj�����'��,U7m�k��[�cE��/K~:��u�����0�{���6������&U8KA���������#G�DRR�X�+))!22R��y��l߾����	���bٲe��O�0?���@��y�Ƿw��Z�B�u�???XYY}m+,,ĩS�Ğ��m�۶m����ȱ�����J����:nђ}��k׮h766�͛7�s�N�V�w��/^�O?�$�ښ5k���'�s�?;v�h�ڵ+�?���0�����������,�UXX������ �9>��ɓ'�����P�&l���b��������E�c�����0(q�	��UTT��%��z�6��ʵG���<7g��?��K\����ۍ���p�~��oRG%�d��nb5��41m� ((ύdee!00���b������˗K"!�&^uZ�I t!���=bcc�~ʴt��:o���^��+Y@'.������ތ�7���(���3'H���x����d]��SP?7�֭?��R�;*:t耻w���5xx86o�,M�!���°}�v��}��aѢE���nkbb��&Lxm���?~��q]�x�����sZZZ����7o�� ���%a����a��^����c�iӦZ1}1o�<�J�Ds�d2q���:�y �IVݽ{�/_ƫW�������lTWW��� ����ڵ+��틎;�y.����~��Q~ȧ���3g��Szz:>�����ٳg�i����޽;�����:�󕕕����E���j{.�+�� ���'��y�h�&N�(��mݺuX�x��q���PNLL����T�L�6[�l����3g����� ��� ������|7n���NQ������۷o��Q��Y07��O����s3�
��t��GD�!���&j��!V���-v6�>�J�&���I�{��wQd��3f��~WUUwww<�\��u �u� �pod�/_F�޽�w��-J'���Cv�&�FS����%d^�a��m�z>��xCDD� ��
#��:�jM"񞐘��[NCԓ�s犝+))���3>|� M�!��oߎ��0����
\�zϞ=Cii)���ѱcG������+e�]�___p�\�c
Z"�}��)SWW�ݻw�W���9>>044�������L��ٳ�&M�(�h	TUU�>}��|�G����G`��(***8u�T�I�+))AEE455�|���ϟ?#  ��A�y@{�Ν������ �&O	w�����:�$�N�MOOo޼����X�"""�j�*�}�L�'���I�CX�𩸬219{��E��#""�鎧1�[8Y3�,g����0%%�&�x�p�	�<{Od�ӧOcРAb�wwwTW����� 	w�$�	�ɓ'׹�V���"�k�iiiB�9;Y`f��	yRSS��>�o&�7��U3���x�����LMu��v��K�qB�!gϞ�T6��Ο?�HA�=��-[�ԙt��СC��ϟe��AFFtuˏ=z��:u�j~MMM?~�ޛcQx<~��',_��A�f�(**�~�����dʦb���1}�t�K9�X,DDD`ɒ%2���˗œ'O(�!	w���<%܁�p�x��� $�N���ѣ>|�Xc=z�nݺ�,%3t`���Q��EiiEurj�vO��#"�_��E|?R��粽��L((��:Y��;���I�{���������5�����~�M��u4��;��ވ����m+JXX��d���:&��'����9i/�'���z�OKM�@DDD��]��U��_�I>��V�u6�۳-�y8	������w�!/O��i~~~:t�4��ܫ����)S0jԨ:K�����I�&a̘12K���e8t�P���{Xj]>}��`������klll,����l�2�l'
�\.-Z�:�̙3R�6����c�JU7���˗/������%�[���ƒ%K���&V�� ��%%%.�;���ׯ������b�1Bd��]k����d{M�2n~��d��γ�-5� ����~���I��I�Y/��ւ� Ə�#�����*�w�~�fff҄H�A������۶mÔ)S�s���7Nh6����x[�SAQiEꇜi�v��Kw,�h���N�*
�,��鎥>\n5���>dO�2���Xs'%%�u��b BM���2BCC1b�xxx�YB����n�Btt4��݋�������I`�엇gu�Y����&&L� ???xzz�y�Cnn..\��#G��ҥK$�NR055Epp0z��	�ۗ���͛7�r�
�=����7HL���ڷo=��k�fff����8s����$.�u��qI�i�ҥHHHh��	�n�z��w���Ƒ#G��۸qc�U�����	�-�������ĤV{dd$bbb��ӦM022��6~�x�.x ��Fll,����7~�x�߿_h#m,�>JJ�I�CznFQI�����<�;y4c� S#ݽ���t�R���B��5
�¿�lܸ3g�k�C�a̘1҄�Ю���p'	�F�����X��l�c���кuk�u3ǌ��g�>L��C|B�%��z�/�,�;y7�;�e��MV��*Q�EiD9y�����D��K�}o���X�n�4�D����{{{B]]yyy�������,�N7�SSSBUUeeeHOO'g9D��Ѐ����� ��ϟ?#++���(/~8zC022���)444����ϟ?#??999��l�� 	� )���cӦMb��p��Ҩ

,,�>�Ƃ��AyyeMB���n�uv	ݱȻM�ᜤ괣�v&C�,�,���iv�~f���
^�x�V�ZQ����G�"��u���\�ۄ��K�зo_��6'O�����S'�W3����T$&e��>x�ݱ4%�g���׭,�E�n|w�ž#W������۷o��^�Vii)������GiC$� � � Zmmm$$$�yFQ}���жm[$''�7"�z�p�6������[R�s�D�ciJfL���@猞����r`�+��(Nh�^�z�ʕ+b��~��	:u�$U	�t�$�Nj�7��C���l?{���d���*Ǝ�%Mh�}��'�Ն$�.�N}\��q�����cm��Nps~�Q^^,X ּjjjX�f�4�AAA-ԪU��J����lwv�����%۫���/ߤ�Z��qs�l���g�+i��KH�%��,G������>��7<(ּ;vDHH�4�����b�իWptt�<�ӧOhݺ���>�mZ[�"L����῎��˖�g�˶u�:�g�+�V_�sy%~��Q�������K�ЧO���x<������ײ� � � �hlll�c�ݻ��ݻ]髮��G@S�n���3�}bF���O�Ks0m��,{�ߔ��jarJZ���jj�����ś7o```@y޴�4�����9z�AV�T�����l��+W��]�խ��%��J+��L�!�v�ٶ�����r�����t��o*����v-��|L�:U�7p&�����$� � � Z�+V��l��xYVcT���%�?��g�Y�d��l�s~�˷���}����,���Uh���|,^�X�y-,,0q�DiB#D 	��b��t�R�����a�֭B�hi�b���҄&s�
��w�t��X���{�
~���븴3t��o��f�ps�����"������KAAA�B��ى]"cϞ=x���>m��б��r���M\ڃ��5Vv�"�����}�s+L�>��˿��	F��B��۷�=k�e˖AYYY��!H½�����^�s/�Ν���*�}F���2G��d*)%+��)��m��t��\1�o�vf��ɿ
�J�؆�����7興dggS���``ժU҆FAAA� �V��ͦܿ��+V��GII��{J���x|ľJ޷aۙ���Q5t��\��?Q�\:�Z�O�x��X�`�Y�Sh���ٳg�/F1zccc���� B�.,���� �� ---�cbbbD��pw�� 7)�����ү��񔻷�;�O	�x�4ᒙ�^����/�ɤ�EE6�5���y��TVV����<���=.\����Y�IAAA4Cmڴ��͛��������q��%�}Fx���L��d����_&/۶���t��DE���y�6��������x5����
�J���[o�>���	mڴ�<���+�m�&r�o#J��� d��po �G���%��555�7o��>���v�64��{��~K�7�9<Ϲ��y���R�VVr��{���h�`.�Ϯ]�����s2,Y�D��� � � �fl�`2���RRR�q�F�},�����Y��d���/_%/ؾ���cii6l=3���b,oP�u�����>�-�˥<���!&M�$mhDh_!+c'���@ll,\\\(�9t�ƌ#�ϐ���O>V��z�vbӎ3At�ђM�7�}[�c�"���yX��1�x���������pvv�۷oe"!EE6��`h�Cmhi���Q GQJ(+s���QQ����Jp�ը�V����9E��.Dn^1�kȎǖ@YYF�_g��U��Q��;������Tr�Q^^��
.*���/(���Bd�!��X���|��)��@F�0�ׄ�����Q��wF�����TVV�����r.**���[���"d�����rD4,m-�>���`��%%�(s���(*�QYY��?�j|.�Dyy%rr?!;��ϣ��t�k���`@WG������9
PVR���"���By9�ܪ���T������Jvn>���_�h,���02�绮�����e8�XL|�\������
E�e����(;���r�2��155Err�X��N�0{���u�?3�6ƲQ*����g/��v���XZ���pic=Y�M��/p��M�}�n݊�S�R�3%%vvv����6<Y���� dA~]dJ.��������)�������3�����������"��d�������5��8`��~�۷��CQQ����CǮ�������`0���S�Dݾ}�X�t���`g;SX[B[K]h�8*x<�򋑘���w�O�@Aa�l&h�d2`n�;S8ؙ��\�*R�[]S���"�O����t�{����rDLЉ�b����vf��3���TT�?��˭FfV3�������������OE��������01��C=�R�����X���tĽKGRj����NUE	��&p�7���	���fK_5���i鹈O�@|B:R?��̀��*��]���1�4�Z]�¢R�~�A\B�ߥ#3+�<n$?����J����{899	M,v�h�Ic��"<�T�� �Uʜ��6�̘<0���*��8x<~��1d|̯����1�:uĈ8v�,B��u���\�����+Wлwo�����#rGX��\����]���[���/s���~�\۵�"��i���cٚ�(/�?�1x�`DGGS����VVVb�JP�d2��d�vp�7���j�\7'���}��'�HL�HnH�6\]lб�-lMe�0��2>����T������X�EE�wW;�����ƤQ�x<�����T������&!�Zj�����X���,V�W����Fbrb_%�ѓw��^bd���nh���zb�m�TE��3��y"�=O"��kKCx�9���9���%%�KHǣ�	x�&���l ���HKK�ܼѣG����������KB���.�%�����y���b��Qˬ)�N;;Y�;��qiظ��>6l��Y�(����c���K�,\I��%���ڵCll,��\.HII��������z����R���-ʉ�l�?S&�F��خ��w���ǈ>w���>|77ꥑ"""�j�*Y�G����:�;�k'GhhH�*YE�x��n����"Zc!1��6BgwGt�`%%EZ���U�{��p�a��Iyy�d2�`g�.��Ю��R?����x����
Zc!)(���l�.����B&�L%������������{p�r������ۢ��#ZY�z_TUU���q�Q<^�I�ǣ/�N�Zj�Ю�y8��T��X>�W�ū�{��w�B�={6֯_O���7o���!@|�t@�WY�'��/�wn�}.��8As�y�hoF{f�/�3�    IDAT�-ш{�^�놆�HJJ��
����={�ƍ�O�A�r�����ݻ1q�D��8�q��	�3{� �v��64�dd��s�-֯�"��Ԍ���\Z[�3���*,�� JJ��5	ĉ'(ϙ��sssy:5�Ib0 gk��s���!����WoSq��c$&�;���b���|�t���UC������\�������p�խ�y����.��*ܺ���~��Oet��⩫+�o���ٽ-���RZV�+�cq������ơ����}:�s'�Y���K^~1.^}�;ޢ���b��������}[�F�� �y8�1�>O�dޥ�`0����V�ZQ3~�x�߿���9�]1�j��p4�7qiW6l;ӗ� �zED�dW�'Y[��GRJ֭�Wټy3�O�NyΓ'Obذa҆&�� 	w�Dk�]MM���PW������U�x[c,�(��$V���293����g3h�i�̀�v�L���ūOq���z_g2������-�I���8u�,�kq�:[�����t�C�������/^%�J��f����|�a��Iw8"��|�|���1���Cw8-���"zvo�^���Dw8"U������8{��QCu����z�о����J.���W��S1yP��L�t�ۧ#:u��u�U%%�~�%._�EEyP��lm��ۧ#ڶ��}W8��Ÿx�	�<x���CB}����˗)���̄��5����>��c���,XRJV�O���%U����CuM����u�]i������Mj��[[[#!!,�����ann���,Y�(��h&	w�[& �� ��xhh(�'�/]��_~�E��!}���!mh����z��+��cڂ (���vY1?\MM��+���\w�EEe�+��|>�|>���(ϩ��!��Q7{[S��Do�v��l��철���N�aok�����������3���K'G�����灒���wq���6�R��}�!d��d�W��n \���D��'n3S=���**JHL�"+RGQ��<09�����R�]�l����ս�|>�S�Ɋ�F����Qü0z�w��g�G�����	%����̣;��@O���`��.04�j�v PU����5�]퐝[�ܼOt������Opvv���ڵBKe(++b�8_((���&����cA��A�H�D9��y\����5=�P6�E�;���6n�{]��EEEpqqA�֭)��d2�����w�_@�R Կ�	i"I�Ѻ������ر#��>>>�t�R������g���-��"Z� �:ڧC;g�G**��h/��'Nߩ�u���BO�ZME����������J:�<�87������p��KD�{@(k z�9��N��.��Jn.��.=!�5Ks����E��1#̧�2�:s�Ǒ��ĥ�5FzBW���#���[�#'n�M\ݡ4K���AC�C�	�%!1GN� �}76��>������������������Cituu��������2XZZ"?���G�W�Wr���W)=��t�� �}7�w����Z:�E�rwww�Ç)ϗ��;;;:\Y�.�h[����*���o޼��y���#��9I�.��3�o�����ľH�hl����D�]o��&��~�e�+������OOOJ�1����2��y���3&�����
�ɀ��<���S��\�HV�L&�};aҸ~�~���ł��)ڵ�AJZ)!CJE�
�BHpOhk5�3�(q��b;�K�Dyy%�!5Z���n��};A��Mw2���7�k"�}���C=Y15�Ō����l�dv̈����.�P�( !1<y�'+��f�5u�\�̎Q����\n5RҲ�G�M�6M��һv��ɓ'�}��fự���(�"<�<{�����w� !�����nem��@O��z�Z����0���333���ssj!�������HII�Q�bKA3Y�N�2�t�Rt�ԉr�5k�������n�����zж���SYe�Ǌv��ǑZMP실���L��j�q}6����
$��_�+))	���ǭ���q�FY���())"4����H�VȆ����N���Aܻ��rT�hk�!|�@tvwh�qť���nN���!��ʀ��fOg'�f� �[z����	9y��1���p�<G{3̞:��t�"s`f��NnHN�FaQ)�!5y]�1u����.�o1�������ޥ��3y�'��>0~T�f��[l6m�,akm�7qP�%%��{�n��S����]���n�ѩ��,B�HRJV¦�g� !���.�g���s���^�MEѧ����`Ȑ!��d2�����Ex�HA3I�7��l0�L�j�WVV��Gݷg{ڒ�<��>��r�O��	+�*�WP\A��{{�M�%''����<����t�"�КK,�?����A1@/�v�7s(t��NM���l�F�ֆ��q���b"��+�B�7��t��������ݡ4(%%EL���`S<X����db��.�3m04�=C���h�a^�P��n�,B5G��E��>�(ҷ��1X��c����ޖ�P�,MU̝1�]�d6�?:'s,��쿧IJ�z� p��}�x����O�v�M"�J>W��p�m�&����Q�))9t���K���c�PTTDy��C�BYYYڰZ��vGA�
woooL�>�r�cǎ�СC��������}h�"�&������rqBf�<I���4L75�B��ee>f �c��+++Dy���R����"�f����N�Z��@��RC�N�H�����b��i2`��B���͖}*��t��j�7qi(-��d��f�:���uk6[�Ea0 +#�v���W)du�TT8�5e<���!��b2pv������J�ǣ;�&C_W�f��Ό�P��n��PVVě�t�Ӥ�Xa~x L�����SVRD�N�(�\IJ�|#<<=z����ʕx��Y���im�>=��"4�<��h۾�i����/����:h9�q}#Cmܹ��uw���������(���p���c���_�����p'�>|�X�w��%�����%C�>�r���\���=.�K�xJ��=�?9>::999����<���W;��lv��o�����S���ڼW��
��@H�7����՘z�X8{Y-FGQӿ 7Z�hgmi�Es��@_��P�MƯ1v�L���.6�>�Y��h�ƺ�?+F���q���S&�o}6's̞6��-ga�L&#���� ��ݭ>��������"**Jh�]�H���>��9t�� d*�PyXVN!-��X,&�u��c���b�)��Q7�p����СC)�ONN�͛����*<Iِ�%d�ݰ/��^B���_RZ^Mǵ�̄&,�\.������[�n��Ic0��A]1��g�X�4·�U)M���w�|Ѓ��y����쩃��ي�P䚪��Lg'�C�������Y�C.K�z�X0+ f�zt�B+kKC̟ -5�C�k���X0+Z����eI��� |�?��)��dx�9`f�?�8-��S/�v?�O�<sG\������������())��u-MU�8[�"4���sy�>�����D�����&�dM�먱�[�e���s�啾�����]"���wm)y{{�u`������hkcL[���Ԭ��/o���D�9x�RN\B�6:��`���/����Ś��?ie0�>�;��\`0���1�ǝ�P�GQ��"uc�GQ��i���y���T��9���2�;������g%;#�an���s����Iw(r��H�gB_���).�V�5e��[v��G{3|?}9c��z�`��-���(]:9",Է����>�رcB_�ֹ5m2�&�޾/&���f����2��qm]u�v0�G�܋����'τ�Ѳ߱e���_�����E%'Juu�?����D�3��<;+���b�]=�~9�w�RSS)�7hP�>�=xhwtqw�;�3�σ�����DX�/�mM�E��XLL�mZӳ�I^)++bf��-�PeeE�O��y_��-}=M̚2��Q����:fO������&��%eT�aia��S�[Թ*Tx�9��]�uqu�AhH�sNF]�ɽ��������u��n�~�  /����\u-'\qqY �[E�:wQ�2�=*�|�&��$ܥ$����D�v((�С}+Y�%������\�G�ŉ�KJ͞Cǵ5�U�$�I+��ǉ'(�gnn''z���߷���[��!�IM��a0�1ýIR�,SB��������w|SW���f˲-����`c�b��`H#ɤN�)��ٝ��}�i��vfvj6�JzL��C16`����-Y��������K�p�su���|���sb�{t��<E$�xiݔ/22����z�r��  J����zNT���0����\���D���^�D��HN��KϮ�ʅ|Ɍ�Dx��G����ܜ4x��EL�bcc!+���{���s�)Iz�1����ҳs��;#�9�y������]Ǚ�=3+�k&YSS\����U�Vq��C���?III������ۤ���Ԩ�;ø��9�����j�С�F��(gA��̪U�f8�dqa6�_���0���x��O���  [7.���v؂X,�o���"�vD7�σ�Y1e^��F��W��Tʩ-2K�b��W7@d�P�1�a��L��n]�
��� �s�ޘ�������H�%)!^~n�/�⋥�fes�q֬YC��ΗL���1����0✃F�����&�W(���^?CE{���0k���p�f�ڵk)}���^���a��nmC��w�=�Ĉs��u|��&�g&�P8���ʕ+�����VKlZJ4<�u1��`^zn%c+������R���?(R����t����a�L�s�/�Щ��V�?5U1����s�d�$=5�m���� _d�~��ՠVM����`~:,[<uE�R_qH�"���
�P����Q�\�����s�&}���`�Lf*��������jr�b׮�C�M݇���+�q�����Q����p��C@E�����I���B���Hè�aw8<V��Y�9����~����Kگ\&����������g]-^�BBB�Z���q����$��s�@(�z���z-<�w9C���y|��`���X��k�L���X�bj6i^^4�g���fIa6��Kgz���c����l�X8%�V�x<xaǣ��x<��z��J��B�H˖��W��ϼ����5����=4�����L�1#8���e�F<�=cz��̲��:hnn���T�.@����BX�d�ߟ?~�8�ݓ�k�	 ����oh����:�;�`��ޡ�1�w�,�Qǎ�ۖD"��>���'�1�!d;���eC>�� �D,�W������ ̛�
���QB5!��ӏN�ºU�^"#���y��ZS���mE��b����I�E���Z����/?��Ռx��\���8�B.�2%xrssA�V��y_�\�ΥXtt������'��zJI�
>3`�;���O�`G��N�Ȝ9s@��_�%&fg�ol�v{`d��m�9�N�59Q�+}D(�U3;#x<��J�|��g�p8@$��⩰���Y��܀Ju��0<:f7��&��5�r�m �H$��D�R)Ѩ�@)��Ȓ�P��7o�0="<�u1D�L�p8\0<l�������tY��X(�K�"�D�V(5*E��!l߼�[z��{�顠����gWB�"pD���6Y�6���t�;�.�P(���X(������(��*�x<x��G�'����ƙ:2�^�J`eY,V��Ș�awY�.���tY�B�\(J�"�,L"�I%�c$���gW����N��A'B��g���!��=j0�9.��崹�n�H(���B�T,�k�JY��2ц*a��Kᵷ�Da3��ba��yL��x<0j09�c�&��eu:]67x�B�@*
d
�T���z������sa��r���
�@+��'N�����䵗�Q�}ՆП��>q�2l6~��pՓ�钝� �.�N���������/[B�rss�̙3to��	�HAA�ߟu��p��)���� �䯹��c�G�/w��8mm���#B���O�Jq1���9p���***��P�9��#B�������duwt����>7�����Ζ��Z���ի�Tr�p�J)��U�������у�xj[�5v��jgb��L��B�����9�{�GFM�Mf��#c�������y`Æ�H�P�^"�����&"� v<�~����a��A�΀��(F���?j���1�����t�׿Y�>7I!�l�h�u:�����P��J%��M��>c�?I6�͇0-s}1<t���F�ǌ�F�m���������B��m�j�Z}Dh�>2TFb��#.F+�́�'�25b<�})H%���p����5828d�f3�6ٜ��������	��s��r�x[�&dEt�6-,Tɘ?wV
̝��nw�-�H �<��Z� lvtt������wƝGO��4���g���b�J�]�,6Z��R��^��\�z�!��h/7o���,"\�:���颩�g��|"�o]9�~x�A����K���9=�|���?Ӝ9sl6H$�55/,,����*b_UU���O�<&:B5�S4�zG�H�)G@`�8>n��L&&�9��H�Tp 8}��߂{^^�D"p8t/�x�x	��	��������;�V� ����{9v�� �~��_��S�U?��۞��#}�Ҩ�au|��<Y�
��V�K�щ���ھ��?e̼��_Ju
���7��6�.Hф�~��>:JK��RRB$,*Ȃso�vM�J��.`ķ�lu76u_�0����R���]n���lY_0_��ir�~�.LE\���I����@]�W-��$�E���-��9�Z����xߡ�T���CWn�����7���T?���Ǆ8�v�<�\Y�CFҮ�1�4��ˈ�޾kK[�����:Y9yX�}ع� ���7������,��|���-��vM;����� X�<�� �����cp���ؿ=z�R����v 8��P\�%xt��yqZrt��>�O�o��g�Lb6��� ?���f�D�l��'�<��w���~	 ����K!1>�[￼��f����ŋ������Xp��Beѿx���L��5�W��;�>���1�nfg��!�7;3�~6yt��we"r�f͚W�_�X��TȚN6���pAM}�펮��8r�6u�С�A � |c����Iq�MK��%ʹl�(����?+���>ǭ6ϝڎ��}�/�;z�  (˧�?���5�  �6/���d��#�?޼n\��c��,R��d2�ڴ�hv��u�z�ر�ߺRd+ ����H�IO�y�d3��d���?��xO,tx<<��H�	0��:�i��|�ꥯ7J��#˗�c#4�e��n�(���D"!l߲���#�\E*ö����ttZ����s? ��ƒ���7ׯω����ʚ�L!�{��X�j>�9XF�%Q"tjX�HQ�@cswoK[�v({�.�_
�� ��aM��h����sH��IM�����XQC�')��� <���>��g, ��޺]����<�W���Ԯ�����uj��v32&��xW�����A ���%iP�����x���?z����F)=5�a�D�ֶ�Ғ����2�5�h���')!�b!����2QQQ.�~�E,,,:�]"?�6��44tl�{��,���.~ �lۼ�������k���̑?�0�y�܁���S����ڳ���u��>�w� ��'�.�����kC�c
���χw?
�������I'���rAUuKY����//�P��tѫEEEߋ��yk��億�(��͆���pG�EY�A̟�j�\�j�c�w?����©S    IDATS� xb��&���͞��T$"s$���3���*{�lX�j��$���Y����?=�]L?�U���M�$���gg$d���Z^4�.�BO��
'�䉭d39��G��j�������������W`��y�S�����Dc��Ȗp��,)�D�� p���s�|>LK!������w�P�u�ש#�3͇�H%�Q�RAVVTUU=찦�|�m̛G��˅�g��x<HN�?�(3f����S��b��g�i������>7�P]]��s��1��bIa6�SV��s������#����|���[�o�VT�q�%OM����D"�H�f�< %�L�3�o~�^;��-�O�������5���Zn��0��� �5@��k �䒞���S�7׽���BL�}"����]�y�������]�p��U��2Z��P �V�'毹�o���s���bL�}"�NU���egKo,��4��	 ���{H
�ZEɕ�]�^w�ҭXl�}"��������٧?�����1"u^>lX�K�Q��D�_�v{�ꍆ���j°����=VQ��?�9{��/�+�݋2D��&�(99��455AOOϤ��bt ��m�`0Z�V��M�N9��q�N�=��"�[����2p���Ф�.r|'�? 3g����]]]���>���(-���5*����Q�{q8 ���7�MM�ި��M+�w��Dxt)��rwϰ����e�R�"���]��+=_�����ƚt�v���@G�	���D+7�����\��ɞ�&��N��<��������_����w�|>V-�MeZj�F�U�[o_������9z�r�o��/���v�Ӊ���Ka	A��y�Q�G+��n�\�p���D�����������4D^��t��Y86:ff%�;"Ȋes����nwxΕ����vp:պ�tQ���s�ɵ�$�͝��H����Y�(���q��:{��;��}b١C�"N�ᣒ�}~�����"��.�	Rip] S9��:G�0�0����zII	WY`���'�����GI�
;y9��������Ɍ3�֔����l�UW�\��<����Ξ����A	�y�?I�������L$##��ੌU��I$������v]������|��o�U����F/������i�4s�`�#sA�g�����v[uō��Ç+Н���������M���e��tӪ��c�'��reÁ?�~8{��D��;��Zz��{6�]F}t�lb�&���<X��ŋ�邲��_���Ī�`T�8t����[�柿t�M��I���P(��(?ݏ�bs�]�{��O�~ݙ����ݟ�'�]�)�����`u] ��� �@��A����n�'{���3�?|�rե�ؚ��ɣ�hB.�@���Ũh/�J�2���,#�# ��9Nڧ�J�/_��'�S�� *��7oz�I�틁�d�o�N9��?>{d�`&]|��D��Tj*u�$	����0*����|��������`"��p����Mim�l_��RʉWo4����f~Y#; �{��`����CԲ��I$�G@fz����/����NlBuD�O\��;�b���z'I���:5����)�P��>>�}TGy����]���̈��H�w��.��^�a�`v~~�ΪKJ�AuD�;�^Z~�v?vfD޼4Ѕ��ڕ��K*����*�f�=t�ד��xq��mCJ���[ؾ-�$�bZ�����:G�$�������E�)G�b3����O_s�J9�Y�f=�p���N�B)))~����⁁�4����D�r4]=���р\.�5z��p:����������ѴMݽ�-�2KKK�����c�*:o�vd�􍠦�NO����0LDXT��M{�����o�X����{����V��U+�����G��n�=��˵�B���(���˵/�TYlْYAQ�{�8�.8_^��O�]���䣒��_��v�U�3	�B,)�-�d��ܗ��o�w��g�����?�����Ә>�|~PD-kC�0gf2���A��굺yG�^�Gu� ���:âϪ��l���T� wnp$Q=�ݺ5�}�B.m��a�D�������]v�|~ixd�hW����T���p������'�S$33�|��l�&�@�}$٦l݃<����Ќ����=��i�٠���=rVVCb�Z���Ɔ��c����S���K]�n4/���N��9&���?��w�D�]���!�d���+�Ř�B�b!��N�2O�Dsf�(� T�h<��G��Cu�|�����������E�Ԑ�H>s�N��ZH��@��� �U���ӽ���v}t��˯������J��:3�A!���w8�P~���݇.CsBo�{by��ۘ>rsҀ�g��ނy��C��4�Y\�7��:YI4��
;w����cfKk���`��P;�uvv����Vo�O,��M�K�p6�=C�Y.ц�@&�<x�Ju���^H�	�IN��V�l6Ccc�ϣ"C��ߝ�Ȩ	5��}܂���M�M+�w2PQ�� ;#;�lu߮m] 5�}r���7�^�L�ϛ���Ckr�"#�.k��Gm�흹;w~!㇤���}W���c�<vG���NAM-oj��N<���|����*o6�b����f����oV7_}�ӳ�EuBop걚��,�|>��Q����reîO�]x�	M��t�vv�a�ר0=��e�0E`��W�7�k ����C�*-U�m�#�xe=���E"*�|���鋁}��q���8~��?�fw���A����A{!	'�S$11�����׃�=�^�Ct��1n���S��歏?�4�7�����555~�JJJz��0���4p�c��Je���{���vﻰ������Z�Y�<5Q�۝PU��X ��������n���;X��Rc LK6�N0�����QȆ˙�\�\���?�e��T
�S��ǃ<����!SG�4�5X��sqkLBR���k~Y[����G��Es@3�UZn�j_;n��E��8j9)!���h�+o6��d��ߠ9��#G�4_�j�V���E�	ۡ����zOl�!�>j0;��{�5�/2X��w�u�9������I8��"T���f�ϣ��7 ��i������:�`���Z���}��m+��<������=�~�� ��Ngqg��	�>[!|>���+qr���D��2��t��:���;�ǃ�,�Bը���f��͖�>\р� ���JG}]��'�P!��f,a�����n��kھr�P%j���{�|��;�?���*Bb�3'-S�b�z�:W�G�����oT��`ٟ=3���01��}������uh��d���U�i�Vρ�sRP�^ZZ�'$E�^��Gۉ:�`��/k6-���.�O5�$��N*���%����o�#ꐃ5�L�e$��*���|m�&	r���Q1�B.��x�z���6OSg�F�Ȕ��:��t|+�'s:;Ӳ�#�������b���=q��fUZ�,�Η���h�r���?�]�}���>\^Zu���~�t��_L0�y���ʽ�v�9@����~[�Љ&�d�v����Zu���_�Cs�HU��ӝ�Cf��R���'k�{< 5��̶˼�4���3�YP����������x���	4��`4s���e`��Aҟ��OEp�r	��	2���ڼ>'�������X�γ$���BP�L.�Sܩn����h4A��N�g�]Am���?�k�D���V)XU�>/Z�֝��<x��,6�}z���=�("Grb�D�*Ě/@SS��(�	�����ȁ��b��Tj�f�{�;���'Dk��v����t��i)8�4�ۻ�ϣ'@ee������X���SL0�\��=�����(�	p�䕎;�{��cf�aR��A&�DC������q��C�`2Y�Ja����7*��NNp�H\���?�n�H�8�[헉:�`<��Q�H���6�����n��m+!���� x'���4�Z ���&VS_6�bX�e`�h���'H}c��1�DHN�c�FKkh��.9pa�qB�8q{����3���PШ�ѐJĐ�b�Vm{����(�	������.��{i�1�k�r��vmC�;���h�$I������5�r�==�}�;�[��~�f�æ����ⱹg��{��.�{v5
.�a�9X�e�N�̳��O���D����p�;�r9����g�������p�&ꐃ5|�A�qxd�h-�p�z�g.�:;;���ӑo@LX�oM]��G˼�ٰ���eG�{{1l��"�R���>`�� ��]���A���u`[j�N�v���1�Ä�6�`�;Pn�����|>�����C/�n�:;�_Ű+�I .���Y���jl�~�8aZ��_ð�R��4�H󥭣�P����(�	���Ѻ��3��YxAs*绡�!0�&o��+n�Lׇ{.xo��1eq���I����TN�=z�-���AX��l��)@U�����Y�&��-���7�O�N7�0������1���߶غ��e�ML����G1� �݃�0�&��j\��Y���A��f��;����W�a�m�%�rf`�`/���(�	s������Ul���5_ZZ�{�\�l"{�ª͍���k=ln�r�ҥqㄱ�y~j��h/[���Y�q��4_:��X��~��~��ѩՄ�6��uܩh/�t �P��Q�er��c��������hy��e``��-�j/L�	��:����&}��=�p(a��JJJ���cR,�V�MuC�k�M�=2B�r���3l�{�� ���������b�}S�V)@&cO�V��斾�G��d0�Ȁ���V����ok{�� @�"=�#(Q��H�Y4��KO��{(���c�(�ݨn} �0��a()-55�t�\6������C�����nw�ؐ��h7�{^����?�a�M�e"T�w�t �ڋ�l�� �1����3j��d�NF��w�b�����w�l�.@Np� ��e4�֠V��o BƱqNl����� Z~�N��������3t	�0C�xq��c e~F��GÚ/������}/{�U���X趫V)X�Əu�6��0C-=��h�@��Tp�\`���v�b��������|שh�;4dt�=x1h�  �Mc�e��%\���~ɡ���o��=�f����R�l�/�"��:7��^��m��F嘒MI!>ށ�����N:oY}��t3>n'�Bs��݁�V?
��H_��Dغ�G"E@����&��.##��1�b��`2����A&��7�U�&QL�0V��ꞑs)��c�m]�C�s� ��=4|>���P�{��N����e���*ʇ����)U��@@������Lb0��t��c}���qh�T�b�A�cV�� �e\݅jwo��^lv'�sx�j��/vЀ��;0�&�w
�T�F���g�yK���fwp�;�WNW7I�6>T}���TU`��v�ln�;�L�(u��$r`����փǯ��n�aF�,�0첥����ژ�A���޹h�I�4�æ+v�rA�Ӫ@(�_@4T�n4 �����Z� ��4Xb��`>�b�A��>��;b��n$��.X�ell<�K2g�?h2[i��eSp�Dh�^�N�;��/8��ns����i/��	��J�_��f�=�����N��&G��qy�oOM�jg[,�W��H$;F��8�A?t���rL32&>g�;i�J�w�EBç�)��O�b�8Oa�e�|Q)�(���x#�F ˸�î�U��V��L�2n��b�a�L��m�x ��fQ�j�h��JQ3��h�=�5T� F 0�A���q'J?&ٹ���F�/hزw�*�;_�F�gn���p�����"Z�_&��>M�	8��b������ �r����	��q8=Dk��JG��M�ʻH�6�FsP6�)--u���t�eKD!� A��5��DKI��`]r8迠a�|��e���v���]��� �q�-�����jw�\$���TJ�|�x O)� ˸��n�<$b��[
Ƽ5X�'N\
ʳ��4N{{������f�����bs���:�`n��hГ�w��;4�j/L�	�`��t{�.╃^x�%��E�������=h7x&����;��F�X,B�f��A�\ZZ�5������bk ���B1�0�Fq��C{�T��q�������İ˚�� �����`����^�a���ߣ�1��v�¸�N{ [�ʽP9�Z�#x�\9_��<�%1hF�y5�`G�j/L�	��5��ِW��#C9���Et�q�;Jĉ��=5P�;��t�d���$�:�N�{Hb�;iolȖ�q�N�#����R���]q�zo�c�x< �!(kغ��7S9b�fCHI
\n� �]�D-c�����Z��E{ �)hz�����- z��`n���:�;2'�S��[V�z�����>�.�Iܢ �i��tz�Vpw:�b���s�v�=A�� �t8�_D��-��"���G���栽Q[�
q1��ܦ=�$p](	e�0��ݴ;�A+��]H�;[����p8��\���i��dS	��P9�\u���.����M{ �78��Mp���4*7�>S�	�2�G�4GP�ӹ�v|�On���3�Ͼ������1n��h@�� ��ol�;|>�o xE�{����������@��vӾO�d}A�|Ĩ� �\��>[��y�v�|�xp�M��_0����`��q�����E�ө���w]�����Ȟ�|�%L{	�������IC���H����$�O�w�����$�����3�!�x<`w��~�$
�
�mZm����ptN>��b8 �����Y�,�/v��"��P ����7+�{K7�X,���t�  
�Qvٲ�`�k�XD�_���1�e����kJ"�@F�� �/�ٗY���=���W����~'≂v�r��'��\�����;�la�/��FN���Gp�vQ���bբ��a�+�U�D"!�W�bX_�b8 �}�|? ��/HB(� �XL{�[1������Ͳ�����z�l�/6��"�Vp�avY�{�0_DB��v��H P�m��pR�^h�}�;�F��ȉ:�`B��˂ٱ!�`�&���-+�E�/ �Bs���GTp���`�>
��DI�� A.��~a���s���	(� e�t�F�#��X��b�a6n���(�Ak���7�0��E�,�l�/�T(������QE"A
�]�d�aDV+�R���$�E�t�dct; �5��k/BA�fs��OV�s���Ҥ��p�Np� ��p��BAЖ���Kҟ������C�J�Z�]�Q��mMh����i�r�4�v���2�2)��,�/X�IEsP3�T(^�a�-4h�E,\�b�a�q.�]���E(@�º�v�@�L2�.[�/�ՆH���F����m�-k˽���"\]����c��@�G)76t��!��p�{����P�e2�Vv�>ub�0h�p�_(�}��_6���}4[#܍F�؇iC� ���H>ؼvA�\N��j��;�0_T!��<���G0쎱d����QzV*�i� �bq��1�8�Y��Z
�\��PH30쎍�d��(v%
������m�l����E(@���z��� 96�u'B�|���H:`B(=Ws��P�Rnl2|]~����[��l�;�c6��a��[i2��T�EBQ��C���~ ���l��\�����d2=�p�o`�v�r���غ�մf�B����~��,0�KT�V�re~�]ȪBd�1�e�8N�]שi7 �jB�1����`�����Q��P�"(w]����e˸�5�X�:�Vʖ�f���M�-    IDAT,q�>��^X�XcU*$�P3Ȧ5���J���e�r/T�w�΍f�N�
�A��Ab1Y�ݗ��K��_���/,"�&���؃��~V���%6ҍT*���1Gp!�������M�ʻH���1J����Q+Wa��c� �3V�H j��+�f]�z�]�w�>������Mk�rh7�0Q��D�m���Y#�:N����/.��>X�,?&ZJ{�hV	�84�:�ڍ2�+t�L&�=;�-�y xs[�Q.E1� j������ٰ0��%�`G�0��C�!���Ě-ޣ�����pC@{�� ��U�A�SX�5�I��ܕJ9׸��+2�(��?__���Up�:�D�4���͋�Ң��cD�cуt`
	�(�5k��c��h�ڷZ�(e���d�*�7P3�c��7�jB&߰= l����/2���sj���0��u�W�|��Ol�/v;�M�>T�y���z��((lڻ|�AC��ؘ��`��ӆ)Wb�eӅ�D��I;���2^Q�Ȉ�X�U搊�B��|@����)@E����^S�H�5�Urqqq1�J��A&�D���k�C%���� ���߰j^:�qغ����0��n�V�H�h1�:0�$�s����
��HD{F6�R����h�&�����]�	X�%2BT4Qz�v��X6_�7���V�s�3HB\J�q6E���5�A�R��B��i7��WD�$�1l�i�L������\A�!�P�dr����b��J��s	;�3��>�����P����Ȋ<B� �9D�r����:ξ@R�e~��0¨���|�C�>R�m�m��(QWX�w��M��UJ�@�	{�v��ۂa����,�H�M�ݼ� ��9irrrD�I��1l�v�l���7%I��zu�
�8a֬�MKN�D��˶���އb7!6�|o*x."\-��Ͷߣ�6����м�b�B�����"��Y�v�0�m�T�_�;i�E�������1r�����ނ�����8�vFSއ`�Q������cc'/�m�Xa|�l�]���(Q��a��"�N����98�}������F� �5t��M��q��T��I6�.HI���a����,�:�Pl'Ć�0a6�]�%1>%E��]Ţ��,���5><���?�n�2R��Ѩ�/' PWϮ���[$�Iyᡊ?�'Lld�kB!����rASs�v1�G����k��[�(�	��n��(#�����g����$nY_� �8aR��°[��n��4:T�w M�;4<Fǐ�&T"~�x%�`6� �א��v�axd��*� 텋pPP���==�o��>!���e��9XC�M�R�HH��u���'<<BBB�����.�t"uH�Vm�R�S���8A"#�oI�b��Y�2A o��$EEoZ��8A����@%B�_<<A���H"^Fz\�c��'�Ν����966ݽ�5A����%3=��")�qBl^Q�������lv�z�Ɩp:](����?F1L�-
���F'`�f��k����E1N�'�팊��ތ o�H���n�?+ .n���F:��7<�04;�"���[1y�xKJ򿕟�h�	�җ���Mkk�ߟ�)�^��JYP5"��TH4���v{m���ݹ�����s`Fͦ�Ǿ�b�L�<	֯�����R��fs@+RJ<&��%9!�?ь`놂��R�Q�Tuuo�EX"�D,�����Q�����wQz-JfWmc'��U�k�h5!��h��(�	��X!�����(���N�2!ɉ��m����b|�;�u��Xf=}�`�i:��;��eΊ���i)��ò϶`�����S���v~4��`���. �H�u��BBd3H��;R�^�.�|�Mp� j�8����Y�]���+�1eP*$D��e502��f@ _�HkA�N-����F1N����2�%����\.���64u�ӅU���Զ%��b���"afF����  5,�( ���@�=#31�x���hY�f�~VvZي�:n��˜�O�Y���� ������JBNj��`�{Ff�o���:��'�.����b�1l{<V^�x<xzb�R��{P� 1V�^�^��<q�4���ʶ���n�����88D���*D�K�!k�j���4୲  5텀����{@ӆi���%�����<�}Y
Q�� L�F��==>�~�-��T^o@�=+;iU��|�ikt���E�f�ǡ�WW����1��p����̬��[��� ��ự�aJ,�W�QL:��|���@���i��g�Q �yT�R��nw�\p��	�4:շ��f�)m��Ky��Q�#�s'��SbJD"!���QZ�'l�^kD���fNS�ND]�2_����vq]�Ѕ)���hZJt�S�E?Gs��c����Nގe��F#xؘn5*缄�U�z����t�T�9X��O.��P��Y�GO���`�� ��:{^F���8����t��I�8�x <M�)G��c�
Ed�FC�gW���\ӦM���w2P�t�ͶD,�쬤#
���?��ϟ>/g�o����fw�5�
b  �W��l�j��I�r4<�>Ӽ٩Ob��E+�@�
���S��ĝDs���K�Ϭ��9X�o�ige�! ��1kz��g_�74t4=�?9I�e��j=k���Եq����ś��Y�bzRxY�N�v	y�
�~��;m�kcnδlݘϚ~eEEE����N�d8�� ��RЩ�t�^"t*��O��"�#��E;����I�5����O@$���?�r�(��~ATntt:DGGO���{�x�O�J���G����xJ$"���x�e�1���f����7m��h������L�y44�zu�dZj��R�6)�W5�Eq���V+�-x�ִԘ�g�Z�	���ha��Y���8ѧ  e,?��_�C���LY�������F�lXP�7w�N��< �rb �z  �rR_yl]�T'4�uc�+9sR�c�����|ș����"z��e�ʈ���=6���l�2����+�����d^FZ�1��LO��&�Gh�����;X�.T�y3g����|�#�n�W�:�xB�2�}����|�Zu�Vl$	F�����;w(}ޛph�ىw�և�z�%�r(CdO����5y�;�χ�,�+�P}'��"���Y��Xq��C�s'��2o&'��0���\@u�\���  ��2�=�}�Q�<$�EE!Y�QU��j	���r%�@@��1�Gl����0w�o\��e@k��͝5�\.E��-T�n�2O���N����a��ż����[V�-@sB��]�� 7㯘Qhm���#�;й|��� �6T)�7#�چy�hNh��͋^͛��UL׫��7}����X�*-'�.�K�=�mɛsf�b��>W�������N�6d��[?�ʰ�@��m!�#���P�'��d�¨�<��3f �X���,߇`�Q�\��������i�"<b��=Y\4��S��F�Cҟ�邾��I�����B���^UU�b��u�Q�y9i�}�7P�<}�/bF� �����'r��j��σ����{|�W�<8����f��$!_�ܮi#���so�ڗHļ���+ްp��d���q�g�TF �z  (�\N'��H��/��4*�`��ig7�����?([7���f	����Ηᾗ$0���Qױ�a�̔�[�6�&Z��_�7<W���B!n�h0̗��>h�@�����&U���:�Sۊ~�(?�y�L+��e�Ձ�s�@ ����I�����b�cX~�M�!G@�L��x}�VMҧ/�ї^9��L"��''i��!i�v@e��U����.�ѷ�;�Hvl_�꿺M�^�����q��A�n6[�\�-T<@An�/=�2�"݋����|y��93S�#�V	n7;��N��kn�iE�!	a����=��#�z������ִԘXl_G?����7���Q�R)�L?����/�:�Ⱥu���fN���
���t����.�q�\z$md�FZ� ��x�j�i}���y�υjxu� �`4���D����^�>91R���ֺ~}N<�#�l۲�d�%���S���hh��tA�c�U������m�ظ~}���޾��E�����N(����L%��������ߟ�&z<@�̎6T)yz�ED�r,��[����4���h/����v�vH�`��	�����@Ep�;w����=;��#4�;�H�R�1#,Ü9���knn�)86�  '�� �7:���?wں����z D6n����6#+��:B���z:3I�����B�N���O/��b[V�-�?szKJrZû�5v1����������ˤ���rk�/ѝ�������˸��N�cN+j���	��
��q/� ��JQ^δ�[7����߲�GK��jT
��6�O]C��'Ew�0ܼՊ�'!.B=fF����Н��3O.�U�0�W�b; ���W�]���&��ý  �H�K�JMj� ��Y�W�[uaQ~�W�|ܭ������I�r�(��񩽴���)��&�# 	�i�I��u����TWW?�p��+)� �������	Z���PZ�����ǅ�?�tQ*Q��>RC�qY������,�d�b0��b����3�f��J�|c!cQ�m(xz��̦i)�z�N���Zk�4ͭ�P[�_�������7YF�\�>���:4�u��.̾F$+�(���_��!}c�b�hQ��|�k��l^��֢w�-��6T���E3�`8  N�� �݉�G�������_\s����l�/Y�:U�ҳ+�/]<�g2�]<5��p�<8���r�P6�>B#]�8��3O,���a͚���|}c�¼��5����9 w�P��D�x<p�@�; @r�>li~֝�[~�����j�ܙ)��9sRI9]�l��A�#�P9�x}���AL�v)q��O��fiy< -��guH$���0��  �NH��;  �L�q�ߟ��x�`��U�Nz-�{��� �~@�)G��T����a�$}z< M���5�D"�?��>"�&�܍z�9  �����¬�_ر|_QQ���S ذ!/�kϯ���h�{a�J	�#���8  �L�WjrTԒ��ۗ���S ظ&ƫ_���h��)CdD�-��=PST�=p��p�$�  kz\v����} ۘ��_�[<�dQ��b1��  ���E����,��E�(w�/���g$?���*޸p3�_R�i���s�F�ϝ��JӰ����J��-�ii��;dʮJ�b������on�ذ&w�_��֢_.����L�K$����
Ԟ-LPQYﵟ��U
��E�����$Y����H������(�Fr���y��rM)��ܼy���Μ9BB&� ���G�$��B����Ҁ*��A	_�C��̾�.ݽC`�X'}>o�<�H$~ۣ�.> � T�xd�qrT�Z,�n��� j��


��ѣ�>�o��D"��CL��1 x��S��"$D�R�˻�������u��̙r��UN.^�Hǰ��18v�6��#�O"���Mߔ?:��v8���@	/.*
�G������@��D>�w��EI���re=��ɘV)�EYߌ������>�w�/X�6<Z%kFV�
�?��.n�>��9)wD�P~dAB|��j��%�~�j[[߷����׺u�����7�3r��N�b���×��#���!7g�UdZ��ǆ�c���FDh��z�^��ڍ����&Ć����Lr+��7g>�` �O�����X ������&�G\�G��v��x���4��~%)1��ɉ�:,���v+T�n%�n�>�s��D���<���839!�E�
��?���#G�����(^�o�)���%Z����7��@�Ҕ����Y�Pyyyp����>����1 I	�t�/�!�� @Q�E�>�I�>}��RY��p�ի�zA�A
V�5���vCEE�X�¯�z}~��V-�^o�nb��T�<�Ⱥ]�>L�1G@�� �?�XI��-�OT}��;�����k�`^:D�k���Gh�������#{�瓁Qӏ����^��5�3ta!�HO�]C�6�ܮm������d�E���R�����������?�������ᱟ�:UIK�yK�#B��[(�I	w� 8{�:�I�%���JJ�_�[�.\y<���b��Sc�%%E�tv�WC��w������>�>�����d��f�� �w��׋d63>n�����g���ҁ@��Yى3�2�*�c��{����o�a��<��o�D��czjl<��e��%�Ui������`�J�3�Xě7{��6{c�>�J��'{_�<ʉ+V�T�������jR�>��Tp8���s���Η{���䪜*�2~~��mƱ�����S��#?:t�
-�7�(�P�J~���#ZOVh�"��d�#I�_������Iw ��5�����ȅ���jɟ�t�F�1G@�d����2�.�U��/�r"׮]���C��"�$	V��f��ŋ~� �J�j�:Gcs7Xmv�Jȉ%  �!� '�OA�}j�7�)�N8�B��ƢE����������R@�t�����ۄ"&��FFh�u8��NOַ��4�Y�8p���������CT�g#�C�%%D�c7�����`�`4Á��}�r��������}7#%�nd�t�h��ǯ�ݝ���H�vnS��O�赋cct*�͜�r�o̴��ù�۰�0��_�i)�Qi)ѿ̙e�E����ѱ�����>z�����aŊ�
�B��Z��� 2BC�ֽ��[3W��â�LH�KԯP ��������7ge'���c�b�h�;d��M�ro��9�j��P�bcb|��P~M�ɸr����n0���*!w^:������Hļ93�s�HVV���{��h��'6|PRr��k�'�e���ڐuɉ������G?��RU�����O��R��y9i+�nϊ����޾�3F��=�. 
�6�)��RI_�*W�$��bC��/���V��.��\�K��W�eɒ%��l��j�`�*r�  !!2�ؐ�� ���9�P��?HWp:]^�����N�� '���z ����(Be���rX�x1�<y��].7��w���t�/RS�r^|��7�8=y'��$:2�x�t��	M]�>�D�t��=e.\�@ǰ�۵�DK�܋H$����xH��ł���4:6f�۝]N�s��t��x<!_�W���T"�S�Ȣ´J5�Z۾8r�*����$g�WÂy��J�܋L&���L� �=xuAn�}�`3�����>��ep��<���Z$�drI�:D���J�%c����`���Ͱ�}�/���$Шɔ
��J!�=#i. �u��;��[F��bms:���{��t	�|���W	E|�B.MT+aaJ�DL���W\.7|�i)x����=x< �|�����D @�N-ש�"�������-F�e�l��8\�!��ep��������b�@�P��*�N�S�H4���l����W�^'|XR
�ze0uq���[ �l6���3���g|���t:��.����B�N ��bad�B�Q+t�0���(r?zz�����5��#� |Qj&)!R��� �.,�v�c��븣��t�]n��6��&4b�(J"�ׄ�h���� ��vkPgr|���+�/Z�BBB�d2��yk{��VP(����F��p���cǎ���(�5����^����V����� d�$Xw|�e��r�"����t:A(��O�jժIw�/Jm��%1��� �u��(;�X�$)AG�o]C'8��Q/\��� �Y��^����" 2�\i���(��� t 0����C}c��Q���v����v�Ɉ'��/x< ]�J�S��l�������A`���b�7v���~c�.�q/|>�n�3;�    IDATfM, ��~�*���~��A�޾�x�y�����X�DB��k��zm $0=�x ���4�f��B��5�p��:<�t�C�D̋�օ�F�4 ���x���p��w��38K�˙s7!}Z,̞���P@!��� h  ������h�w?>��0СR�],CQQ>|�D~��w�:`�\�KB|\��Ǘm���}Ds0���	����UNf��Ք�]��ޯ� h)OHD"�����l��4�ׄ�y��n�QR�������j�L ��C�Q�������{Y�Z��o[�>�<8�N�j��S��E'cc��Ʈ����L10h�]S�ЅAW�|��<�� J}cW��{Ŧ�v+�*���0�r��m(��w�(�	�<snT�0=��9x	�Zz�+�p����}D���·�`h8���`�v{���N�ш^W�q.\� ��%s|i/7��z,{%"\�kFs0����D�&|ߠQ{�����^��?>(AM̂;�v��	�?;}�tHN�<��`4CC��.�h�
���{�9a���촔虤��\n��ccC��ƍ$�����vD�?:<���g0j�ф����_�l<Tlv���q�۝L�8GO^�;uL�U���NA�W��/��Bo���`-m}p�Hp���n����	0��߿���\�� ��0=�X,6x���r��
�8x�j냻/�]�[����[�f'_�>59*��'W,&^����ua*⽆���a`p�`q�N99�9v���EP
�,���:�֮]�����3�&-%�ŝ�=�X�1r����c�띺�����D����������k8{�&YH��G�ᎏ��̧��Cc3Y���~��LQ��������)���lx�ͣSVD����[��2ncz(�`d����1p��f���	�x�$'��I[G���Rki�O�M�L���zU3;U��0�BE{IJJ�z��۝P}���aQ���Ah����sg�Ν��D�w��}�G��u����LH{	��`ܻ  Uq�r�
���_�s۶m^�_���H��Z!������c�<����i�ь���Uy��eﾣ�>�>�g:�tP@Q�`��hT4�Į�i�h�n�l�1����+��X D:ґ��H���a�����9{�0���0�<����!K�5�j��_������	����7������{�y��J���^����L��`�ۀ]�/��+�
E8��������9�ŕ��?#'[���
@e����I)���#��VTYy��X�=����AQL����3q���v�{%뢟�����:��ܭs��'L`dr�6yY�?[Y��{^��~,y�e��R�WWW���PE�jI�'���	my�PqZ�H���`��>]�ti�y.�OҘ�����n��gZ029Q���&p��^�|���<y-mF�Smm-"""��
E���:�\� �q:N���s�K������)'��Q��t���;\������g�Ц�_�r�q���Dtr�u�|�hWy�%y�(�ϷɃkJ�}րݿ���K�� p�Z$��3��*(���G���o7g���PX(}
ޖ������hX2c�X��d�����|����:}����O�%~�355Ÿq��Ν;hjR��� ��JZpWеkפn�b�0g��m�1����H_K�X|��ɉ�-]4aaw���-���Gqq�u�&S��� ���%<� ��\EQq%ӡh���<���St�T]S�����60��	���+��_^eI

+�۱���K|K�]���)L��Q���w�n��e/�P(�!� �g��.�&���[1L��q�������U3�F9s!���O�QyE-v������9.�e:�޳gO���7�<�/��Gi�Mf�]�햾3�3F&'*'��2�h����a���̙�CSSf��gJ[_p���	�\���F�sy�������k�1��;��ɉ�x{{��X�!c�R�k�M_�+M p�\��zV׈m�/ 3�N�����__m�yr%).��֝�PJ9��v;$�����$-��]l�9��M$㏳w|7��P4ҽ�d��k����U�%f3�F:�.��ɚhr��������_�t(G$����C�'Eŕ�y�T��1
����O�ڷt�:,<I�p�ñ��V�^��X D%�-�˭����*���k1U�,k/"��.]R4,i��/fm}�=	*����r$u��C��ٹ�����Q̤/�p�`����X��f�*�F�lcf���%��H�,��f�R�WWW'ӭ�������_�� �G��u*W�t(����v�o�9��b�?�!N_��d���=P��sOB�=!��E�=|��ݿ]Ac����k����D��1�=y�ݧ#���-��8q�6�2
�r����. ���QQQ!u��J,��_��y��f��0��
�029QK��::ڌ��=�N�X�s��;v��ㅄ�Ȕ�IN ��}[_p �W��t���,+V���&,<��+���֫�N����Dٖ.���ͥ����,�<l�0���I=���?����Ɏ�x|�z�*"�S��1��q���K��I����@(�珛��f?�)Uaq%������校�����Xt�<�$-;��g��fDE%?�:O7Ϥ� 2�|��m����Rl�A7Ϥ!���ܥ��6}UlB��D7�����q��E��;88`B�I�0wʽ�����oO�X D�V.����N���?����˖-�Ñz<Y�9p@��@��
��� [�
eggc�ڵR�Brvv��ݻ�]$��k�SWkXYvTf�R�hb4Į�����(���2a�#K&�n��q�D�ēǛ7oF�~����Ó'm���\�b1b����C��Op�%�M8z�&B���SY�B<�N����ڀ�4S�VY��ރt�TFM��~kˎ�dc�t8j��_�]�/S�U��!*&N60�h�t8j���{~���*:y*���*$&?�K;�1�ڄ>H�!� 44��!���)FNn	�\�BGG�Ţ�L$��H��3��v�KCC/^,u{}}}�)I�J�0zxoF^[l6��f፱�m�{�n;�Vj>X:�����6#_�3��p�Ft�ϳX,;vff�}�X�j�:;� NՓ0�=��Pi�ź�:��	X[[�7ސ��ƝǊ�%7C]v�NC(�L�f�N6vL�?<u�͟�066������q�\�
�b1|7?�:����+��O�J��/g��t(��@(�ًa����϶".1�o;���b�Ci�x���u��I�<m+"�R�Ӯ�t�TN�U\l�}���|�&�H����{(�ݞ�WTn~���YƊ�ScG~��3w��{�*$&?��N���z\n��v�nD���Ryܽ{��ҧ��5k����}����e�&;[����S�@���X/Ը�>c;�7nK^??~<�u�&�xw�ܑ��LNb 7T=	���	w�� T9Icc#�~�m�ۛ����ϯ���+j���&Ɔ�Of&Ɔ�2��8�2#�,�?vx��N�jii1�i"�q��&�뛚m�l�2���R����.(#�6���QO`�FO���b�
�Ǒ�7𬎙��mIIi5�g����L;0����B\��3�������#)%=��¨�F��o��_0�݈�U
��H�(�Ӽ2��a]ݶW�����������MYB!b�2Q˭GOg[p���W���2�:pi�k��56��
��m�j�W���bׁ�((�>Oy{#�йsgxzzJ�^KKeee��~�m
�+1n�;���9�jin�fmi��8>+�� �B�[>e{o׮3������χHL��e��R�nܸ		*߈z`��'aR��+�z_ �I�hii!;;���R����ݻ7���ϳ4tPO�xw��B��@ G>Θy�/�*cA�-_�F��ƅ֖���~���>͟Fg�XHLLD�^�������������怷掂�9#�r�.7�'υ�)e`� �A.�7{8:�3�R<I���?CP\R�t(m��cF�����i��b1��s��˥�<e3���S�`�Ⱦ`�[�W�P��{	�x5BbQ2"��&��3s<�d:�hh����H�	K��<��l��^c�ݩӡ(EMm.\	Gx�Δ��������t��χ�����߻�=#<��n�l���9�U��N�S5�Vd�;�G��w���a���s!oi���!++���}v������-���bs~ ���'aR�;F�zE ֪r�X333�5J��,:::���o�MqI��	C]e�)6��22ԛ�������Y\F� 2�0�-���%c�d�b���M��6�=c��]+��dBB���M�+UIY5B$A$���c�5U�Є��8q�6��U���r܋H��6]�[퉱�:��3�.ݣ*"�����1鰲0��3�f�!��}��VHx<��
|��)��Oʁ��E��힖Q�__ExT*�SV��&>�g!=��]�aԊ7��r���?�S�(%���r��a
��k�ݱS��M#�p'4�]GNn	�����4i�ԇ�����������?�Vä>�}60��4��'�ٴ����֬�n�`gc��@�b�*PS[ߓ�$n�nܸ#FH_��СC�)��S m�D]��V-�G �r�.]� ++ZR^�ljj�������yq��E�+k��������x{{�7��������b�2��1�5�޽�ѣGK=�ڵk�g�ECk�,-L0m�@ܳ�\�nl��nX"n�y�3:u�N]�Xa���p���j���r�q�N,�%��G�N��ͥ�OܪN��U�zp�>�S�j�b�0d`L�8�U�=��-�ՠ(�%f3J�����Q�zcҸ��j�&1�)�ވFfvӡ�+�z�0�cG���>3�d%��0&�nDӍ<9-]�>>>R���$�ͲE�9�E����}nߡ����H,����99�tg2���Cq;4��獍�������ׯ��T^�4@UO´V�uZ)T�V 1y�d��o޼7nl�y6�����T��-95/t���ү��[�hªA�1��*����g�_��M�A�!**J�1akk���Je��n��v����0��::��s�������t+�]��d���1y� �6[3oH���#8$�C��2ú;u	ѧ���n�W"(8���h��A,����'�c���1-#���b���-1'*Q-��pƴI�4�F�X$$��jP���	e&��jc�G/L�0��:h-
E��I��Q()�f:�VM__05�~�d�ر�{�n�ϛ���o1zHI,#&.�?}�0i�'kf^���u&�1TV?�7ߟ�@ l��_|��~�~422��%m>�оܻ ȁ���o��._���hyy9��Y���쁕�')#<�<��<~����L�A^�|���n]���t]��I���Aۜ9s��K�i���e˖)�����q����s�0+��QO���&������C]1tpO�i�)C�H���<�G=ALl&��?`��jo���<���W��K�F��$�<��S����C\0�o7���ohBLl&�G��	e�f�ѿ�<�Do׮�*�����^D
���P�&���`Ȁ���N�5b#���ѩ����jJ��,�v�)M�k�0}�t�m�}k,FzJ_\R��q|�[���e4�Z+O�2x@���~o�;s���}^WW���>��%K���+#�����LӀ??j	`�*'`�XHJJ�����}���`˖�70Y,��|�m-���D"1b�2�>����@�K�[6�Ww'�XcCF�
�"xo=)�F�޽'ӉY5]ij��v��砞4���:wYy"�����2:��X,z:��s���q���zS��#"�	>JGMm�Z�&��hi�w����ޮ]�����b"���E�z�G�hh�M<M������N���;��V�@(D�<DD=A\b6�|���t��1x`xꉮ�Vj]Lmj�#6!ѩHI̓HD�x�����{b��j�1���я�����6���1HOO�#�����'"""�}ެ�6���7��=k<y�;�Љ��B^�zɤ5�ܻ�g:UkiY56n9)����,SZނ�899��S�g� �U(V�����������ǁ�n_]]GGGTW7���ݩ>�d.�;���	�k�RBm�v��.֝�R,�ԼZ�7���ܥ{�\�x�gϖz��ׯcڴi��F�`inמ�p�i�vJ?���6 -� )�y��*B!�k��l�m-���ݝ:�G����S�|Mm2�������䧨��`��͆��\{����=��u���/)e�HI�CJj���SJ�VLWGN�6p�aמv�bg��v"�ye��*BzV��䢱�6eZ�F�pt�Aw�N�^�� /��WP���|���!=�P��}��L��ݩ\{��ͥ��:(u�&Y��HI�CJj>r�˨h��z{��͛�4Ir���S�`���ӔJ����Q<��X�c!��%���v8�����:�C�O�i�y===ddd���V�1���Kl۶M	ѵ�@�(��E�l<���(===�����Z�ܔ�����B9���M��~��d  �����G���	y�����٦�q��%�y������P���l� ::Z�/�&L��[��"��͂�eG�X��ڪ#�-;���&&���Ӂ���+'V�x|45����GU%��(.�FqiJJ�QV^�п�����N/^+V�����`��]]�W��76�����5S^Y���*�V���Eŕ���S�m���6:Y�����k���֖���}=]����~��D}C�߯�Ҳj��V��S���J���{[e`���6f�^^�M��Ӂ��6^.�(����CC#��<����ߡ�*�T�{fll��6f}n�+SXXCOWz�گl�"45�Q�Є��Ɨ�[JJ�QTR>�j��U�f��?�X?��bce
3���ц������@ Dc�<p��(.�B�?�&�TQ��Z ƌ����f����`��шt���ƌ��>G�e0K{�r��Y}�.��i3��,�I.v�"�������/�H=&��E�.]$V1  i��H��w �0CՓlڴ	�}����kjj���$�0��\o�/��'fp�7�7�ci������e����r�fȩ��a �bμ���E������͆���/"M��H��h=��%�č9B @[�mm-��b��@Z�bSO Re�"}}�X,��J!DZ�bS���/1uaVhh(F�)S�ѣGKl�)u���i�C����t,�ѲE���v:c`���b�H$���Π����6FFF��̄������ܹ�}��2BlI�1�H0�x�u �V�$IIIX�ftt��f���]]]5_p���G=�K-DU���,+ˎ�;w2����|�t<��{˦�r����071d: ��/���J\p;v,~����]�n����X,�/�/�D*"�_���O� ����(.��P���B�aD���.��H��g]J��JKK�p�B��w��111HKk��maq\�픞zH����+����f2O{�f�e����t_l�[!�z"����_���655aѢE��Qˍ�o���#�xѨ�5 �������퓩�G}77���݌FqI�"�)�������5+��</>y��eS�uw�ylnj��t,��E��Oݖ��EKK;w�iܤ�$�=KE�	!�B!�4��ի���Ν;������b1p���9\���H�����{K��d:�����S6�q�zTr�@E%��I~����cÆ2�{�����*��� �W�D��=�p00J�=z���>���+>�f������'O6�F$�i^�{�*�����l:Y�z�8ێ�4�w�ޥ�Y�l��^.]��3�S�/7n?FDT��6��V�X!Ӹk֬Arr�"�B!�Bi������J�������o�ͳ�٬�    IDAT�F�X,�8�)#D���h�-,:�ekc��y��xڲWM�����S--6�n9��B	�d �����ׯ��c666b�����U4<i����F{<� G�|�]�����g���L�6S�N��&+���%��V7��cj��\�e�t,mч���ֿO���r�	 ��k��Pb��;b���2����c\�xQ��!�B!��7nܐX�u6n��m���P�"�:�hk������f����&�Jy{�4�|�����j��>JC|b��6Æ����L�8p �����&�#�HSh�+H�LV�$&&&��ʂ����}RSS��������`�o���Xa*MYYM�ӂ��|�E2K[��^FF:��;�a:���ر�R3$ggڽ{7>���ƞ9s&	�B!�BH;2z�hܽ{W�>ǎk�6v�.V���y��Ҙ�o ��%i"��]�.U3K[�f唾���C��L5�imm=6�t
�gͶ�p8x��!���/��uuu�֭JJJ�fK"x�c"M�SʼP�UO�b�|�ĉR�����X,Ɲ;w�m#�4��C4#����z:��;v�B��ٶ��KV/�2���$����X�-��c܋���e�С����fK�������ꫯ�B!�BH;���Sxzz�{��R��ׯ������ᚚ:�D"��Ь����Yb�'NN���fd2Ok���i��:��ٱ��F��{A,�^G~�,֯_�ŋ�4��?��ex� @��t����2#���'���Abb"�����#0x�`���Jl7k�PL�<X�U"+�8�%`߲�\ӱ�6k�O����~���f�����2l��'���p8DEEɔ?L$���QQQ��B!�BH;��ꊸ�8hkkK�';;}��A]]]�mX,>�pzjH>�
EH�*<ol�o�����S'�%;vx�f	��ێҠs���3�$�qpp@bb"����=z� ��U4Di� p P�d��=�p�F �U=�P(D^^�z�-����l0 >>>���C��Y7�.0�h��P�ʴ��9�����Mѣ�����5�t�t���D��������qo�M<>v�,�: ��?��e���P$<B!�B!�Tyy9,--1t�P�������� 88Xb����
mm��a*�͂��q����ս{�މ��,b:�����S�t�oog�]�
+p�x D�����ٳpqq�i�>�@��4_������Zi���m�[�naܸq2�Y�~=v��!����1��a>�	Oe�b =� �^�4y��k�Lǣ����ٕEѿ:w��������^;qѩ۸��"&&zzҿ�\.z�쉢"�l@!�B!D>fffHOO����@ ���'���%����	kVL�&.� �/'�東�����w�;Q,�u�̴����N�FhRz�jl�a��s(*���n���8z��Lc?|��*Q�. ��c2M��O�� ����ɢ����{�ɔ�z̘1�r��B�M��/�Ё=5*��,`nflmbd�������/�^?w.Y-�ݭ��w'�11j���i$GO��p;4��b$���ֆ��?�v�*�����T$<B!�B!�\CC���1m�4����l�7>>>��xͶ+.��Æs���U鴴�,+���ƒ��\��GF�>b:&M!�U�3y����e�N掚�v<?�z��M�eJl��䄋/BWWW���x�����h���຺&�4�}�x���C :�����2]o�p81b||| 4�AY^Q�X���S�m�mia20/[�Υ�}iTLz�N3���Y}ƍ�����a#}�*��oYE8���wA�n�
///��NMMŒ%K ���B!�B�FLLfΜ�N�:I���������.-� N6��0Q4L����ձ�0������~���
���I���VL����m����h�:��1�'���A@@ �u�&�ؾ��ػw�"�ɢ	�B���� ��y�G _�c"CCC$$$���Q�~�v�ºu�$�a��5+��_��fJ~ayYYy��^;�t,��Ś7z��9ǝ��r�4�� PS[�~9���� ��Q�p��mh��o�Ř0an߾�h��B!�B ���QQQ2P�ٳg��������anf�H�j!���U�P�شx��k�LǣN��6���x�mg�.L�"���<���J�y�7mڄ��N����������rEB��> �k2MD�ϙ�y.w�lQN�:׮]���X,ƴi�ZL������?��.v����V�������^���B�M5���3��jk���h3H��N��_�\�ӼR�����[[[��?x� ��}EB$�B!�B^�m�6|���2�)//���;
%���dc�/?�}�Sz0I(!;�8����v�a���Q�WO_bjl�}{K{�c�VQI~��'��$�1b�޽+�AG x뭷p��EB�E�� $��q�b�OM6�y�\����âE�d�SYY���#++Kb;cC|��<��vP$D�+��yVTTy���z�ێq��G�b�>\=mIGc���[jl���������%�c�ٸz�*�L�"��EEE�ի���	�B!�By���>���ѽ{w�����c̘1��K;|��L����/��@~Ay^U�-::���-b:&e��^mPV��M'k��,;jn��ר��c��?Q^Q+����5=z$�A��ׯ�T�@	v X��	5Q�Y�S=<?�.})kXXX %%2�{��F����F��l;�㋵s������J���=�+}$7�:p�*���c�ot��?�v2�i��H��x�q�|(n�Ʒ�����_˞�iΜ9�x�<�B!�B!-?~<n޼	Y��۷�rF�!.X�pZ�ٺ��r������Y�پ�r2�����f��hkor�����������	�}�Ed?-��N[[�n��ȑ#e������yyy��)�g ���&�h�o	*�5��sW�ٳg˵����w�}��v=����{3�����s�VUS�X\\
1~�y�r0��H��/�Ꚇ�-�;��dcfٚN��[`p.�?h��o��K�.�������X�t���B!�B!�ٳg�T����l�2�����n�āxs���i�()��(���724زeǙ4�c�d�ǳF��/��Mǚ�v0`:y	�"8z�I9-�ݽ{7>����X�t)�?.Gtr�
5���t�wEP5� d�Rׄ�ªU�d������-����5+���+N��>k���T%�7��v�0��$o����R����7�9�%�f&��&�x��ow�p�ϖS���� 22�Ʋ����B�~��嶉�A�B!�B4������лwo�����cĈx��q�mߜቩ��F)��喕�D
���t����3Ϗ?.6/̮X���;�ƪc_��#q�"�G�����-�]�h���d���ٳX�`�<�ɫ��JuN�����ҽ��l%144ģG�гgO��	�B̞=-�د;V-�6�m��]Yŭ����7�But�n�spY��/u����ۛ��Mrƭ����516t��21o-�O���	|OނX,�v������e΅'0j�(���+&!�B!�"5777DEEA___�~������*%�[sGaܨ�򆨑�B�*j*kj��ywM�uM�<����b�;��<���(����mf�����ب-n|A,~?}�#Z��3b�ܼyzz�e*��χ��;*+պ�����9�&kC/Y��@m�@xx8ttd˷��r1r�H��ŵ��s��,����I,��������������g��Lh���u�sll,�:v�}֤%l�o���yB���H�f�E&)Y����"Kԅ�f;hs���tu�t-�:u�p�����E?���߃ I^l���ǭ[���)���������!B!�B!rY�nv��!s���$>555۱X���a�g/yCl�"�������W�������"��)Xx������`�-��#��,>�#�
���<�zn�qNi���/�*���lt���v��ն��A����Рm�[=��w'��zyݺuCxx8,--e�C$a	�s玼a�#� ɕ�ۑ��*V�8 ��9���ϲo������-����ߝ--�<!�6,2:>܂H$�@9��ƹs�0g���		����!
��B!�B���B@@ �M�&sߠ� ̘1���,�5{$&�q�7L�F��b�������ʛU  ���{|��w򄨈Y ��{RM��{�F6�~ \�5axx8z��^�d�	566Ƹq�p��466Jl[X\���2�ۍ���B�'���wZL# ;w�Ĳe�d���� 'N���B!�Bs��uxyy���T�~ݻw������[l��$`=���&icD"1������)-�544������.��MPPV�Z%�����_uN��	��9H [�$!""nnn2������I��Z����kVN����<a�6$0�.�K�O}������oe����cܸq�w��}	!�B!�e�۷/���a`` s߽{��O>���I�0{���s�������@�&d��VGG�.]�ԩSe���ӧ4h����	S^B �$�s�րN�7�
��Ꚑ��!88�/�� �����s�εxũ��	I9����z��'m�H$ƙa�v�T�?��S���r���G�r�%�B!�B����999�;w��}�
mmmܾ}�Ŷ际���w��`�)�@{TW߈�����墻ZZZ8u�f͚%�<����2e
233�	S���{�ր�%� 3uMXQQ���4̟?,�0;::������?[̓]�m@��t������컺��j��q�'Q�R�_�f���#�� |}}�:O!�B!��JBB���1t�P���5
<O�[�y���.�{Ghks�	��Re�ر�r��Zl���???̟?_��V�\��ׯ��WE ���ߺ��w��x~-b1Ԙ~'%%<�Ǐ�����3��뇋/�xҽ�����48�[���D�pI+RS[�]�� -��"�����}��ɵ�P�TB!�B!��͛<x0���e�;~�x455I��^^Q����������JZ���"���*���ؖ������X�p�\smٲ;v쐫���eb�ր�[��ϋ��ͽ{�`mm����ܷgϞ9r$Ο?�'��@ ��Gi�p8���	rb&�DFVv���j����عs�\�홙��<y2jkke�K!�B!���H$+W0u�T�����	���Gppp�m����.�t్}��þAhl��VGG�O�Ƃ��ܹs����]$ ��^ݓ�&��*3 � ��9)��A@@ &O�,W����c��騩���}�>�X�h"��)�{[� 	���@���_~�%�n�*�\���6l�����O!�B!��K�Ν{{{���߿�1D"Q�m�l�O��˕��h.>_�S�Cp/<Y���p��k~����ĉ�ب��.5 � H�:����n�- pZݓ#,,}����tt4�O����R��w�1Ú�Sacm*�|D�4�����]DDK����fcǎX�v�\�544`ܸq�����?!�B!��n���C�����Q����-��}a�{7,y{<xl#�*jq��u�����)._���#G�5_zz:<==QQQ!W�p���[Zp�� o�{R+++����gϞr�������ӑ��"U{mm�����Q�b�{�[�#'nH�BFOO���r_e����3g��O!�B!�0e���

����\�o޼	///����v��w'¹[g��#��QlN�����&��;::��իpuu�k����9���r�WP0�I Ԟæ���T٘� �=#���#44r����9sp��]����t��E`ll ל�b1p'4^~ u
sss\�t	#F��kN�P�w�y�O��!�B!��'N���?tu�+n����3f 77W��,�F���Y��Ѣ2��Ic#'υH�Q  ��+W���Z���eee=z��j��
�;�<&&omh�]v��������*W1 hjj�ʕ+���'ucC��`�{;�5'Q����~�6�2�O���ꊀ� 899�5�H$����q��q��B!�B!�b�ܹ8}�48�\����1s�L���J�Ǳ�5�.�N6fr�I�+%5�����J��}�̙�'N��@�C����;v,�������X*�m��.�	 OuO\YY��� ,X�@�_P��9s�����nݒ��GSQ1�x�_��m��G��4�H$�x�	Di�t)d ��7�D@@�ܛ8 ��G��J�E!�B!��KIIANNf͚%WaSccc,^�999HHH��OuM�����ܭ3�l���$R�oha8{1�<����ll޼��탎�|kj\.�'OFLL�\��������5���������7o�D�����
����Q\\,uC=x��!���]�����S��.� ZZZ���o������\,cݺuؽ{�\�	!�B!�M�p�B?~\�� p��!|�����[���6fX��889�0�(_TL:N_�� u333����2e���VWWc���x����c((�  ��'�� 7 Q ������7oބ����c`޼y������C+,�3�;�=7Q\]}#�p',"���*,,,p��)L�0AB!V�XAid!�B!��Ys���ɓ'�>��w����w����03� ��DqE%U8{1I)������8�<�O�\ZZ�ɓ'˔�H�x �x�T �-�+f ��+Y׮]��ݻ�=�@ �?����B)l���$�P��{	�r���U�_7n~��w����=?��âE����=!�B!��L�:�ϟ�����-��ʰb�
�����OG����`����֦���$�!G��U�Va�Νr�k���bL�8���r�� 8�d �-�+�W<2���7oބ���B㄄�`���RW�~AWW����1���O��UI,#*&��QR*}�v ����?���>�L�\p�7o�]�&��B����vvv022���.���O���e:ME!���Ӄ��������|��ٳg(((@AA�T��!��;v,._���?p(���~|���hh�>-	 ��c���ܓ�XS�B�p��c�9�������'OV(���,L�8YYY
���? ��d �-�+N�- #�
���.\��ѣ���k֬��ӧe��1#{c�A��db1����+�"e������+������_�8JKK1k�,�S�&&&8t��+s�������d�ѣG��?|�{��aϞ=��=u���_|���˖-�8��3�x�����ņ��e�����?���a���J����W�^�9s&&N�ww��~���������ٳge�\��)S�`���/=�������C,���${����?��O?�����077�i�P���ڿ�;??���x��	�>}*W섴%,Ç����1f����5����؈�"88�O�Fzz�\s���4�\.�\.���������$&&��I��E<x���/=����ڵKm1BT�_�~P��8 $''cѢEr�	�07Ɣ	1£�lZ�S&�@�����H�������7���#G`ii�P>�o������QP< O ��A Ђ����y>#���*HGGG���ﾫ�X������'s_#C=L�c������±�g"�1q�~$�B;���������===�b�����i��������aĈ/=��?��o�Q�|.\��o���cs���ŋ_i��񠭭�����կ|����>�۷o���˗���GΨ_���St�����лwo��MH{����9s�`Æ2d�\c��b���k��?~����իq��a�b����t����SSS���"�Onn.���2? �������8x� 


�6.!�ŬY��i�&�����?((7nDdd�L�֯YD��    IDAT_�_~�E�9_�ٳg

¡C�p��M�m�������_y������\.՚#�-�ܹ3���1`� ��ؾ};������({6f�2q �w���xWDc#a�I�q;5�u2�733Ö-[�z�j�c�t�-Z��zF׹� ��d��V*G1 /</&���%K�`ӦM
��1c�v�Z��*=�kĥ�|��~g�J�Xڣ&����$�ʵ�޿DFFb�֭
/�?x� ����z� �=��c���+�ޕ���ӦM{鱒�(}�۹s�R�!�1`� DEE��ٳr/��O�Μ9<��Çahh���~�嗗6�Z;ggg|����������������������.]�{� &O��`۶m/��S7###̝;AAAC߾}U6׿o��СC����'��(,,��ѣq��U���p8���/����q���Gq%����/�}�������V����?�!��t�.ݗk����O�<Q�b��={0w�\��Ex�F��D��� �Z&�����Ʋe���!�'�ڵw�ܑ�D�?��"95O�'Jڂ��j��� _m<.�fEǎ�g�DGG+�� ���7n�����;w�jkk_z�k׮>|���Z�p�+�;������J���LLLp��1�l$B����#22R��`b�UUU۱X,�\����{)}�����q�ȑ6�ޡ���������>:wf�"#!j�����W�bѢEJ��f���?�ٳg��p�2�"����H,Y�D�cb���>��{�)}NBs�={�ٳg��_Ux�nݺ!88�9=�ע���Ƨ/����R��2�H�(���o<߬�.�fE�=p���={V�2|>~�!֮]�	�P�@E����O>m�o �P^d9?~���8�<kԨQ������6���T��"��b3�(6��0tP���f�iK!��� 	O�� ����;＃��VVVJ�K�o��?����c�uuu8s�V�Z���-½{��:׿����מ�W�	&`���j���*���۷cݺu�}���#00W�\�ÇQ\\����?�[YY���	3f���Y�^��ޯ_?bĈ����T�?M�8�W����GYn߾-�K���6���бcGI�x8p BBB0~�x�r���~��g�;������p��!11�����311����y�������s����-[����WFFrrr$�166���!���`cc��===������H)e/̛7�������WW׿vwwǰa������Ia�@ �G}���p:tr��b��z�j̟?[�n�Ν;��ɖ@�����!q����V9�C����v˝ہ��&D�f�Nh<
�*��cǎ�ꫯ�駟*�dii)�z�-ܹsG᱔������h[ǐ4���Lbnn��'ObҤIJ���
?���\o���f���l�A�ѿ�Ky���"���!:6��Y2W����c�b�Ν
]�����xyy�6e{7t��WrWUU�S�NJ+�իW/$%%���ݻw_��e�p���}��Qha�r������
[�ly�q�H��'Ob�ƍ��ʒz�Y�fa�֭�͇~��A����-��\��\.���P�Qe�p��ח�Ɵ��1<<<��;����~����x6L��	B4͋�U�N'y��y|��Rn=z4�=���0����СC%���r����غu�T���]���ӧO�'�|��Ty"��gφ�����J�Q�F���_|�e˖���~��	�
�B4_�~�p��y899)e���4�_�^ᔢz�:p��A���ͥ8�R|1����؄,D?NGrj�B�O��8�m�6���������EEEJOA� f�|M�H�R�(��
<O1è��
L�6[�nUJ:SSSlݺ���X�h����_��HN���nc�7ǰ�?�E$����~y��HH������� 2E������ի�}����CBB0p�@ZloFdd$���_z���S�LQ�K�.}�1&N�SjB4i�$���{��2�5
���L�� p��e�������<�z�j��"�С�=�*�;jkkq��,^���'O^iӷo_���V6lx峽������^l��>|8RSS_z��ba���J��%B�)))��_��쌝;w��]��f�ĉ���Sx>ggg�9��BCC_)t�����#�h���X2AAAJ�G����Gpp0<==�������T�z�*�s>#6!MM�OU�.��QO^�7'$?�{���ba޼y������Ǖ�ؾg��;VS��ZlW*ZpW�F o `�ʤP(��_�I�&���@)c:;;������X�x�����!1�)~?u_n���m�q��R3
 
�/S��+q�N,v�u�9���p/<u����wss�ٳg�JaMy	lڴ	�Ǐ��KU{�����c��u���o��Xuu5.\����e5~�x�X����	i�tuuq���W
��������ߗ{l���˗����/=�b��q�F�������KuZ^�%$$����?~�e˖aذaDE�j���`���/=VXX��?�X�C;%%%X�h���,?i�$�Wnjj�g�}��k_-�ebb"񶟴�-[��&�g��ʂ����kVBچ��
L�:�~���n?�?<�͛71x�`��jh�!���?r�>���.!�V�+�Nm�	�B2��p�j~��,6|{>~��K̆@�ؚ҄	�s�����M)񖗗c���X�v�Zj�I��4 5L��Ђ��T ����@  88���Ǖ+W�6���+�?�G�a��
C����r�`�ދ�h�A���Y���G�xV��B�*�D"<�+��8�	�����-'q��=$���W|�`РA8{�,�����奴Ӄ���9r$���_�bD^u�ĉW>@͜9&&&
�=iҤWNZ�����Jyrr�+�m߾]�_�	i�>���W�$755a޼y���Tx|�H�?�/=>}��צ^h���;�mۦp����`�ԩ�lD�X,���E���y\T������.���
�r�����&�Ӑ�.h^
�LS13\���.Y.(�y�\�J�T�媨 X�W�M��Af���1��x��� ����y��<��,���<��svv����-::�NK'%&&���Ü6�Xww�Z�Y[�lAhh(�}ҤI�ݻw���H$�eb~��7�����իHKK��,  �A^D�c�6m��������~���q��e>|�N3�+�
��}��^���c^�|���������(/7܉�ee�HI��c�&`����t�.|��G�8y��?���b��ƍ��˗q��)����r�ԩSx�7p����YGy ��}�i�覩�u��3 ��ݴ����`�ر���Ŷm�`aa��~{�"33��=�oߎ�O�ֹߊA�{�����  kK���A��l`��-^kg[[+��ύ@�J%����qd��AV.������N�UE$a�ȑ�7oƌ��������ﯓ竩����ѣG���]�fjj�	&`���u��՛�����ҥK�a�κ�VVVسg���u�4!�z�����3��ח-[���D�'##[�n���P"����7nԪ���`|��W�sG�����#G6�s��Ǐ����������ѧO�3�	ihڵk�k��Ȩs�Ą	8m}�����ڪ��G������Z�<5jڷo�i{������s���ҥ<<<p���Z��0\�v}��EHH�̙��/�D"Ǝ��c�"11�7oƁ ��}p\V�)�����w��hۦ%��l`����Yî�5�[5G3I��_^.GN^!���AVf��aVr��2#����'O��ŋk�w����ʰb�
�_�J��Ǎj��h���!z@��w�;��T�z�K�.aǎ6l���upp��u���;wb�Ν���?u�? ��!/�I�39���`kckK�ji	��h���-Laan
c�f0qsV�f�^�
����x�d��\�T����R�>�"/����(x*��d�-���s����lIW>|�ٳg�7�JXXg�P-+S�@ZYY��w��]�rׯ_�u�ڒJ����Gll,�C�[o��3f`ǎ�V!M��ɓyk�޿[�n������8Z��#�J1m�4����e�F���?�۶m�I�B9z�(.\��[F��ח�I���K1���JHH�����2����d`��d2����i�8q"f͚U�+
���8.++���p���X�r%�s�̙3i���&@&�a޼y��_��w����Ag}���`�޽X�|9�n݊}��!??_g�+�Jd?�G��|\�����E"Z�����l��ЪesXX���]^��بLL� ��F�HT����Q.W ������
KKQ,���X�bi)
�#/����(,����0}�t��>�.]3p�A�k�B�v�w2'������DD"���e���L_�^����������oC���۾};+..���T*YDD����wm���,33���*
foo_�>g̘�{�4������


j���O?���Ã`۶m������u��Y���޽{�>nݺ%�sG�zΝ;�{�͛7Oo�;z�(۷o���X�v�j�~Μ9���y��mڴ�����"����'��;w�Ը���_ޱMMMu�8�?��ff&�D��f(���w�޼�wRR��u�S�N�y��o�`�^-�-���*�YFF��ƍӺ�֭[���2N?G��m�٦���N�)JË��9[�n����.�d2����鳉166f^^^,22RoωT*eAAAL"�����2��l'�Q	�7IB��8���c���z9�T���c[�neC��ɇ��'''�d������� %%�<X�߷�d�ʕ��x������󜾊������F��z���7��c�O����S(ڥU�V�����)//gm۶���T7�nnn����x??��V�※��+))�C�/(C���+((ཾ�/_^��{� ۼy3��7oֺ������?~<o��ӧ��y�P(������7n��	����ƾ������M��א"����Yhh({���^����ֱcG�g5��^�OH#� ���Ƌ��'�s�^O<�1���C��d�}upp`.dW�^���]XXȂ�������wcJ�x߆_�~�V}u�҅)�JN_aaa��w lĈ��cl�̙�E��v�����������T7��2�)
�6�|���0�w ,66�w�)S���P(�����c,::���ի�ꨏ�1c���q��e���y�&����\fll����ʊI�Rζ<`͚5�y�P(�###6�|�_t�ڍ7�ҥKY�.]������+۰a�ߦ���_����@R�{cB�! �A�7/FFF��ߟ�����d�cO�<a������_�K�j$	sqqa�����իj2u�b�����
��'O���_]�~V�^��gРA﯏w ��o��mS\\̜��4���)����_��sk׮���SӀ; Z�s����[2g͚5�?'�.boo�
y��
���l�ҥ���E�W��ǀ{�Ν՞������>��%�o�>��<(C�P�!���lӦM���寿�b۷og^^^:��dH���`^^^l���j?�Cqq16��U՚�4	. r �OmZ�n;��{��g��\.g.\`�W�f�G�f-Z��q�m���؀������ÇYQQQ�=���fD����84�L�<�����WZ�!�Xzz:��������׀����{�.o���]��h��B�.111����ɓ���h2�nnn���q��Y��u���O>�c����?'��2q�D�>�?~���߿�����N�:鴆�p�H$L&��ckk�q��=o��>{�9���ɓ'�)��qvvf�O���ܫKR����İ�>��4�A_oii��~�m�r�Jv�ܹz��1�}���������I1 w��� �¿�L���ف�^^'���$��w߱iӦ�~����W%	�֭�8q"[�v-;s��������<==L�J���yW�ܻwO��_#F��=��~��Vu�k� sssS���5kV�Ǡw
E������k�������ɀ; 6x�`�玹s��xCp�4i��O��9�Pt���{O�ϱlϞ=l�ԩu�h}�`>����Y�}����ӧO9�޼y��}�b1�����T*��2
�v��E�ο�RZZ����XHH�4i����n��^�����}���S��-[��k׮��$�
J��ޗ\�e
 !MTw � �����ՋEGG��R(Ց��,55�EEE�U�V1???6|�p�����ڴi�����&O�̂��خ]�ؕ+W\YRR7n\�]_Ȩ[b`ذa��ٷ����n�Z��9��mٲ��mqqq��H�w
E���������u�M��o�����T*e]�v���:�����;ƥK�N(]�gϞ�ܹs�׻&
;w��5k�֟g��pW����5���>��`���[�jo�����|S(Ê��'KLL��9X�d2KLLd���lɒ%lʔ)l���z_�V"���;��C�2___�:Ē���u�zU�;����#��D�dxD0̈́.� �� �A�̌A�u�&N��>}�`ɒ%7n$I��!�HЭ[7t�֍�3�\���l<z�yyy���E^^������s<{�J����(.. ��� `ee�f͚���666������:��ܼ^WM\�v!!!����R���&i׮]�;w.����gϞ�q_�?�����?#''G�5�UPPF��.]�T�YXX`�Νx뭷��:BKKK^[ii������cƌ�u'N��͛7k���K����]�v�l377GXX����ޒJ��6333*!D�n߾�aÆa�С���Ǆ	`bb�Ѿb�C���!C�a�|��X�f�={�窵��ܪ��yڴi�?��r���5�w�^,[�"������˗/�L&��؄������8q��� ((����}����������獻���A.�W��KJJPVV@��Gccc�D"�l�FFF�1�m���������w��R�DLL���K\�|Y�r4��@��ub, ��߂iGGG�i�&V\\,��M���癗��h7�\�r������k��ԩSy�mU�̫��g�U/-3{��*����vQ��p����G��Km|��U���w��sG```���w
Űbcc�|||XDD{������L�o__3����x�y��7k���ɉw�oLL���={�,︾���?�
�p����"""Y:����d,""����C�ׁ9�%���B@*I��U�B4����y��cǎX�t)����.�ѓ�d�믿����رc4��@���q�ܪU+���;5�7u�TΟ333q��i�֦+������oy�_�5g�;!��*��zY�UXU||<BCCy�k׮U{��!kժ�-??_�J�_yyy�����;;;���.����QXXX���:uBll,F�U�jF����ӧ5����Ǚ� ���Wݶ�Oiz���=z`���j��#�����^�;v���/����.IS{�P�_hD�h�ݰ( ��A\g����/��:t������ �˅.�QIII��E�СC����֭[B�D^q�����p�|||�ݧS�N6l�-,,̠�XX�h�޽�i377Gxx8�b�널�R�䂭�� ��ֲeː���i377��ݻԹ�eK�d!M	iLc�~�:6l؀1c������%Kp�ҥ*?ǘ���СC�E�H$B�-x�5�K$�d���|;vL�cGGG���7ޠev	!�KKK�̙3agg��� ���]R��T*�I�&�C���/�����������B^�5��& ؇r)H��)66�۷Ǵi����GGG�Kk������;w6�5���BDGG��׷����}�  wIDAT����U�~���8M
�{���{�uQRR�?�qqq�����0{�llٲE��i����ѹsgN[׮]q����)++CAA�Fۚ���}���R����ܹs������!007n���u��Ɔ�F3�IS�P(������|��Wx���Y�f�б����͛��ޢE�������~�m�������������弶�3g��?֪BH�TTT�;v`ǎ�۷/�O��)S���@jv��}���c���������(��H�!�!���_���ٳ'��J�JJJرcǘ��/������h��C����ӧW���;w8�;v��Ǯ�5�_ΦM�x�J�RֵkW�v��;��]BCCy�����������S�k���6��-))aݺu�lg�k�:t�w�Y�f	���P1�ڵc���=�co��F������#55���"##��>�PXXȬ���(JÌD"a���,""�={�Lo��"''�EDD0www&���4 �@Rù��i��  ��Qk�o�Fpp0�v���cӦMHOO�,����SDFFbҤI������"""h]��ܹs�s����ee���н{wN۫���ŋ��2��Abb"�����X�|9RSS9mfffسgg满ruu�%$$P	!��ѣG���DJJ
�g�Ǐ���Q�^�r�J�����b�ر�*	���5.GH!UQ(������/ڶm�q���������4�q��=l۶ÇG۶m�����X�^ҵ1 ��5���>T�0����C||<���''' **
EEEB�W�����m��'OFTTop��$̰a���������??~��Ǐ�4��XZF�Pp��9s�T!߯�����߻wot��A��t�biu���@���L׮]y�䕕�!))I��э��{��׿�_��/_��`%%%X�l����E'�ז�����/�|||`ll��� ���!�����d8|�0|||ЦM����-Blll��ߞ\.G||<-Z�~������g��ٳg� ;���`,����po8v �`? aK������u����0x�`�����������%�\.GRR����3g�����B�E�$<<�V��\T$a���		�������ޜ���٣v=OCv��lٲ�7H��_�ĉ���������ҥK4hPe�X,F@@��A����ŋ��o��g�q�W�^��Ǐ�2���-..ϟ7ع� P�6�sIϞ=u�eҩS���H$�lk۶�N��[[[����{��M�6�����S��5o���ќ/7������F7B$��R�Dbb"�֭[cذapssàA�зo_4k�8��R)p��y\�pqqq�q倇 �8-t!�4FV �C������X�>}؜9s��ݻ�իWYII���|�H�P���4͖/_����Y���<)��#G�p^7n�����ۛ�s�R�[�\����177giii�~���X,�5�)�Zd�ԩ��T~~>kӦ�^�W�k�W��Ԕ������x�"�H$����������}�_/J]���
���:=Faa!�����*����/���ʕj��ׯo����:���/���ݷo��	
��tbnnΆΖ,Y�"##ٝ;w�\.睛�L&c����޽{ټy󘫫+k֬������ ��q|�մB��L,Tפּ-G�
�]��k׮U�I$t������ի:w�GGG8::��Ύ3kF�


������ddd %%III�}�6-C�w�}�������֭���  �&M�l�̙;���S�NE\\g�����1w�\+#��:x� BBB83@[�j��7�����2ݑ�d�������9�7�|�~�����7s�L޲>����駟��ݹt������ǎ;t��֭yW�fgg�om��ب=Ǆ��W��������s=�w�ƨQ�8m��ޘ?>rss��?!�Ԥ��gΜ��3g*����УG8;;�G�ptt���amm]��egg###���HOOǭ[�p��M���5��qJ,�I�B�vh���p�> C�E�
RSS������(��LLL��� {{{�i�666�H$��� `ee�D���B(
���������999���E^^^e��������Oi�,R�'N ;;vvv�mcǎ����ann�ѣGs�oH7KU��ŋؼy3�ϟ�i_�v-o�fBH���ʰr�Jl۶����ルW�"44T���2�K�.a�ƍX�p!�}ժU�LK��ݱf�^�����Kv�(�>}2�����mC���ѣ��/�Թ�q����j�A�>�D"|��w�������`���U�gff�)S�p��r9<X皎=���\NM&&&���������?!��Fiii�24�������#ڷo�siݺ5Z�l	 ������1D"Z�l	�R�gϞP򗕕A�Tr�[*���� ##2��^wt��4�!�)� X @
�/q�P( [�n璷�/2 l�ĉ����fnn^��	��LELMM��۷k�􏖔�P4�X,f			���B�`���N�!���ٳ�T*�G�K�T��Ԕ%''�x�jI'''v��]^��=bVVV��N(]�������Ǐ��]�-����y}��ٳ�}����D"Q�tc�T����o�'N������2�X,��B�P(�E` ���H�$� Rg
 ���I�k!�@u�0c���@�0a��v���k3$e2�O�N3�	��R	___�Ub�!!!8r�jݿ��Ν;��[���ܼ���^��2�v�022���ѥK�σ��PXX(@e��ǪU�x7ooӦ�����;�ԪO[[[�����ޞ�~��iܾ}�ֵj�G���߰`��Ϯ^��]�vU����d����ݻw�ڜ����ؕBH���5 �kؖR���@�o�(�&��g�rf+-X��={���ֻwo�K���j�X��N�h��#G���JKKٮ]�X����H$��/+++����._�\������W�^U����y���W�{�����ԩ?~<		a>���-[����P��5k�T�����aÇ�hֵ��%[�h��������s֧O�j����V�Z������@v��I�T*��NYYY�C�������ۿ��P'W'�uW4���ς�&(
�R�y
`hbt�Ak�7>Q �0��m	!z��C�w{�/��VVV��r�
�_�.Diz�|�r�3ݻw�B�ӧOc̘1����? ���}�>��#dee�ܹsHJJBvv6�R)D"ڴi�Ν;���puu���q��;v��M�V�7����z���~���9W�������������?"00PW�bPV�XWWW���ۼ�yzz���YYY��?p��]<y�YYY022B�6mЮ];6����+�?��s\�vM��.\�3fT�scccXZZ�E�����///ܿ������ �8m?���ίNܽ{7\]]9mcƌ���=<x��cB1H?��ЅB4��E�M���bff�


��-��ﯳc�w ��7�dr�\��L3�)�ڥW�^,))���I]=z�M�2E�Z�1� �߿?+//W[_mg��R�d_~�%��Li�133c111zy�X�B���pץ۷o3''�����޽{�����u���lْ�����,�k�B�P(z� �[��<�T�qK �`*�G�BH�RZZ�C����T*���빢�q��%|��7B�AH�r��-���`���(**�Y�Ϟ=Ê+ХK�����Y������6Z�:qqq2d�,Y�R)t9��Uii)�}�]A&�����|x{{c�ʕ:�.u�_�~�믿j����;v�=|������k{��)~��G^��3Ь]�N!�P�@���xB�Z!ud @)���BiquuU;�j׮]:=�!�p�LLLح[�x��w
��iѢ[�`�{���:y�_���̙�,--�>��f�U�;�s��B�`���lݺu���U��B*���l�֭�^�W����~�zfmm��qu9�=??�EGG�)S�h}�;x� �����Zo���#��&L��@�P(���v �A=Q͛�F�3� | H���Fo�ܹ033�>|���:;�!���2���V����+�z�-NۡC����������1z�hN[nn.���t�?!�ٳ'<==����_NNN�ِ2����q�.\��_~�E�ٝUqqq���;�-**
�����e�z����'�-??;w�v�Y�f���R����r��� ���HNNFii����X������C�E������;;;��@u�IKK��˗q��)����꽤��
!�J������d<|X��pabb�i���DFFF����H$����y��߼y'N��GBi�� "����� b�h���r��G��wB!�Q������%�b1�������joJ!�266���E�\EEEt�!�Bԋ�9 ��N4p'=���m"��@!�B!�BH]�X�Ѕa� +���B � �jؖB!�B!��� �� ����ɫ��	`.�V�B!�B!�B������F;y��IU,L�)���B!�B!�B��x�; [ �	\104�Nj"0�?�q �	[!�B!�B!�N	�"� � �
[1T4�N���  p�B!�B!�B�-�A�� ��� Ѐ;�1�����\�r!�B!�BљR ǡ��~�\�rHCBLx ��j�|'�B!�B!M�SP��g EC*p'�dՌwo��-�-�B!�B!��*� ���Ba�!��}� �� � }A�7B!�B!�"�t��c���.���� (�/� F	`��?B!�B!��O� �d��=a�!�������w �	Z!�B!�Bi�ҡ`?��� ���&�܉���jٙ�_� =�Z�B!�B!����@5�����@��EB�Đ�t�� G /��	��`�B!�B!�}+�j	��� �'T��PU!U�w�P� �A5���-�� l^�9 ��4�j�1��\/!�B!�BHST���@ы�b�f�罒\ 9 �@5��Z�40�C�evn`6�    IEND�B`�PK
     B"BY�ʩ��*  �*  /   images/9a88a734-d46c-4092-86bc-e9f7b966a1ec.png�PNG

   IHDR   d   A   '��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  *NIDATx��}x�U��;%�w �����& *Ui+
(�
.��������R,tE����{!�t�{f�罓��0�	��������[&_��w�i�9�ܫ@���h4N��#�h!�O���6d�#W��rl��\.c�P�Đ���[�o���P�i���>(*.�(�:u
999u�B???>_}��#����!��w��d�g��?���˗;�XN�[ޗcAu���>4��4>}�s���A|\4rs2���D�N���Ǿ}���PRRR�~�70d��ر7n���
��9���	I�V���cʔ)��@�JKAJ�M���5���Æ�,^������収������˪�SCf�1mҤI"͏ bӷ��f!��;��`(3 .�
��C�����5�:u
nݺUc�ƌ�aÆA�բw���3		������v�>��?�t���-FƭTl^��>���t�P���c�#��/��":v��>�l�0#_�Z�]w0D8�OT��Q�F㡇����&pr�Ei�!R�q]<<��C����#HL���%_b�c��H�ӬY3���������8w�F��^�LU���lٲ��F�>}�����L�?]�tARR��D��� 11����ڵ+Ξ=��j۶�j���U=�w�^8;;�^�z�~���͐���U�V�][`ێ��)���E�O�(�zw��((+3��˙������������!�0y����믦��r�X#Cd�g��?��SX�|��l�צ��������Q�-�l�׽ۼi��+�by�"^x�E̙3[�өS'|��((0}x||<���� 6jԈ�QZr��m\�tI�]�����`�СX�p!}�Q������V��'CZ�n��5j�b8��x �����M�6U�\���f����۫�|�._�Gn^a�5��t�2�M��l.--{5�e�+Q1Ɉ��j�����₾=[5���2<6�E�ڵ�b�0t����tUeH��Ə��#���u3_� mnaa��^w�I���<��̅���/O���3�˚�5���~�7%�X�j�w�L��$�W�X�3f��TνH$��k�Νj𢣣�4�_~A߾}�V%$$�{IԀ���C�b$5�G����UZ����M�6a����t��e��)3t��5 �:O��gl^�����?=����[��g�+��ps.�j5EE%�����ۇ7�޻{��8o��z{aFWi�@u�EM��kѵc��i�"��㓧��O��'f��/N.ΪR�2QVj�%64���[�8�.]�b�֟Uc�f�B@@�Bg�`��S�⧟~���#ƍ���O�FiW%���ܹ3�]�����5$<<\i��ŋ�&мyyy)mb��8j۸Wt����������=�TaII�?�]������O��w�s熜܂+%�es=<\g_��B�N��	0Գ&�4���P�՗Q;d�J�Ҕ���-����0������DH���۷sNx���KdAxl���tL�0A܀����+@�ҢE� J��ٳ�e˖��֬Y�$?""B���~�M1����W�\Q퐙d$��IS��xNP�mۆ?�Bڦ�$���E�b�0m��Ksߛ��[���s�kx�����{�hoK��;����������{�X�Y�!��A��1�3R�$�Њ�ɭt�%[�ڋ�����i�N��A,�Ar�t�@Ϟ=q��qN�O����o��6lؠL�%ݼyS�����L{��:0��իW+�\Pc�L���	/��������Y(.)�`��RR3�@��\��^���0Rh�*XU�98:�N:ĠM�^��hN���t㜷&H�6X���v�C�C
���쏘ؤ�{�\"+�(�ڵC����oj?��]��Kt�V�� ;N ��ѕk7��|��D�&K+�#3�za�A$~Ů��Č���;ڼe���#++���2��ɍ�����/>�";Gl�����v�� B����v]�c㦭m��j�J���y��w����A���[�(}��ӧ�o�O�	:�N�:}�%�͎���;yyypwwW�6�Q\���Y��#F����������|�w3^�B1 �v|}�i��*�O��_��JQRf�Ɩ&�*Y�y�DӃq��f�i�?&.�}a����tA��h5HK�U�J"�E�2�Yy�b��e�NV���ٺu����8|��r�DYDk԰aC�9sF�:2�E��~�w�ׯ��:AG���ѹgee!88X1�h�ϤH�&���"���g����^0㨽��8{Oe�=��de��`g;Ⲅ����d�-���=eZ���hР�kI)�	��Rl`�L'��@y�4"�}����130��J��U_�������c�̙�aֈ���!�$��)��^##�7(e�����I�QԠ�/�?A��[o��5+�o��>��6;EP�wl�#K�,H�D�!)����sF����3��Wm.k�̗���e������D�������r��Ek4p+=�.&a��4�ٳ[=K/�L쪣�'��Ʈ}�*ڦ����j5�*,o���5"0��$�Yc����	:y�$~`2�/Æ�KЪ������L�V�Wc�~\���"7�5�>;��o��!���&>��>��y8y|��ٰ��h������?�U��88=�6X��ҕ��b��>��lN����3���L�O2�L˖-EvN6&N�;�ُ�'/I�PJs�-.�o�:�M��+�Jd�W�VG5��ɔqO<��C�`Р��SXT,h��l�uќg��73nVz�������[+�\��[���6�_����7����^̫�d|߾��IU�*YK.*dD���Qll,�H�ƃ6�g�p�)�P(�a�v��p����	��G]����O��  ��1�����ԇ�J�T0{dTJ��z����d&I�0.]�W��"kܸ�u!�'���$)����D�&��;	���jKw0��F�4T�����2���E�7F�	�֭��g;�����䌷��A��#X�v%.
C�^�V|�Y\�9�&�ٹSS�������M�#>(YL�^T܈�����s�7Z����V�`��^��7�|�͘�~�����k�A;
<���S�����$�׺wig{�&���Wga�uzswwCw0��=//G`�	�$'Se`��)�PT\RP��2��]i�|��E˶��wɽ:���'O_D�H{�h�N� ;{�����N�h�K��b꼥�I3j��:}���3���I�C���ʞ>%@�Μ��ҩ]�t^X��ؿ�^f���B������ ��w2����}E���jLy)����=~�t��F";�8����Q�e�L�Y�q;>Z��Ԕd\�xFⅆ�'��/^��D;j0�����X����1/1ԥ[_t�>)h��W�A��#��	�����(4���Y<2�Y8��b��t�\U�@```E�.л��;��_�]�Ǘ_"XN��Qbf��01����psu����k��8�e=J�8qFB�U�B�/�1�c��_?�j�]{D�mx(z���۴a)9i*�ИP�N���SڦE��H�<��k�������6�%HUflæ����兵�) ��냟���T�g-k�y��O�p���9���%ތ��G+��4������c��!9E�vT�	d�4XL�s�#ZTycġ:w�ĉ*MN��y+qQ��s���[�X�ɧ�J�{q�I���pr�8�HI������!�s���E����m�7���-��2?�Af`j�!��,�9�YWz�!oL�����ƻɱ��by#r�j,Ŷ��بY�9x��ء��H}lI~*bN��d������cԜ�2Jr-!1C�)�<sA�-!�����B�kRS"�fi���L��>�w%_Y�x?���q�&@՝�����W�Іɪz�գ��e��1w���U?��������NM3�"KSV5�)++O6QX�`΃Qh���Ei'�3��<=l}���<m96�뚊�w�;���X��G%X������p77ԡcO��uW���d���$��̺�"��r��i9[Vq?�*�S�A�,!5]�D���q��i���`��#�z$�{�},Y�G����h�B���ͫ����\UP̺���[�^AE߫Pk�׋�h�`Ҥ̙S�_�>2���A;C��yJ��-0X��1i���`=�ή�<g��̙�z���qèQ#q;�&���_�,�+N���O�6^�L�¯�Vj'$���:��%�~��&� ��'"�r6o�U�D]ށ�7U�Bԥ툍�"~-�~Y%��;bb8u�Q���F"8�+�<T ۻw?1��x��Y*��ƌ���Ʀ�W�a��>��o��ݻ�o�0aE���0�A!��4�A�_M�jr�T�8An����T:Q\���^cQy������)�w�S����.���8X�b���Rq=�
b��U}		iʄ݈�Dr����W���B1k4sj�NG�+f��D�������
�^k B�2���TP��.�w����Y�b�X2�M��u���ݍ��/rԮ�wb�`���oW���jt�T1Y���CZv����u�pա��\�� גno�;����>@C?�*c��g
�����}�w�`0���ZM��?��Q��歯(�X�a�����}��">�f��J��2e��ଜ�AOu�є!?����A�Ӎ���>d��Y
w���1�����VX�}�*3���8g�GK ��9�̀��������F���ġ;QT�(ݨJWCB���hP����ExSah��r�T|c�����)�S>|2���GTt�z���T�%z,��U狊L"�����9�кec�m�T�����OSS,{�K�2�6;�`�K�Ȑ9�,�f��r�u)�fmԺu?Ht�"\�k�OE��׈�T� &�f<�wU͘���
�~o�E���0sѵ[wU�ǪKrt�Ep#_A��0�H�[$�":&�#��7�dD�@#�#q����OO�V���?�m��/y�<�2]�%�������V*M��H�p"�1ʙ�t*��	�����M��Ŏt��R"%�B
�n#;'�^f�;�d�FANK�� ����@PkR����Uk�c`W:�����6l�3 /#7q2r�fk	��{E��Μ�AT�:��;))g�+*:QM׍�>c�{����@�(��C��}�}n4~�x=z���Ř��}�_���9sZৈ;RPm��=�5'�+�G�����ߟg�@ػ�@ڵi0�G��2���M��W+5;�E�lÑ�WQYF�5����ɂ��WT&"o�������� v�����[�����`�r�  M"�W���ե����w_9RT�#f+���[���n�$���T�!�()HF�`w� ���"?ARf>��j�v� �꬧=�	�9R�66��׿����=*���_�asg�Ȟp�l '�����Qi���_U�Nm�bh+*���d����@^_��/��C��)ӭ]�_��S����!,^hԨ!<ݝ
ar�ێ����@A%-U"QW���-�˭�� O<1����W�fȸ�\<o�֑I!���C`1w��6Ĺ�1w���������P��C���pķ�?�6�կ�o�􌳣ڶB���h*�\�̬|1��T0Y�0��N�~�����s�U�]+�"PA��}�ȑ�$�uC�fM)�L_���p�F�Q*ǝ���zH2ea�Vl�(P��Pj�����b܈M��}>�ݥu�"D^ꤣ.�ˢQ�W���4An9x�q3f���dA)3�ο>8����-
��gJ4��ν�ɩ��j�ў]�jeP�E% 9%�����-���"�:B,�z{���Ѷ���0�v+����ph�Uaa�*������>�l~�%�>�N���CGbȠ�X0�3��i^|�U�S�nJ<���� ��>m1*rJm�g�B�(Δ���y�q��j�:|��G�g l%�/c�w��E̘����J���/Ŕ�Lq׈�ͪ<�<t���ml\\�]_�%b|�h�x��C�PkL�i�pS�}�������F�����K�1q.\�UZ��,�I�D�&m(+V���5���ļ�(R�
�������_W�{,���|�9���^}�m$&&)��<�����d�||:e�vX:s�p4
�/_���)i��e��^��e�$���q� ����X���7��R��4yhѢ��^�xu����-��)M�a!@Yi!l�U�$_ ��t��Lp��H��Q'ƟǩC��Wo<u�{$�������B:��h�*|�f��&?Fb�������DZ#��H��T������)�}u����.g��i�0N�믿�P�����駡�=�(@ki���}s�Sͷ�M����������K�n�\t�X�r~O�sY��DF���|zF���*�MEq7R��~g�$�)	m��VZ���젯�/:u쀃w!&6��3�7��֜5��U_'N��?�����JcSu��i��DSN!�L�����h���}x���|X����;��e�݌��������\B�;�3a+�L�i���g�a�yʟI}z�B���)'��m���pw��a]�a����)��,����N�w]R�&2�ı}��.a&�Զ�Y�X�RU;,���QVn�,�:� h��47�%'���k(.5���	��5����ܜtU4���#���UɆU��%��r����J>qxp^z�e%�bv�/�c�>���?���yU�Ú&T7�X�����Uo'CXm��l��\O:����Ŝ�����л{Kx���hq?V�}�]�TQ�sw��}�=�C��"''��<U���`y������Mp��	���µ��ѤYc���u;A$8k��XX1�K����غu����*.�G�bj���>�����jKL��6i @!q7�,/�!C^�	R�����_z8x86��{��(�R"����,�SL�U�Z�i�k�$���.U�Yeʗ�>�C^�Y(.�f�e�n�A��pt�A��O��p��Q4p�ţß���^����rM���p�,דp}bm��\/��Y���DKn��EA^ܝK/��	.7����Z<uEB�_��A��H�'s��Y3,pt(����th\�[z�{]SU��ұq�^7V�M5�*=c4��T���\2��Ѡ�Q9e����34YL�ԅX\�r��
Pc�P�:�A�1}~/�+���z
T�J���	*_��Ӂ��XAaa����~��6�ɪ�����j�MUHbd���`��x�S�`A2a�QJ�N��/zU��,:ȹ�41G��?�+��E�?��b�q���;�$ �V� ���j��7jJJ�<s�.Z�v��B�bE}բ��<9s7�B �=s)pfV.f�[��|L����BB�In:�<c>�^������ީQغyR����ŕ��Yt��{��;���~������=Y���Ж��m�=EE��&=�@���ΒY#.�{�ı֊Μ9*��ة�rtb�0�� o?pZ��VSޑ�k?
�t*ٲ@M�)�#�Y��5�\�2�vd�.Hd�j�ʊ� )�F�_�E���r�ڊ�TVMǛ�G鿙X���!m۵��>$�|}Ȇ�YbI\%��ǟ�����c{�֫T�\A�dɗ�VPQ3>[��ҔԴ��gr�ws��������Dܘ����-[�T�\N��7�B�lnP`�bNEHH�Z'�~���ps^e��I8zd?���μ�
�T����F�����|w+����p�z�Ih�"PTЇ�,�&��0h�D��{���M��Y�W��V����#��&�8�Yٚ>�j�rC����ue����gJ67+`�&f<��D<���V�|еCCeE`��0��v�-rS�&=;u����U�j��떋B��~+,*��Pf��h5N��zy�O�������_�U��Ν��ݻk�y�L�\S�:�'�8�*Q

�^�K�f����ի�j���GmNP�US|V�sW�nݻ#33K��L.�;yt��*\2"O⩅C��$YZ�&H��Nl�<hHJZ:6�]��>�X��X�G��n�D3E� 3
�?�������8]auڃE�k�lm����40b�*<3e�U��|&48@!���س�MN�EM`P���6��`��;�iGG;�����tUp��l�6��5/��ֹ�@oWdފsh]SYNԶu�B��.�4:�wR[EEG�sǦ��p8�Dm@S�L�>Cm��=ńi��%�����Ԝ�V���NN���s
^�������X�x챱��֊!t�'��Vf����gVTt�����uqqD�@_�tQ����nN�()�Ę'�HO��I�+A�׀�m��/�@Bbz9$,B��!�4n ��Ӥå�����n/�8_��?7u(�[(c�,0�1�Z�]J�	c���z���]�:-X���߫!9�O�}�v�q��N~���Ɓ×�u:a�sS��a}��#)�5>p����Q!�>�>A��:z�Iul���l�����Wa ��"D���Ҥ�������{�v��tss7-��������2c�K�+��������mϙ��u9P�3<.&m۶�`5�_�62�/]�7�Ip�&��7�ޣ�7���c��"�-)i�������}��aݞ�]z���T����$�m�>v�TϮ-��z_�o.\�ՙ�}�&b6ZC4w�H�a�����4bX�&_|i��rqv��Gzp�؏¤�"_����u{A�afy��C�"��o<�w�lԹ.�N�w.�9z�T��m�n�Gÿ�;wۻ!�nb>yob������Avn>�����)H�-��n�Q�!U�o��(tJF����⠸��%���r�zi4;g$u]4<#=K��L4S�&Nm~���J��l���-s1��ʎz���Y58O4$��'�����������dc���~��l�wlJ�B��saM�33$��z������{�hgo{A�Y-�������y�b��g�ۦ��oǱ����� �%�k��lN��`�@|�}ש��BZ��J���,�:���b���Neɧ@��mo49��������!�DZ�O�yN\��`�írQ۴Ƀib��C�h6�z[���^>C_!���������y��mX���0�1*Uo'>`�A��7�-3�9�&�ζ��
�--����}�8����`�G���'��8�Pa�5/7�k��p&-I�y*�G�^��f/���x.��}�A��QX4-5���5��6��r��2����7q�/ry���1��Ix������������8��u��--3VLU�c�ʐ(�Ԑ�R���E:���3��9*��C/L�
�HII��:��÷A8N����&t����u��﹩��tU~~a	�FsWsj�{Iqۼ�{��'�'X��d?����j2�L��9�����<r�g���2أ22s���A�O��WW1y��o�mD�ݵ�lEJ�ol�W����¸t���~ґcW+;i�<T���[�e��{y��E��סc�����#ѭ[D]:/����Oi�`ow��0k���1w�{��TBiYك\ӗW��[6�y�J��*CS Ϟ9�h�\����s� �uK>{���Ξ\�MDQ_zF� ��%d�}� 9r��1����mx��>o��g��s�ڒV��#����C�&Ә��x9"UB4'NG�5#�o������R2�1��f�L47�/������{�U2cߡ��+���9	ʚ�P��Ֆ%9~E�q�i;���ahb�@֟U�5��|�ŗp0�MC`oc�����-���8q��U�\Ѻfb�_�};[m�p-�y��J{�Ve7$ٷr劾˖-7�J���,v4Bl���f�zE47b����)R��6m�C1�j����+�0Z�`������VE�9�J��\C�u�խ�bތU.|۱�l�z{�P���
���Fm���ɸ�nG������ܕt�Ͼ�,��N�îDF%���x�>(߼@\���s�jW�ӹ��D�[
���5ޓ�/��3���v!1�����Z��H���i����|��W�Q����ر��:����tt�ď�M[������-.qX�j5�\�p��5�n<T@��KW�Ծ��>��R���;t��M4�8�o�E,�ھ�\\8gݺ^���ƿ�����F����C%�eAwKKL�G�6��)S�����؜)F��+1���ty�r_������e���cz�ʀм}�S4�yQ��"a暩���u(w��٩ϔ�l�{�ʝ��<]�p^����L�;�ѿLW|_�5e�c���K��C�o��fwv���=S��n������3@m���koTJp��K�f/d�!L"2+\W�p�ivho��,�At���}���!�������r(<2�nw1������)S0l�3���.>����{���ys窝��VJ2���Nͫ)�˝�O��z��	��!\ć�u�(�V]ҍ*ɭ��d%�ZSW2k�#��\7hf��s��g)�0�s�<v$j	��0�QS/Z�˗�}�J���!�u��o�IN����֘A������S"�e�e`G��e����?��s��y�c�꾑��o#%��Ɏs?E*۬K�9'�v��U��9�es���ՕhF<���?��Wν��q    IEND�B`�PK
     B"BY�U���? �? /   images/05596fff-4f8f-4556-8b1d-73ff55b6eaa8.png�PNG

   IHDR  e  s   ���   	pHYs  �  ��+  ��IDATx��i�m�u��>��[��=�ٜ)� �"��h� ��8	0� ����`8@Dȏ��D� �A����8q$�(�EQEJ"�j�j��f���o��{�9{gk��>��CU�z﬇z��sϰ�o��ƒz
��Zz�t�#�N_�T�=�i8*U3s[=�s���on�|�]5���u�?�<?#�W�{]����n��������ѻ�}�����^?�8�������o����}�?o�=�7�ghH�i�|4�7��>�k*ߺ�ߺgܹ�Nۿ�"����0�Ø�Ӽ��xN����$�7���56��3���o?g�]������O_E����1�-�eYV��l���;���p�O�3Gw�5�񶚾�������Cʿ�W�}���=7��_:WO����T�i2(�%ń|hf毄Q��i����cJ�Ǭ2����.����	jx�e���L<zJ����˧��(����}�p&�!�j�z���\�j�1vC��[[eͿx_s9�y�� {}��"��7<���a��*�9<[�WX��5SdeCCD|ZА6q��Y�aLa¹P��e��k-��t).7�<�����X=�VK�s���(��)�Cߥ��k�����Ũ]
�4��5�]��w2��4�3�U�-�q����K��׵�ֺ�iO/�3^��a$�&,�7��΍�M��*�ea�'G×�s��'?�o}䙗�!�����o������O��7>��?��O��o��&�l`�n���,�-B�{$��[�ʕ�R`�s����ӱT�䜋�Uf�=��\�<e����q=ض��e]'P�U�KK�G~(�B89ϫRF�� ���6AMR�����Z�-��Iy����E�h��w����~~�>���.;���g⪝=���foe�~�����.�.�D.�K�������U�\���Q��{���������������w�D=4����Q��/~���s_z�}�Szƍ�<cn�>�&yఌ-d��X�@�r ��[��v� *�$0�:	Qg��u��p,6֟�1'0_6�Lp���s�W�q���|6ܸ���z*�o��e+`d�eo�LoE�t��jAІ�n�C����<&��p�m��e�Y(�P.��ش�@a�I��7�gwf��4�f^Y��tqm~_���.���>6N��+x��)�I��'~P�-�`~Ƹ��go�}����~�'���w����kz�[t��ڃ�?���?������_����dt|k�NF4�����:>a��"�����A`�f��`�~GW�m8��"`@���F\�������«LB�/�J�#�_�4�x
 ��G�|�|мcxk芆��yL.�gP�`-���Q�|1���J�E�(���r�l���Z}�:�l�s�Y������V��O�Z�y�?s������QB�{�$vHTk�]��%��ӎ�2.���>;e����|09yvp�Ƴ�<;��_��[�����o��/��w�ӵ�����_�G��W��Ԏ��G���%�WD���Qy<���p	,gNҁk��5�xrY���qT�.�n@#��P��ֽ18��vQ�2�ΓY�����xxb �au����,�ݲ��������8	+H-�ËiW�Â��p}XJ.�n�:GT���:4_[�n�A���HL�tE%�R��s�݆c��s| -� �R����/"|���㚿��F��8��9���!��sU�7��8N�Em2�00��>& t�)`4����1�'O����������?��o�������k}۷�ҵ���������_�{S���xB����q7oޤ0����4C��UӉW�-��2u,[$ڍ[�*�$+���S��+��0Jk���m�Z(�RD�6�GP�_"��cU0 p'6g��6��nȕPK9ò[p�ex^�]�dJ�����(]9goc_�S�8��d���iʏ>.R�<.���0�Gh@�0�I3��Jlv������G�ԥ~��F󤯪�[��0�m���`6�*S�ֺ3��$�����koE�o���7�{�rt���0�I�[�����	vkG��8��N���w'��~��/����������^�kF����^�[_x�������G7牉�g�������L9�7n�4 �sS��`m�0H��u�ՙ32�y[u������&�tvz�\��q(��W����S�;��
B^�<H��hV����1�ܾ��#�n��0� ,֐X'�/'�ą�'��
y'�'�{���=�o��yA�%0a1@T��!�LY�9������Q֍����U�VC�kʞ�,�j���
���l�u��O�"���el?��(�uI�7�sr넎n��q~ӛ����W5~}�	�v7R"���;8֙���6O���`8�܇Eh��x<�� �[O�;����K�������/��5�k�������?��T�c,��q���[��$�[����7):�^ �1ѱ�5�̨�=��p|l���W���x�%\&(D�Q��뀳�=�U��b0Ӊ�{w��hd���Mx�@�NO��W8�h��=��,x%`ٸa��4p����`�m�fp�T�#I?תdkۑ�%����+E��Ix6����.[��:c�9-bQ�#%��h��"��x|N?x�F>���l��,/s�V�ާ��J%p	��SOo�q�a�!�������r7]�x&��Jo3��I���z}���-�@$��u�ˊu�0V�V~�������?y����/��ɻtM�Z��?��?�{_���0�znR�m���8L�f�c|�lͫ(��Q�̿�͖
.��q4,�4�=�Zm��3Om늖"��i��[�c�[]�����_��C^( -f|�r5�n �`���ƶ՗
Z�(�sӘ̑�g�5�������Q!��I���2k�2��ʱwT�%�\��((���9 js���*]�F�<�ʸdjy+��x�k,��1�^��)]�8F%�j�72�;����/�a1���P�Nl�-��̟�ꗿ��3��Eׄ�(?����?~�Oأ'Bg�����v�kݓ~��H�X��X0�A���v�!-ñLB �ڃ#�$����ȵyeۀs�>�+�HVʁ�bP �2���V�������n^�!1����`�~�Rܸr9��L���e���@<�%d��$2��ل�n�]E���c�=[P֎�&j�aՎ@Z���.�8V�"��5]��8��kkR���kY0��؄�@Wli�]x���"4]M����������QK��˛(�%�wvT�q�?�q�D�!X?`Fm6z�=�������>��s��<]�6��������ӕ7C���h�� � qSto̶�&r
&�����Qv,3+AD:����ŭ�OGJ�� �$�T��YOH��g���\��j�.�\�ԇ����D�ݶ���JH�/si�2�$R�em^� "������B.9�m��-�U�ˀiDQ�2W�g��@��EMX|���Z�0��YIw>9$_�x&��|M���|Y��c>�Mrd�b�[2�����z��������]P��+g�����έ;���b� p�q\Һ,��*����@�o,-�U��ps��2��$}t�}S�dk�o�+��"�A�ilE,(ںf~ճ���w����eۼ	8 ��c�Q����]I�hY �P��L1�t�����H\)�˒��*�-�a���U�,#5�ə��3��F)�ה��~u�Ȕ��E��9��r�(/gC#��c?9+"k���s�M�n�t���a(�_�!���+�~1d��"Ȝ�doܦ�w�}���W���s�"8]P���������/��F�jhΫ	+�X�����Ml�s����" /�C&e2Y�!��%�%��d�)0AdXb�>��b�[��s�.�uM���Or�J[���\�*��;89H�Y͕>'M��s:_�F�]_c�ue���R_�ʫB�x�J��ߚ1���s&֕J
C���Ij��3�)����n�k4n���L�~}^\خr��9��+� ���n�� s(I�z����K�IM�IEe	����W��j��ҁӵ ��~���{�޳�ֳtvo�Q���p�n���g�/�5�.q�׎WQ�$��%�ƵX� '�9q��|A�B�7gM��+U�6�-9< �\c1�anFֹ5�w-�}�G��KV��T6�F�h��n��QRE챩�>�^��7ʁ�?�[���M�Y��R��n���2��?���X��q��G�9e~gG�Z�B��;��.�s�'^��R�g�hǲhg��E�P��MB�?�c����'z���֕A�x{��R�eRY�Ѓ������[���w��Z��+���jX�N��d[��lU��^����xܶ��pǚ���:�ʘ��u�{(���m�*Um�����3��	�@�Z +v�c8ĭ������R�:QJA��`���gD��"��b�oW��(�.���G�yb�<��RqQ{�w�� J����0h�����,h���N4�[��Gv�L,{���D�呴�e����()�������K; ?È��0b:�Va�w������cʻ�?���?������5�M<M�b$Ȧ�>#�&:Q����ޫ��E�uPnO��>�Ҷ �~P��w�6*��kW��g���^�4hY�:��"e�zӹ '����gh��#�u��@T��=�v�#qپ��/'׼����|��06)J9B6���l羙��g��}H�c�S޸�5�0I�6M�|&]!-ڥ6V'�_����5���ql�s�^=��+:�z�y�f�������_;�ǧD�ԮB⊋��:�ΧYm���E�``5�AT�E���v�w�{Oϵ���햞i�מ���9����7.�_p���2�2@���
��G�r+f�DS�e79�N�2�R2�S;�q�~{H�7*'��ݠZY�.;fW�x�>LN�~J�UU18 �����8\��dpmK�=Պl+.���<���L��M&fo�K�P�����8��M��y��KVj~�6�ۈ�h9�^�t ;G��ڽe"n=��0�l9�����,(����mD@�(hZM����eW�q�-���h��Iur�,��ns���z����-�&c�}�V,��G�u��d�)"��U�]��Y/%3D!��qq@����H),��qܭ��?��?a�t�t�\+, �ߪ����Q#m���8`߰e�4���$�錂�����%�N9Q-���&z��䆳\� ݭ��FN��Gۯ�Ϊ��zTrٶ)L��1��7�í��.�"i�?Je̍Ǐ_��=(oK�S�\z��"*�9/L��xt��mv���hbv�K[T����ꢩ��^Oj�g��Tt�ˢf׺��Ԥ�G�D��-)p8��t�t�<��<�}Z���8�D�����<��vsv�*���W͒sW��${�)x�F)�'�]4��C�}��c.���˨+�]���ݹs~�k�B��x\$�US?�d�Y��=��03���CnL����8ho����U�s�w�]NOc/<��#��Tq�c�h�v�Ϲ�I!��l�h?v9w=g�|Q7�p��K?��T����h?l6;�#��E��6O7�jS�=(�Dp��a�����B�"|M�#�|�+�HY�U�^K��	o��LPW���=En����|�<���^Q�k\`���%��d/2K+����[��؊�1��jѻ�d!�u�����$�R0�%�OX��L��ˣ1�]��Y���:�~�	Yn����e�S���HD����;�P�ߩ��&�)��aS_?��f,/x�8(�Ly�ʨ�墱���䚇Ly�C�5 s�S��tO稤��ěϤx9�j�<N:�bw��L�Gi4|�OuS�i�h�7�<>�!O�EM�9�4o~�˪G�Qh�<�5�%>'Y�p�q
�̨s4����g�KB٧~̂ßX�2g!���[_t	�R�����=�4eOD���}�N�ZD��&�B�W�jG��A(B"��j�qM�毛hC�I4!@����\DN޶�Mk��'^�0��%+���1s�ކTF��4yvo�ĴZl�C���R� M��asYٌ:yG�Uq���e��y�����z�����%�2�>�GH����rNRHj�;J�c��j���~����Q.��+vp�� �6f�v�'fR\���1"�p��X$J�d���P�q$<�r@��;ᙅ�9���5 �������8���ͱ�è�S$��#|�*(';�ֱ@��#Q�8g�wx���iZ�[?=<t����rCQ�mTABZ�~�]_�ѐ��!����\s.r�>�B��C2��x��)�-8� ʃᐆ�GTd*��ρ؝��,��Q�� Y��yL)������&�)��su!�;+��tS�u*�FI�3�v�<����W���ɴ�hq|��w/w���cU�3g�F�S�w�������8�s(/ۣE��L]P֭�NL�žzI�݁38�4�p��U�����n����]uM\��i�I~<���c*��ֽ��.�>��\��Y������g|>�J9�8�v�!�!���D�nh�э#Ŀ�kNڅd7"�"��'��{����ЙEBt�1��6�`k5��[�f=
ca03����y4���-_P�9�yD9b�y\�K��a"Ȫ�J�¬l�����rj���X:�)��O#p��� YD#����gmA��ʪ�V	aQݼ�\�`x�D]�\Br�.̭��ѺB?k݆$����{YtI����� �a}462P�j���|���+�J���BfC}�T��c�/�`m��Q't��6�|�l�c��Q���Yi�;0�TÒ'�Q �2�	�����i�C��Q�<�V��-��T��]u!V/
�x�x�NNN�w�*�]{���6&s0Kñ�Y>�`J��g��� ����vM�F�t�����GA'l�'��LL#5�f<4s�z����㝨�Z�At!�[ ��+u"��G��e-������盱��aa,�цﰿT�5L��Q7��� :��Q�����
l�QWmPL���c<�i�b�l\-��d�k]���%D����k�2GW�f|�$�M-�R~���u6���=E,ۺ��L��d��v�(H,f4���/8o�)��@�C����-�5���O�=@��KV�7�%}���{Nyg2���o�f)������56�UP��]L�e��=6A���E�"��]�;��堥��Mכ�?xP6�p[J���Mx��^��z��G�����7�����Ay)�����(=T��U庬����PʻRm�����Ae�+���L�=]3:xP�U�WIK�|{�멧�����7)TVO=���)Ӯ'<(����zڜ�]�B���J=��SO�S�!/"cz7���{ꩧ��7��Ay'��rO=����G��RʻP�)��SO�"Xq�{Ny7��s�=�������=(�BĄ驧�zZA��)�JE/S��Eƛɸ��-�)?�1�{ꩧ�0ԃ�.d#�,��c���[���ѥ�6bӠ��߿�;O[�w�0��n���q���w��L;���d���X�#����s�;�<E_� ��SO��u��:xP6=3��v��6�ϼe��[��n�Aw`+�ڭ�gL�D� ��<brFӞSލz瑞z�i_�=�����%��<���N���=��f�;XZ%��n�%�]��i�~��d���w"�zP�I@�����v'c{����⋍hs�.8+�_���3�nݣ�K����٬��]����;���b=wM�j�s�'&Ѝ2d�k���]��[J�A�i&�1Y1�y�b��;F��\��A��G������RS�ݏWMy?mzl?'�~g���tҋ/z�@���ع��|ye9�����DEYP�Z�^gj�ԸG� ��{ʽ�2<���
@W΅k"��=���x<��Tn��+*���Vp���s�Fˏ>��f1b��������Ёk����֦؞����ó�x���uC�M�S)ɢ��1G`-3v7؛s?QMe�0�<]�h�9�ӡP�ך,Փ���}`�������A��P�9�& z #�f�l�*�g��bPRQ,)Lxb�f�cvf�QV��P��& e����Sq��u���w�� �e�W�����.�R�\X�P~S�n�|E��j^$\�:�輣�U,�o}o^��ʡ����}ZτwT5�>���X4䩷������ᯞ�<==���w PiN��������b�.@�KãQ�ly�3�l���u�+w� ��;�IEg�����z�}�u�:>>��������9���XsL��΍�r��!�&U���Oǡ��x�a��2C�����SF�`�����Â��N�p�(t��+�z�P�-��7��ݻwi2�0��dP
�ⴝ��������A,��)� ����	?��6Pw���V$&�v�c��������k�a��t��*���w����qh�bOIFs� �}Ǣo:��"s���&g�,^b8�%)u�),4x[�r4}~L'�O����=�|��kL���(�~�N�=��`��[	i2�=�`ܞ� 
���LU̜ �1XB�Z�������ѐ� Z�m4����E@�l"��Mhz:��-Sy�Z+����l�B}
y@��p,N���e�M��+�NC�+�6�&�H��N�BS�zA���	mW��{�������E!�5&S:;�a� =��s�\�g�ל����a2�cG���$�V��:H�ibC���������sSW�|��&ʡkπ����|4��	d��}��E+cZV#��U��i�������ÿ�4��HD	;+.ղ%�/T�X�^�ܴf��8��s��Y!�)���~�]Qh�O�b�X4�6s�c�vC=�t�l��~)���)�ق"i:��D��p�-�B_��)�j�yEv��`��g��\˰�PC�"�(v��,��K�VN �(J�_���ebװ�5����BE�)��i�u+܀�C-h�]���e���J �P�z���C�1{d�`p�>C?A�7������t�t���)/'���%���I0� hS7m�-L�>1�k�.\�po0G��6�$k���e�9`�?�� �Lj���yyjBP��v��g���"_���£0�-�V����;�.���#��n9���0G4������ƅ��{�K���~�����~��ݹ#��ۅ�yhhX�2�]b�c90&渚���zjy�g�"I�Y��®�#x���&;���JѲ�|NSʺ26���ID�|p�V�"�Y�h#�`e�ku�zJ�">Q=�Q�4&HP_@cR4E��.}��k��X���9���E�k�j��!O���博�E��A�ѥ�9�&8xP�c_,'�2�˔C���R���#`Q� �#�N��"<�؋re�]{�3�S�����M� ���MAtZW��Ny�s�ϣ��L�%���eQ�V��h|m��A�zNy%�2�܄J��?o�<c�Y��Y��RW�b:���f�2��܇�ԃ�4�S^���5`��_��m")�|�r���kG�}��崯��<�:���K!��������sO-�s��J�7�[J�_�;�}]i2�}�6�-ҧ�S�~P<(S��ۘdo>�z@>|ʭpelcӋ,VS�bw:�<�p�}3�Jj�r�h��%�^�2�������EO�k�E��!r�m��!u�o������Z�~;��w!�s�=���������zꩧ�!�9h=���r/1멧��F��f��A���z�y�=��#ۃrO=��'��w:�9�]���v{z�I<���[P�|�)�F�_�E^�L��k�˂Xr�=��������v\^K�cϤ��Ds�j)����|�xʳ��߼�{q�։3lw�������!<�/(e��~�9�sFB�����Ϯm��Q�,qm�����؉���S�N���ي��itcDggg4����c+�@�YI�(���)��v�>>�m]L�T<���`D4��R�����e�^�8iif[�)�ʂ��#N;B�c�o�,��I�<�̱(K�B�a��Lu����c7�4�'�{�%�8�u%��Vp��a;�tdG��aN��4==#W9�'S�V��y���r8/ L
�%�dW�n���xȋͤ�r�P�3�ϔ�e�?ī�D����eC=(/"L�[wn�x8&3,i<K�.s�xe�L�5�P�0��1@6:[ r����X@�(L�c�l��̀��F�t��Y��4�y�n��ץ�z�x=��gų�#�$�����#}���Qx�1��~�q���8�샘w���͓���8�����IXP`�=ס�K�g@-��刊QX�F��@0r;V�̡y\����b'�~���G O ���0pb	P�|p�n�MG���	(���9����^��!��f�He�m9 f��;;���X��Ep� `Óc��" ���=���K��4 \7�[mA�����pf�;�Ue@�.d�A6�S1�E4F�He3�,�6t�lz���D�L��٥ˣ��4ߝ�5�iFvۉ�\�K��)rR!�4�ɮb�.����;���f�@m �	�<:>�:/(��g�&�/�!��k��'�Z���rUv��J��d?.�(>��=�C��F��fM�쐺Zzj�8�w��s��	�J� ���ɺ3)g@��x,=�)���E�D$a����Pu�@t3��_�W��{E�g%϶mX<�]����� ���^d��e'2�6��\~�y�x����E�C��r=�ϼ�@�3����V�G�DWb`8n�(��rv����#Nʽ��|J�c��r*SA����EY��lc��!��}���]�s���} �z��ˋ�Ϧ~6[�<�Ĩ�G ".��Yڸ��}yRn�Ĭ& c��lexa���G�w\}d_X���ڕ�u��w��`r���T뺥ܮ��4&��-e߄����[`SG{bq�Z$�K�eU����)Zy��̯ eM��=���,-r�j̠k�j����zaY�|MA; #�޺������+�,�/����L�*C�>W�>������A��մ(?[�HZ�%Y�=j\^�'�$����q� ���oP.�z7���L��5��XT~%��,�}�\�6�~�{>3��1�eʚ�֤�sM���G9�-��������濣�\?T+qZ���������t�l��|?�"9��U�~�S�L@�_��(�'" '  
AjrU����*����&���/��y�\:�LF�+�vS,��0�U�N6���.U^j�^������]/�U�z?b�����}�8� (��f��׼s�/똝]Gbn����2���e�;���K��5��q��re���y��t����)�;<��י�|:PF��^�,���q���_�����ȣ����uH�=8xPn�h�t����
y,��y�a���{ڎJ�+�v#G�i!5���<���]�<o����<��0�ao��尗���9��w!8�QO=���#Bx�z��e$�,7��hq�f��_#�-�MF;�]9���w��z�ך2��to7Nv]�GW,����ɩ�.{닝���֤�X���ߚ	͏�,!;�G88�g�Wf�?w���=]=����������`��!`�����s�J�ؽ���` R}�h[U��9=r$7�st�TM|�h}�������Z�-�|]h�27�E׹qSo���-�C-:�n�	<�-�vc�}/V��b:xP.�t/ �O&�6�q	m���Uuл�K&��Q&衍�C+OOO���ʈ8�Nh4f�,�A9,�x��A������pd�)B9�[��������SO=-"��F�2����.�����^y�m᧯ҁR�����nއ;[�KІ��1��a+vք�F��r]��|���óq4�l��|<�} W?��p���ը,��3x}p��ӿ�;��{��T!pX��N�4 ]�e/WG�T_��<x ��%J�8S|��/�����o�w<=����a'^+&�*F1�ƀ}�������r�;��G�sxf�N�5��ǜe����y0w�e�_��_���b\T��`��s.��E=kK	:	<0�LC�'��������o>���{3UvD�xC�y ����䰧�z�L� 5�~��Ti4��(��}��3������/���?6�}! ��q\^��XO#���y�{��f]�]�Ӌ���-��3��	k�h��T�Cd�=�,"�sJ;R�%�$����SO�:u�4�3�d,��J���X�3��|��;���|}FA��S�������
򽊰S@ci6����Ӛ���h�"930�+��ə��;a��SOYޑ�q�������4�N%ӻ-#��n���^]�g �eT��dȐ^��ۚ�cI�n9��5���h<�r�G$���޽FO==ڴX� �y$�,�0zP �ǧTFW�)/%����_�C�#],**?!_��������4	����n�i!�j����SOKIv��%F.����<�L&t2�n�o�Jm�8��I�b��w�ʪ�zZN�ݞb��P�Ls��_K���|�ܧ�Rۆ���=�t��+V\,�`㟿V���:�\����>���l�k�<k=�����!���ƈ�(�lV��_.�胄�F�&��e�=0y�r�37�|_2���pE�Iw����ZY��'~�i�oȞ~b9r+��%8φ�=\0V*s��!�2Pa1���L������2��|5�|�ZR_t�ȗ!Wγ"���OE�Y>X�ṍ�|1��M�]�JkG��M6Y	ar��y��̇�=[��mU?i�\��ȶ�k�#P�ts�����"�K�}��6�����T�>]o��_q�hy��=��;9[�i9 �1�:�֙�ϙ�1s��0J�>=���?�{�#��(��t������t���,�R���r4�e��S�1�v�Dݼ��s�ٸ�r+�4#d��V�a������k;�*=Z@�g�/���؞EJ��r���W1�*+�	��xX�-�C9�d�x��J>��i��|���A�D]/��G|�p�/���{q�ա�
��̘]�{o�w�,cWے�bSr?y81�6��Z�0�T��y�Oߧc��|�Gl����X��`�"��O���n�"����p�r|F�zJ�0���E�p�e��Y����m@]o偎G��`����\B��c�<��Eo��Y���>t��&+r�lU��@$3�sG�Рu墈����U+��j��1�Br:��!���@����)M�Ω>�0���&�_�xS�k�i�|P�(�4:9�፣�P����S�~���D ���U5Ua���q��ɔ�PG�B��c��i�E��ⲍ>�bPҭ�n͊y��r�-���X�
�(xw�31>�����ܸ� 9i_P~����w=�"�g�AAG7����,�{"i)�eN�`�B��{����S�6.�ҧ+w*;�� ��)��"���2�]���d�a^�N��MiW��E(�����ի��Ruo����n{�\�+3�OX�m��ѐ���|Ĉ��(v� ��:L��1���� �H3v-�Ş�(g��߻}���ă��# 2Ħ�0��,w�1��n�*�,�.a��d���N�G�"��'^�. Ou(ZtG�ߝ�9jX1,�8foR�³�e���W7`]Ó,,���T���Uƙ1h���w_��ޘV�~���G��e�S��j��Ghc�ޡ��l���y�����a>b�D�"r#8v�[��,��.;qd��'e|OU�����Fbā��,sn/f��E)ѯ�S6+�[c����?��<�A�`�����;E���`Τ��>9�"1ʃٻ���ar���`6��0� ��a)屛���Z�/�	�����'4���QE�h ��wצ�Q܊8f D�Yd�K�F��,��Ky-9�hK�������S*�Ja}1I��i?�;� t.8J ��ı8`��]t�y���e)b�����~XȪ	���%q��b0�C@�������iZK��W#1kX� 7/}����[������B�y�6,R�.S���e�^�Eӕ�rR�̩����<)|8�S%�f��G�&��O*I�ʏ�4��1(�x��q_[(�*|�T�C�i���ܦ~>�nt۝��,�4�s�(ϋ�!�P���9���X&�=|���[1 +��ܗ#|��Y�_N.�Js+���|"����[���V�W�x��$,�>�Xi� V���i���ń�@4En<��^�
��]b�����b��+����q�sv�7�1ʸsb$�z�b��qh��.�]�ܦt&�W�-�f%Kip����	ٚ����-�d�hk&=��;�����K�4�B�KdZ��v�w^9)�Ž��#����M�f�m3���i_Wc��ŉ���M9����
�X��pN���Q/���:�A���o�rPI�\/;�$�����D!�y.?��+e���>H(� [-�*�Z������8�w6�0�����S�]�I��+��}9|�s��7�)DmtN��9�$�-�x�W
]9��1 @_	�lPj���5��8
�}L*	m �0��
�uj*"GX�� ɖ1��|��4Qp�>���)�(k'\�B��ɁXN����s�������aA�>�1�u�#9�}юl��ER ��*�u�
�/E!4M�n��@���<yr�El��b�ix{���+],5�&�C峼c,Vu��{����e9�z1�nE���ƅҋ�f��@�W��qرs6"Z��}">2�O��*�ס�r�:HPVގ92E^��z1SI.�l���;�l1~�(�� +^��@�A9�L�\f?}Qy6�X��a�|���;u������ᆚs�u����]�����EX,;�c&	 ��������l��g ��R[�ʴ����m�ȗ�y^�њb�\�����'tG���v�v7 i�F`}���۴P�llO=g��I-�s^|G�Wъ�²�+2)ޱl�i?�_m ����0 �EӼ�Y��N�:N�-xr:�JIJ�|b��l�јj�˱�@�X�'�0�Z�<#�GѱO � �b�����G�������Lt�yU�-��"V�b %f���۲y�s��F�J8�E��5+�����Dv��~��0��ie5T9Y�;���y�r]sZv�P���ae�r�A��K��Zʲ�lʤ���l��q�p.��v�B6'9�f,;�AGQ��;;a�c!瘻v�J�i�����;G��SZTM����`P��@#���p����!�%8HN9'�)��2��!����sZ������	�D2u�bf���ʝ�]�p��{�o��E]��t�xP���(����%۬���v衇��69�O���b]�zPNmkn�Z07t+g��� ��w�MA�v�Mk
�s�]wlM�˛9�z�+��ЬɆ�v������lƮK��W�����-�g��b?^2y��ڨ�>>{Ƀ=�\�84���fq��W�+fW]�U{�.�v����~��/�����.2�u̥ ���o�b)�l��K�i�%��D�\!i�5ݓ�AER��E����/I������A�0�N�f�0�bg�E�{�H]�i�J�]o3��_eg*���] p���좆���u�CNA4c(��ü{T�E�r犌������~;�y�l�+I��2H�(F�#((�;Pb#�ڙ��t5;?�d��1��2؝_R��9*���h�VP�0�ʡ^vj� ��H��tI[<CǑ݇���k������NrAxC��)���L��` a:PP^L�t9��y/sV���Ń��d�QC�1�i:G9�b��f���ז:�}�]�`����8U\J�^ǦY����X�{����k���ʹX;��\M���enǱ����[��EZ���u��2�l�}hw�K�|�� AY�e�k7��B.m#23bQa�A���M�(�]�����縹���4�θ�+s�cl�\R���~F��������v;{��4#z�mg��T���U����x_�YEy�ׅ%��ۢ�yܔ�0������M���_Zr��V+u��#5q�П�{.w�V{Gii�5=s9FA>3]0��*ig��sϡ���uį+�p�8�͋Q&+G�aS$WpGTs:e-e~M���&�G�+�:pÓzB��Z�A����E0�'��:��b�C@"J�+D|�v��g��w�ಘԳ��)ĥ����s�ou��.��ٵ;34�an��,v,ׯ&lO�`=c~p���=�r��&�_�袃8wq&iDRF�i�	��|�u�
�r/^�#���S�57�\u��m�g]�/�w���m�%,����d����1]����	��]��vزE?e�Ar��v��<8��S��@�e)��_�ʬ^Tu��`�M� Kr�1}2�%��3�xJ�k��.�ţy�P<�m�"&X�c� �Vm��u(�J�{�-W���Ƙ*�w�k��g����x�6�}G��1�`�Qu�Ix.����8��spuvL�%d7�4>m�cN6:���&HK3@�N@���Qn�f%����Մ��ڭ	(�����`@97��X�0��hk��Lm��3�!�J)�3��8�s�̓��\�l<{����*/5�M�M+����]�9���S��p�'�a�`Wz9��=���Y�"������DҎ$fea�.��p�Ǌ����!K��&����^^1���XtM��4�Mi�N}�~��,nI�C�6k<W�a�ҹ�N�F�$��1=�o~c1�a�u-:P^���4�嵗Gy�/]��I9��&� �gi�=/���uεk�R"(Q�ssx��p�ېƳ�m�q����c�u�'����m��£*7���~��6Y�xC���dK�0����E%���ZF�d�"�pQBS^Ȯ%�~M�Pw�4�fA>_���'�yq9� �L�
i,[;�Ȩ��9���6G�텱݉�����+ٔ�gC�W��^�IZN��k^ %��e���;	Q6q˶��i�d�[X吅a�d�>�f��q���^U�mw�$)�o��pd��0f+Ya��1yG�Ѽ����˰c�!�,d��7Տ(�R܎D�l�G�^K�,�<$�盧�ufc��Z�hE�f=`۞SV@�
�&�Ujʥ���6�r~�
p>P���r�d/�ݟ��k�{������i��P�r�����%�� @G�-�1s�f�g�
z�Aib��zG��H���N50=���wUa◉{6�X��e�*�0�͜�^��d�w��'������lH�A��_����A�����~l�R\���hn���ՙ ?~���͆�3à}�Qkׇ6��i���T��݀VQ�J�dtw�E��䫦+eQ&�ѹ�r�Z�Zwj{ �]�&˾�e]��P�+q �a���M\��a@6h[�6c��S��߄1eP� ���7�p��u:��Č�p�0�u��>�2AKhF�:��9Y�Ȃv��]7�3G�_scP%��V8U�w�%�ȸ�E���Ƕs�֬��h?���]U%�EΤh~*�������	?��Ź aiڎC�&�u~���g~l�|�ܗ��@��� b ����N�͙w��
����P�6����okEO���YSB�}�Q��j%E
�F�+}.�+圚!eS�m,Q#��r��o��nǵu��]�.�����bb�ns�N�E�(�i i��<�[S�+����s�< �ax�`T�эO�iL˴��.�&�0���C��!���B5��E�8�dZ�$r�]��̒����#����UcR��n �!��1=@؁��0]gVy1���&IeV�������HV����o-T�>8Â
7��H�� W|�un�g���wlqģj��#o,ڠ�@�""��f"�_���"��c�Y��
��pP�j��Yc˦�Yq�W)e��dAGc`Y$��Қӵd[�b���G�ip��F�����*Zv7�c�[N�j����`�-�1�4��. vEw��hHb�=Qy<��n��#��.�q5��dx���y���ܾ͞%}f��1�(m�^�i9z���zO|/�W��c��-�b�z�=e�KiQ?6���L�	އIG��Ic��%UI�ˊ��)�B?��8D՝�)�v11" >#�2�u��mz���5�[������/��P�I^����8F�{�I�
L������*������<���s�q���c�9���c��%����׶�r[�ᅃ�\�����qʲ���cz���ozU����[��	f,=�$&mE�a@�*4��V��뮀ۮذ-�C1!F�C>`@n�\�3��χ��9����vP��ʵ��d�Ut�@2X��b�٫)�~���!G�cl�R����LLo�e#�@SS�tu���G;g����Y%|/�x�E��D����])�E䋈Kn��A�vMפ���XV�r&u���$e	�x�)����t�K)���ߢߑ��h�b����"��
���k��K`���̛�LO����EM��M�g�H������/����S���S}Mi[�2��v]8(�l���;�޽{��;���ޠ7�F���>@oy�[������m��cz�ޢ�O>��c�%�
��
����`Wlp��cYn%�<Sd)r.��P8�R��
 � �3)�QNj]р�[
�ø�����9�E�b6��k3�h:ƛd/Y�(L�4[j�v�Q�Dnxag��L˰Q˴�Q��#�d��
rߡ�d�م�X�"-�"�C_�S�9�N���6t���d�E���xX<��$Tj|$��e�7���B�V����]�<{⧜H���*��c�n���{=f���awy�������o����=��w���|����w�`�""��+�������R@��o���o޼I�a��?pĿ�s�����u��4���\��8�鄦Y�G����!��[�m��(��F�A�̪��}?+�bbN���ƒ  �;�W�*˚,?O;��/��5���v�Qi}�I8g|N��Tġ9�(��>��@k1sPqGl%�}��<.^����~������Y'���b���cFC(�`^��m���_��x�9��;�t�_�����Α��PA����,�f0%�5��F�,(����t;�X�H��������w����1����կ~����$�8��ޮ�t�*�y�'��X��z�)��G?Jo����X�ۥ�P�uXոR�E�Q-r������/�T�����6.�~eT�������W�о���qI�#:��}�&�8��,BpI��J5�"��V�%7���|�xiF��bP�$A��L8���+<:��)g�����([��pV��(�=�����;�z�{��=�uV��M#�[�r��^�*׺�p��}�J��\�Z:�V�a{�3��l5THJ�9�ⰃΠd��4`Ɠ��(J���_��e揯��	p� ����������������/�K/����?�`�Ѷ��e5�{�.W�~��}a����󖠚D��k�2�H:xlX�`D	T��[���E� �N''�Ymr�,�D�+M�4���*�z�W  G��2��@IѴ�Ү1�c����S��ɵ��FM܆�h���F��;mi_m���/&�e�]G�e��r��U���3�y���%ݺ���"�&xq>žۇ7�2`��.Z�Z��*)��'�"�xҎm�%�Z������p�bYt7�� �,�8[�8�Ŋ>U�iΩ��� ���o�?��?�/}�K,����N�L�XM�!c;�?�\14����ցAB��%�T-V��<��@��k��=�v)Ή4����P�	�y t1*?��2�ѵ�$�I�������i�����F���\��]��E��'�GZ�$�H�k��1h��E����E�ɢ�4�ס�]���Í���&v�YCѷ�U�JQ� �6'^kl�e�[����m��fM��B�$J�΢6/0WZ��]9���oE'jv��S���s�y(�`�N��p��^"�Rf�~� ����iz�;�I_����_�2ݺu�U�}0*�b�QŇ>�!�!���BE1���U�4�MYqV3w��,;�b�RGNpxR4^_�L ���:�ّXΪ�ӆ��m���.��Q�[ir�;}{:w�ڛ8�((3�ˣ�h`J�d䀻�z�4�o��n�>,'}Q�]��<��2�LW�����Y�]G~ܖ�����(����^�i�ſ+������>�X�:�S���,�9쓧�I �)w�@�it4 s*v�pPRN����� �L$����	������;��.ƛ�JP^%���Z)T J<�k��F��˿L���'��j*qD��FpZ���0��1MB�'4�}���`=����a�����%t�K�1�֝�w�Y-E)�᱅|^&��6x�CR� �� s�L����+e�=I4�L���v�p�}��K�^0�L�7�˫"�%�ZSfQ��-O���ۄ��V�sʰ�L�ޡ��*���.H�oߺ�C�7�WGi�v[�	��-�Xt�6�;��ZN���xrؔ G�A�2�ᠠ��M7�Ӱ��ك{	��Cj����v��;�v�����G>��O~�Ұ����2���Z���/GauУ�(
�+��+��~�eۇ�ue�y� ħ��b`����t'�@O<�*��n�����$��$��6k�]���vȦG�[R�� r�����X������ :��5�Xc�9�0D��
O�2V��]累����X1��������+��	�<x�0
 |����ԊJ@�����Xc���*ڔV��:� 0
�©2����c��q �и��.\� ݾs�����}�ʧ��^-���DϿrF��h[�
���A{z�2��z�:R�d�n����4��3���w�����=��{�˸�������o���?O��ַ`!7�o�	c��9x.��G�G�>���2�g �n�Ɲe��� `(8��c���:�����
�!�y�����n?v�BCX����8����<i5v�(��SO�(��
�8Wq!��%�~T���3ϰe�[���M�2fs X���T�l<� 0����?-�On�=�Π�{� h�����ٛVu���Xa`��c{�#�i�`�~挢�,�7io��˔65]V���z�����Mkv��܎Q,Q ��T��˖�Iozӛ�mo{}�s������x�.����`̀��?���-o�{�����A���ǙcV��V�G��Ice�E@�M�<+Bx/J5�B��SVY��E�ճ����d���zꩧ���^,[4�鰄���M��S�������X޹s���O��O��z 8Dp>�=�=�˥�l���Mi'Pε�(�����p� D������a���rz��� 1ly�|�#_M�v�
�P�_GUQO=�t,R[f�=p���D1���o��"@��������g�O}�S2BG4��g��n8��p%hkPւ�2�~���}:7	Q_r��@�q��?�����p]����su�P��F ZL� �����z:<�8"Q�d�5��xr�p�GQ�� ;,-p�B�f���} oH���v��JP�r����}`� �(o�r��`�ʩi��<�'�'���P�ԃ�f6���2X`D�H�y�������z��L;�?�B��cQ�5^���4����C
��5�*��� ���A\�[�i`�z�c*�rQqA�]�8��]�b����
��I�E�TME��,6Q��e��f�{ꩧ��I�u�<�{ep�`JU���e�	�}���gI���0���Ck�/��#/(��! G!UƢ�L��`�D+��X�]�3'$�d���z�|���U���� �?���k�����n��?�3�!�U�mżE�׵@Y�v�|�!�x��'��B}�b@����&��M[��8�y��SO=�tєK�k�eFX��|�;�p�I<'q=�A�k}F�y�e�JP�_���d) e<\�A���j�?<@��*�Ṯ.͇�5�=��SO[�2�*rU`M��3��_#�DߥH	 M��	�k+���.�/Ċ�w�l Y���ӄ��ZlEJ��IT��k�.���� ]�Xñܰ���93o�dC���pԕ<䴖��� h��dͭRJ况�0�r�<rW��OQ�zꩧ���T��y�uL)p���)�)0�;�er�EL����Ԫ=�����
�\5V��k��<=���(��1��"X�1����Q���詧�i�^����H�G�Y:t����u9\:����^����9`�ju���e�۹�܍'�l�:�@q��)�x�WC��{o��q���Usjr#|r��Vb�:�V.�m<wU���r>�YGb��n���ݛ�7��nqy�����;������f<��M��w��ڡ?�d��{_+Iw-�S��&���kr�2�*�7��ʼ��7@����|�?k@#�vi-;�\8��q��"��G��.��̧.�Q�Fٗ4r��ɍ�SO=]<�Gm�N��;s��ZB`��x*I�����JȖջ9f4�ֶSVR�7��ʑ�����s?��)�$4M�y])���������um����rr+�4;��w�P0!�ڭ������/I3�6|\7���WH�L��F�V��<�gZ��$���oU��(ԫOI�˰SV3�<u�V2e��t/����r䜝� �}S{ EY�?��SO=�t�ś.�D0��i&�yݝt�)k�����W������E���M��$��첵�&�<X�dw����t���k���^�n�Vq��Һ}<[�fEy��do���l�5��2��4	�8Q��hpԴ��e��(�e#�R0�P
��O��9#��p^%��f-P��+Ì�DvVU�m�<p������G%�f���0��g�$\�`��7��)8S5��}6ʗsR��+�P����)�v-5T���^Dk���b�<~h7�mʫ�>6�y+;�{��%9�FN�-Q�ED�E'������_���]Ʀ]��d���)�~߿���˝��-���W⋜Y�c�uk�lVq�v���pƴ��o�C���6��9��ppw�1�f�]I���][f��Z�w����vY���Mݮ��@]��Edֺ",
H���u��|'&v�s���
�+��t���a����󤴝#Slgm�]���)�'ڼ���\�����i��ߝ��ʾ�&��b�:`�`(���6ڷ�H�{j]��5+�{��U�`�(��r�j��s9�FFҌ�U�]�sj:n=7�&t^،X|�M��ǲ�U��l%[u5]r,L�X�F��G��
�a�hdul�����ף|HV�f��'�o?����m^okL\�(=��>��ӕ�p�<.b\�]�}��a�Y���h6$W̔^���o4�_1Kt�+�u�1������4WX�V}m�ϫ���\Z�-:}�pG���$0/+��Q�w�6��e`7#�G�-�f ����l�]�G�{p�>��*'l���{�1�z~�g�PX�e�it|D�7OB���~4*��1���I3�Jy�!`�a��˽��t���ѵ8��,"Z�<6�:�p���y�����,08\�A�=�s������Ҏ����by��ㄊ�`;�d�a�y[R'�ɋ�,Ms�ΐ]�|�n*���Nw�&o@Gx���aN Vj��Ϫص��LZ>^��q���]5�ƒ�6]�9�hVl�e����IK#&�h8��rQ����̓cNp�d�ІS�R�8礷�2Ϝ��`�T�W׼�6�����L>� P���4~L���7��s��N8�0A۲tg�hJ
�ضaec��9 чE+\��O��M�e_�ˈ�0��x��z�N��n0"�+��J90���TnY�����(G�uFW�I\��
aF��(�Z>(��h���
��p@���J����ˑ.�Pkp|�I�\у�<y�Z�I�����찙��D�� ^ 0,:%� N�W�(��O��|v�s9R`��q�9���S���D�e�qW`儞_Z��!s-��h���Hc�N\Sǜ�.8�-g(V-Ҧ𵃒���(�A{��IL��
�2w�Sǉ���yPp?�a|��O�>='W�i���E_$1��6Ď�1c�x<�sv�#�Kܠ�ɸ&�1�B�ٜ�R��*�T��ߺɤ��v�������wn��+
��HX�-k�������0B��)�I��h'ZS���Ƽ����ʹ��* h�w���S�3�D�+N�ޣ��3�*�DL�c��r��%��cD�D���(L��t#l���f�d�GՂq�7Q�0� ��ݻa��H�i��o����P��ѝs��e�S.���PX�M��;��٘�L�R�r;ig�S(�
0��Oxk��%3�+��@���Y�؆U��"�h��>��Q�pŎ�B�X��#gy�Y�V�l�2{ d� 5����}�������dkE_�a�lC-2�9+���/}h�E4�Y�*�e�A���z��b̌-i].�k�`F"B�(�
�d�czĠ̫�L�V�����Xa+	��e�?d���Ǧ#fЯi�l�8�B 
����0�)l�n`?���,����7y6��ĸ�����]��q1q��Nb*[��; ��ݔ��^�2D�+:,:u�͌CUg��x�*'�!c�i ��������qح�CI��gt�}oʛAnm����[.�=3�x�r��G,��Q�����c��C��E�'�}�au�ۏI��x�rd�Ea���S^���<�L����̒ÉD�n�+5
����x���P��b�N��Ш�
rf��z�Ւ�� _�8��,tx�X���vpx���M�R
n+S���3-&L%�)2�����2���P��-�]������'=d�����3Q�. +�*	�J�p������(�-	��S�&�!?��b�u0=!3t-G*צ�e�D�*�x�Z{^�JS�{�ꯖ)��Q/;���L�(zY��
�m��Ke�^� pS� ��<^r�l���� �"")ׇ���P��8�QR�ƪ!�J�C}饗�\=W�iڼ.�������"! ^M��\e&8��+���/�LO=�TbỆ�뽗�]�lU�l˒|�_�L�7i�T|,Nb���,�ճ�&�.':���t5�����Iw�l㚈}�&Ee dQhr����������u���寮��N>�x�!c��e}�]����2o�%�|�s��6��r�JG�:r�2nB��~��]�2~�/�j'� �D����,h<�\x��懳˸fjϏy�E�w��Q��Cw">����q#�?�1�r�����-�H%�X³��_�Kr���ڠ��Tcux�ט%��7?(�V{=������͑Y]� ���௬��,�o2f��tŌ{=2'��S��([#�f@ѫ(���AZ��K� /R�h�'�x|�hU���,o�·��hŉ��+X>W��U,5�v����|4�rQަ��4��`���'r�E�����Bay�K伵�Xہ��{4���Lʂ��f��vۭ�ig�/�ف�\5H���z�U�/�ѵ���,/=�g���*�wn��I��4?
A�h`������3Q�kD�؏�	������OձN��^p�y�k-�J�y��Us����+"(� �Jc,cu@��w��]Q._9rA79q�K�N�]GT�	G�6���Ҹ��-���	a�1Jy�Ŷ�UB]OE�&M-�@lE3-<ם����@�Sёv2o�ٖ۰��i�$�d�6�k{p~��φ�̰ʈ����K	�I�F��@-�ռH�/�)��.�2L�-��J MT�r���
2����q����ّ�kۚ8�`��܂)�ܻ&����Ƨ.�-��ҝN����M�j������K縼3�sю]v#>�H�7h?�4���?3����ωm���l��������EP��pk�cŃ�/����}-e`��
�� m�rn(���ݥ���)�r$F�9�(^�����o�7��M���>�4c�5 ti���v�7'����P#��U�v��t%�"��&�d�D;c�ƔL�:�׽�}7���LN��+6O�՘���E���"�K~�v��8?�@f���|j;1�ߺ^�
�͹�ճ�X���-�QV�1�k����W;c��V��z-߾�o0������<�5p��V=Ҭ&]Z�$.7}SPF� W�,9��H> 1LCp=^����_��(p�H����_��-n�D�0QW��ZL� ��k�}��7=�J�8W}ۢd�T(�>�v�)[Rfq���~�1ؗ[��D b��|�;���{��'UZ�y$J+�ЅXCE�V;1,3 ܟ�����c`VZT(Ok�7�6� �0P� ��$늞z�G@�G��̵�>�xCC��@��/�w�.�_�3D��U� bO�m}]��Z`��?�� f�G}!���?�#N��TYu�eo��]�,QO��y@7�/��Rf_�iy92������U��G<"�?��?M�f0�`L��>`,�`}���|Y�r9Fvi-���x�r̐� a ҡ ����,�*^��/~���w�s��QIA�δ���e��K��}9s�p�K����W_M~��t�I� 8���Zm��/��k��3�oP���k�r�u�w]A���7�g�B��L�����;����,�%���`��^�h������#��g���p��o/���o1�
��b&H�u��<� �2���v/�K^x�Qܹs�W��q���y2
�������?���T������g�9=][��5=�4K�+�������O��b	�C��.D����Vb�'��vk�En��h��q/��"�X>�O$.Y5��K�7�������/��/H���W�Q�5f�s���e\��v�q�<������g'����:�����:�vyu�'\�|����}W˓�S�}�#y��y�.�cl��m �㏯$�Gs6��[k����S6i�|��g.K���r5�S-�r[d% )KY@*�b[�z�XeǰH��R�9�͗K��u�T%mx�_�BR�"(�rɸ�f"��[�E�����{?Yx�Jv����Vp�-c�xj4�6�U��?s�Wo}�<9�ʪ�jb�7YsN,���ģ;��1oV}��j��=[�(&ΐO�tu9ʿ�W�r���p�1����.��(|Qtl��h�)�U��mh/���0�~�w~�e�P���GAQh�6H�̧>�)z�;ߥ������w�3���,�c��y�+���&	:"�+c���uWb˔N։���Z1)��Dow$��� ���ޞ j��m
_�M&��bp��q��c�)�|��Ԕ�\� @� `�8gN�L;~%���PB��=�
�G���|�:(� �ީٰz�nB;�������Կ�ۿM��K��rc�Ayzm*Ǖ��7�]�y/}������M��u�q#�HX<�������_9W�}��~Y��[0��ϼZMl_��C��X����A�L�.x��e���Q7�1�FWy͈Tq�b��񑘱q,�X~�+L�`c�!9�a*�PG0�z�)���A;���LP(4 �\�a�3���1~�G~��[�&a[�13F��5�/}�K��W�����)z珼�n?�V�7z���Q%45����Jy������,K�^Q��EҼ�+���) E~Ud�rFr��o�&�=�X>�^�'N�a<��_�wt�ݿ�z�J9����{i�i�� �8�gBL��>��O��L� b�h/��[e��_�����駟N�^�#F]�o�N�|:�(k�?ȟ�t��3t�����zk�J� [l�9��)�r*?���|�^纈��9=8���r\~�8ǜs�2�(Ɍ٢�lBu��͗��vs vi�y��]��p�hͻxHT�(����O_���{�_I��>���������l��֤IqI��Dj<C@ƶ�������oȘ0ߍ�`K�-��C��4%.���fSb7�{U�%3#����sOč���Ȭ��*Nuv��������3{��z�2g�	R���T�Qmi�3�EQ�m`J=SC_�z�2
�����hq cT�K_������\�w��Yض�ŏY>�`X}pϋ�=G�>�y���!$�+⋰����r�i�s�큔Z���{��0p�))�b� �X`a��s�P����Z�e��+�����	���W�k�,o��%HQI��ƾ���	!��o����Փ�Rr��@��0��s�HCI �� � 3~�� �L0�[���7(���(`\T���s��}򓟤�|�#���`'��V*���A&��Ǿ�]���7N٨P"�bӲ�DDY�pm�N�.oY��Z^g+_=邛R�l�����}Q��
$������G��~�D0�x�x�6�È1��\pL�v�U��@�}8��q��f���i=6<r��e�h���JF��Bbo��V��t��s���Cf�
����1��%�cP	����ñ
Q~~Ɔx�@�4<0�t�č���x4Ʈ�����ω�дN�#�G�G�Q�tm!ϔ\��ʾ�!$b�I`��R�]��e�/|���ԯ�ᠺ��@��/ぱ5C���V���:7T�����ǁ�+QG�i�s�������7��pBs��F�tD�$㸷3�Sa�FPCz��GS��� (&��Za#�(���w�(k�Jr��5!ͺI�%�6��j�^~7�v
1��P�!�D����Ȟ.�&�x��"��M��$n3�SpH��\��J݃�@v���bΞ�D�#?�^�6�C�[��.VϪ��\zd��sGy�3�>��Y1�����<!k:�մ�XXX�9���1䙄D/��R�SޣA��#�U�R�wrϙ���(����3Hs<�>W�j\s.�G���I�Y}�U�ff���9��ƈFH|��ƭ<~�s�˙�UG�]�28�,~�G��2?�1`B�^#Ls��V�˭q,�E��	#dv��O�u����W����Z`�
�hq������{�����4�A7A���s�|f�į�����U:�ܲ�A񄓄�s'.h:!���I2��@�݋^T::dP�b# ׏�\�sĕ��CN��ᜳi�IP�<���	����܅��$̎������(� 6��:���{r�Iks�A&p���1?��tZW�¤�V���r��Qw��I~�����k||��/�Ԅ:�bo���q��A�y�1��p��:?9e���g��E~T�:6����2p�����g���H���x@r[����a��g:N8�D��&t��|)��f]��_����;���狰�%�48�*D�r���K-�n��L����o�V L��O�6��Q!�Pap� gxf����o;��]ky2���~Ҕփ[*��X�H#�-�Gs��r����*��VtO�g�F���C�b/6�/Lƿz�#?���:\YG�-�]5i�`d�p̼	��ȞTM?Wr���C��%
N�.�����JU]�l��e�ȆZ/�x�T#�C����kN�>��8� '���t��ݳ��h��x�s��w�3&2� �i`8G�������θm�^��@��.���Uω�VWu���R���m���}�v��K^`|�Who�8�6����T�a�!�|p�~�������6z�]驪��b�*�E��'�hg���Q؉���#�1q�����D0v��Y@5����
�ˎ��R' U7��3XR�2H(dڙ��vP��Z�[�A���iZ.���
8��#:�>�jnx�7��~Q���~V�X�-�u�����(%�j,4tX��j���u2˰�"�T�6U\�.�_�V��"(��P���R�� �5���aPQ�#nqH��B��f��*wC�:�9(��:	�}�hp�Xm��oз��,=�ģ���O��oy�����s�Go��-��DQp��V�:U��R��E��g�����
9�gɜ��JR�5�Ŀ[(��=3"�s2��� *�MQ�@�kM����B��`�	|��9��;�J�fQV��+u�F_�O&W.�˶\�XZrA\6Tmn`}�+��|]���'�T�""��"x�Aq��Z����O���;���m�A�5����bj!qt~v�1@A�����Ե? �b�� �}i砬Fb�y�q�t"\�{�ohn�Lvr�^�n����㑷�����ׅ6b1� aD��(��v�YH���~��1J��Z���p^AL��MH�����������gY����U��&�ÈGG<�sRv�v�we?�߉�,�Ql��h�u���:�>�+�{��n�
4�w�n��ӑ��+�C���x����|V�xq�SD�d	:w��A�۬9��HJ�����m/��_�QyF�_y�NO�0w������!����=�[������-���zc�5�|��o������yB/�~^�����8" �):થ s/���S�w�Փz�����6X*Ѷn��U`�z��v�[�� P����l}g/R��b]jUB�#���zX��GeeMUO^ܝ��ݭ�	�3׉�I j�·`��Y�U5�K�z쒺����o�o���ǜr]b�!�M��	D���I�y<����cՕ��_�%�oj�m���~I�6��8ߕ��#v�:=�KJxs�.8��}+��*`�'V��L�i�^A:��;�jk��7���*�S�9���ߤ�U�����Ϯ8ʙ%n,.��s w1JE"�P�F!�����D/v���1�D���7жⰖ���*���A�Yjd��L6k��,2ts�Qa��|WܜR#<g�>,�yxi��SV�e�AVU�A��p����1W�W0�P] �$fFQݳ+���A�=��s�[ƈr^ ��i���܅\���o�x��+YIa�=]��b"�c��K�����.����F����O���J�\Y)3���U��X�>g��$߰]��	F�Ņ�/w��^�~VQI�ZR���JA��{ k9�e�pmI�.�\���xq��=~�.�r�o��` �i/$��zdP,y�r��'�򥨕�%����N�:RQ��뼇�6��j��R�&.,�$n�E?���~�L S�ï����ʡm��#PK
��us�A�5sM�6��$����|�*x����R=^��
���~^���-T�~D�a���_v��j}"�-�/��)�E�ms�m������) u)r�6�O� NWJ�XWA�/�.�~�k�6�����a�4�u�� �u$1R���u�,�m96��ڠr]8�6'��k��;Zz��2��;bo�{M�ک�Jf����ӕ��*�ϸZ$��j�
- �et��*K��[}��5��w�rWP��;n�>p��K�	�m/+�Vuy�����*�ZT�T�2�ӧ~��=֨'.��kt�ۢ�����_v{�`$�~t���&��u*2�y�T��w�����|�g�
��P+����p��r����/F|�#M��p�-|���[�h7��[�H=�]���_����ܗ.Վ�`c�Ɯ�)/�����3U�_-Nu�r6%q��rV/Ⱥ��^���2�zP�ŁQV"yQA^s�퇟��N�>��̠[���bF:%��jo��o�E{�4�@WA��4�ZW��@y��z`IAt��u���h��hT(t_S�D3�>y�=���9]�;Tk��@�@y����Y��_j�j]�T5��5'4vm��e�¿,5R|�c����7�ۺz���\(t�T5M�rU�l�������9�����LvMC�,�F<@��l;�UW�ץ�Y7���w	�]oPP�l�_��%�]%���� �ל�yض=	5�O�����5��5%ܱ����r�}J@�$M-�ei��6�M� �~�s�בP��<��������.��˳n+��e�v�Y��mP��;�w�|�i �kN*��JL���N��5��7[p0]��K���zێ���`��K(��e���Ee� �-�Ӽ��������Q��7(N�T�e���� ��-�Mݥ���ݿKqx�lJ���p�KR�|��m��g�S��h=�~� �ך�h\���d4!�{�ɤ��mJ��p�Ɔİ���&ئ�Ϝ}�)Y�Q��ئ���Q�p42����I�ԁ�	�&�e��+�`H����+���9��X��Heꈒau�~.X(_Z@ �q:��;wiv>��,E��]�U.�[6�%h���<�R=}4S:�M=����%M�sʲ�L�'�%ݔ�|��r�����z�9��NO��bS�zIz���R�F���y�6a�?-���\&��P��I`R��wp��	��l��Ih��?;���y��·���	�P��zQ�FK$���oޠ��~�g}âL��D3���A���.lC�s!#i�h�����^Fm��el }t�(_#jo� Ȝ��������T�̢��e��Qv�Fn��~�f�`����@w�my0N2:r7)�5 :��/_L����sPf��]x�?�sBӳs*�3H�fu��r~�x΀&\�>8;=���3����d���'6h*�^4�t�B�����|Fw^{�ʩ�������ye.ZʞcΤo&���"Z w����u�ne#!�i�P�sZ�S 6���8�s[�1��b�{��S�$�FC���&��`.Ϟ{��,p~��K�3mT#=Gy���`��=��l$�۫DrK�u��څ][�"��sp�tN����db��mx���TLhKU1�WF����C������w��1%����4�j�[W��@y�)�v n|�M�~"�K��ۆN:ˠfj�^A�N������$^�v���%O��HC�1b%�� ��kT'�H.��&`����!�-�_�:%#Q6���Nu#�w�(�2HR�$r�3=�5$�����tJ# ��@דP�sZ��\�<�f31�u��o(�����b.���hn"�0���҉�_@���j�j���n}�����������(胃[�n-/EԘ�P+�@�/�
uϖ��e������QW^C/�Zm��t���/Xd 5�b@]C@��ng��{�J/~� ��� g�\!��V�~P����(����IEGl��?_���ry^�9�lL{e����W7���b \><!p�+�C��R�R�_>K���w�D}q��U-pQ��.m��pց;)T&�==?�K�us���Յ����ז�jG� �׀�,�42)��,���c��g6$���3�ԭ��[�v�k�xh1\��F%�����ڬwݸLj���	�B�\�\X��5���R�,��mk2���|��M]Ҹ^�\� C�me9��U�� ٶT$�ղŃ���O���j����P��H,eV&�+��ײGnPU�hm]l��e���\���%�����0 �!"3��w�+k��jk���i�6�8Ǻ��A�T�[��,o�JE���:�ǉo9>P��/�
�G��U�J2pM��uK|y�+@��Q�%B<��#��y��sP�h�k��Y��b0�1w7Ji^� �Φ,"SO��f1\����j�7����ߥr�xa[��16V��������������[��6!�^��y�꧋f���2��{�E4U�h���_�#m��UnU@y����!lۓ�n��nN���9�и��ov�{K(���?-��G���.&����ǆ�����\SuQ3�as�져���w��겇�ske�>ꋁ�?@��S �0��YT(�-�f'����h�<mh��ٶ�3���v$i[Ġ�kI�چh�~M`��h �kN빬 ���&���K�g\_��zR�T�b��V1#��� �ؚ��k�,� �����3�Z�˂V�������"�.�f�RPs���b�6����Jqp)<������]G@�� �&����8�E]�\�w�v���QDKx�>��m��]��l��ji ��L�o1�/�N�=n5��N?���ZWMM</�v5�UxIW��A����a]�������_.�@ӄ�f4��S,���ݚ[T��(^b���HC��7\���I���
h��������FBl�����ؔCa�f�$�8��F<�|.����$V�������5��c��8ߠlw.���i��&n7�~���f#/�8ħ�Pta{8�0�<�g���"O��!X�u��� %YºwcJ�}@j_myȃ��h^��P�&�<US�8�t!Q	-�:�e�we a�|5 ��6TH`"���a��"�w[�zdj9�����x�.��w��i\�K�:��53�뢊���Bcx\��?��@
��XS���A�|�h �=�u:T�s�8v_3N��?Ayw��?d�a��I��9��x.|�f��^��0���T��/K��R�8�Ex��y���@ "f@��z��wS!bm����E�XX�,2]ܴp�9�.Z<�y�T�T�׎��8V���WѮ�E�
��.B(_c��:��e���u�2��n-�4B�6�pM �ʓ`�И�M�R�s�YV�^$]G����DQwT, q���OSpU���4.*&�q���kA�=��`�奬��م>|��� �א��c��:�nZ��[O��7��u��Sf����琙$x(1�ހ��u�a7\� �e� ������D���:jB*��n\8����H~>��+�\�m��+vE�,(�#�����4��DnK8ʞe=}��#�#5|����TXZ(�� �ך<�d��Q7�����\�FXR�m��L���Ax�0��cOlʀXg	�hs��ШtU ~_�8�RY�U�.�S��#���Q��s<#jǁ�|���J����&|�<������%�,B�ZSI�$Y���^��k�^4�׍P�����#�F� �:R�2�j���7q��ޱ���������t�R�	�H�v���-��l�{=��KɎ=X�S6q ��rVu��ˠ�S9�{U�����G��]۟7�v�=�GM�AF��>܂,�H���H|䅼+�i4�����W��K(_sB~9;�ذG�t砳4��y�t��A��ll�Y,��H8��Oh<���`�`���FL�>�@V�br�fp� fH��B���֊��-	�8��|]:����P�y?��98�h�Ok:;9�b;=�4^��e��3�u20��pe$;��u���)��np ���X���EtO���6�T��ɖ�\��ă12t@���?7� ��ܗQ�M�́�L���0�x�Ѽ����>U�,#����w�'��J[JZ+jr��l���b]4�BK�CM�~~^T9�xNvD� j>�KS�(�,��G��f�vzv��d�f�m� �ל�k�j��������==]�Q]}�`v �`8,�	//�:5��.]�����~�b�|����Y�'liN���y����od�̋�n�)΢��-��pZ�.�/Dc{y��x�����J?�fP𧁮�|�I|]լ�d�L�?Y����4��:AY��7�[W��e�B������8���F�u�	_���%I�M��|���i	<-�_"�`ᾆ�*�m|��*�-��(�'����h$����|�I7Њ:���z��R��$�e�m��f|n�ӂ����s�rǑ�*�s�oo�(7��_ۨ�뭶�*���̵�.����g_v���/C�[W�8�� �׎P����$��8�<z� ���9;�dH��? �&^���_�Y(\y۪�"��cn��l ����ڹ��кv0w^���\��7��q��>M�Z)�*,������ �ל�.Y�5+���*�U�HZ����ꨁvbN�o�Cl0\�Q�SW���[\8ѽᐕ�	8+�t����K�aO(~�݆��@WA(_s��0+�i�`����i���+f�/�<�J$����^��J��;��K�3��9���cn.�E_��-�U0�#��#R�͑O���MA�!	<��׉P��T�6��llQ�P�����˵�XM�7��^��j���]�Z�-��v�-����Xv��$��ȢY��_^�u�K���؅~��Д����9���X)l��f�V����}գ:B�^��Jb�m٧V�*��~wI����E�1�[�շB
X�_UEo��SV����Oy��b���Ph���#@y��h�h �h�=��h����Ph���#@y��h�h �h�=��h����Ph���#@y��h�h �h�=��h����Ph���#�+P���9�|iD=��?�����N�ˁz��k��^x�{MWʫ��6��G��(�F��\�p���|^��3d����e7���Y��eQ���/�e�Xv}��/�ܱ�8u��ׄ�,�v3r,�ϒ�؞�W����x��'wR\��MW�`��c��PҲz3����HW�J�Ƙ� ��뺚o�0A�W�8����I[��et�	��X�+2{W�:��ހrL1��v��ۻp]����N����3\l�99L��OY�,���$5A����_q|�ze����v��v5e��G(o����D��Ė�[�=���.>W�g�LIm���_���+P޼k�g%�|)�M^`���d���������^�W��}7{ �͵m�]����7�V��u���w��d/VuM߷��s)��[r�o�w�~�\�t�˨��Z���p;:�e�Y7>�=~꽤�֕{--���=�A�~���T^yٻi@y9-6��Es{��{F���Rr{:Q�G*����-�yE��7�����Y�����bl��QNv�c����.Z���6�����M帺�b��[�o�ؠ=�sv��8�V9C�,��%�m�/��+l�
v�JKY4[8�:�Q�ǋ�ށr{0�hҡ�7�2��������C��=*]ȓ �2vE]�c���MW{^u���v_�z�m�-���K)�OKW�U��yt�y��l|R�P��s��nh�@*k|�%%6��,)M*J9oL�2Z�x��gL��}4�w��僟��LLJ�,�).I�W�G�1u����ǂ�]��g��r�������6�.�^Խ,��Ҹ��n����P/�deA���L\+����=��;y!����s��&و�bF�Z�pY]�h�N�^�8\K|���� <��_�RgS�ޡ״=�Q���]�ɋ��.�ڇ��5����G�5
ƅq�5fL/h������S�FI�
�D��a���i7G�'�!����ɘtN��6���o'�c��+悓��^�r�w&bh@�C�7��`I����6�{�U
=�������x��[.;ZzgET��P�w:�dw�s0D�@��K ����m��4�*<!����YW�cf��dx*#�� Ihh��`�A\�0���.��Ú#K�%�L'�ff�ԗ��S(?� �a'nۈ���Y���{m�`�٥.veT��rk}�<%!S-��8E4>u�GGRYM��i2�T?X��_�r��w,��NU�e��L�#��gf��^�e���$��ڭC�Ȗ(�c�ɚl����}�kXpQ΢l05������\�ӎ�-\ ����@|�@H��j�5�6�S*�-9:F"t�>��>���#�My����'��v�Pe8�o�T 6+X�÷s��0��q�+8�m�,^�m ����z 믷�i0��17ky�-��KF����w�܏ ���5:Wݠbw(�R��!?�<�$�z4Ni^��
������
�6K}� �<X�}����g��H� ��a�4?W��XJ��ĦR@�w6�	���ua��aq)�2<ב�]s�m�c�]}F����k�z�˖��0�1�	O�=c��e�c.P�H!R,��h:���A$ͯDw(ܰ�t&�!�h4��`B���na@���.:&bN��
X�dr������	��7G��N�,�M �x���̑j� ~�I|}2?��'����D܎e��`#m	U����u:��|� ��l�4ڮ��vi��Fcs_��P7y��v�q�&π.��6	�4 ��t����	�����߮c��o|0��� h����1��s�A�S�����sgS:?���A]��Š�?_���<�V!Y�,	� n�Z:�y×���D%q��	�W�+����|Ng's���hz.��`��.v0����Q���|.��̃[~0�Ir�-+�Q���j��Z��Di�,�D��Iq�O��ӻ� ֊��4QV.�ԣŔ��p���� f��<�����l�"1�}|��I%���W-�]�CkP�-˘(�"U�b#�bފA�;^p�$K����E���L,�h�u����tr�./�\_��=�&�����МH�.W���W匹�ۥcuE����GS?�
_������ZG"�8~�L��eS�� �I_>�s��'�g�ꋕ��'�Nb�d4��&f��8?����1�:��%�a�2\���a��X���ŉ�td3��A�p�Θk������=�>�~���>���gЩ�U��	�2(�<PQ�qI9e��bDcu��{�9 P:�z�sDY�`�.0���gX�O�Sf�)s���	�N��U�muL�I1�2���l�y�.��/��	XW�N�^D�_Y7_��<����Ow��F�b��і_6?b�e^"+$O�kM�<N#C�2n|��9��b��xF����$�]���+e4�R;���5a���R��.��2@=�eP��q�5u��]~1�%�(�"��t�� 2D�$趤#������j��r+`��Ȇ?Ap�� q�cq�ʀ(��OgT����dw��0t��˸tQ���!\>	���;&&~��+p.8ڗg�z@YK6���ܘ�%m��T���dL��$c�׾��������:��\��e~�Q��¦f>����YI�)�`0�Qs���Ν;t|pK� I�Y��72��v��f�N�^����/��+�B^��q��j�b�Jx�s?�yy�&�����u�KRwmn�O6{�K�� ����la�p����)l�/��)+�	��u׹z(D�E�˖�*��z�#�(�CCr�Qu͙Ш��'ぁ9���j+n��v�Q�$�U����]/O3�9,�`(�N�#����B�b�F���/V�$\T{(�.e0*�{����2e6p�V�;S�>�\�Y>����cV!���k�:�Bu*��ܘ���]�1���TK9�_Ų	_�̢se���;6��</�M`Kh�Ka�	[m��,.X��`�p��y�ੌ-K��%��?$!u���z���!3���g�vJ�|0>�%����SP��������8P���D:dJk�x&
R�2D��L��(w&M�9�2�3�0�V��&�ڡ�VGi��In�z�x9�9��zB1�R����(c�R��߯���Ck���z�v4�%�)anc�a&�a`��Tō���x�\����qu^0���D?�\��9Q��}�/O"F�mǪ"�wʆ?ё�P�]�,馁�������/���1��t49��ƪ$��~Z�{�7HX`rQ�( �&,Qa����7M�l|�R8h����^L�Ɫ��R���qٍ	�;���P���,Mp+��p���mW6�����B������1v<C�iS�6~>d�ߞ�XuϞ�ނr�CǶ����m�J�!�6 /-!-�e��
�˩��op53l�ߒ�G�2��W���[CPP]�`�&1�U��l�o�Vq��a>�A��_{��O]glo��dc�Ӆ�j)�A�U�Xڮ� �9�-(�)^u�8@V�w�/�k�ǽ��z�w?]wZ�M^nT_���e;^�7�{�	?�t-@y���⭯��"p��_�N]��.�+���]r�s]2�U/�~?��ݠ;�jq�$ʋS�3��F#: �zG�Y�.t�@Y��lm���(��XMҹ�g� �};	o�1�"�:����}����(�ّ:��@=�To1[ጻ�Abpv�t�]�r_PVrn@����`L�$`v��C��}��h�Ay�K�y�*�!Վ���Lq��3���Q���>i���~�����Q݄�`m�k)���>{�H��:����h���dV :�}���a�:_�~���m���K(4�}B�5�1�9Q�fsK��������O��Y�;H�74��@]cچ
���x�4��@�G�=�K�b'�c�y@�]� �t�ж7��:�|��ڃ�XS�� �7�@{@Ι��砢�:�[P���S�qM=q"5�U�K
'Q6"UŁ�9��$�B#hy5�H��6��k:%������F��:�\�_�P��c\����D-I*�ft�Ui�̒��k�c(�2�8T����_lh[^�2�%"Th�I�f=#�V'*���Ӛ%\~�&b4��E�m��hl���#�ǈ�����W�P���P�ڞ��#hwbh��_�d��]���%^qNv̀p[���"�Z�3H�3�#��Z������UN�e���q\`��;N����q��e�c�!�/?�#�>7O�zƚɚ�@���3;����ęRʐ[��,�L')��>�ԿK��s�V�G�x�:�^�[w}���N��qp �\���ߧ��SBb��s�u!;1u��\HY6:qf
c�l�mh�G 7Z<Q�L��r�SrƂL�[˩`T�JW�V����7�#r>�=��y1��.��鼒5���n�tZ��K�{y��	aQ1����$R�p��g�X��'8�}�� e�&��ߐ�	AN�0K����а���e׀���*>�e��F8��䀎oޠ��!%YJsD�����B;=t����;q�!�n�X8I��0дX)^|=dO	͚�RJ�#:8:�L�IHT�ن�_�oM1�^�����(�g2�" 7R�����4>CT���5�����������!�Ն��kcR�M�.KrTd9?��?G�Χ���!�d�Ķ��ӌ.wVƙ1�\��GGGtpxH��I@�E�X�f��l�Aj��/�}t�|����9���&IԶ��\� �]�h����wdu�,a��m?9:��_<8�?͚�6M�i_h�@����w�A�V>��c��t>���� �����#�� ���3@P=�u���}_���s����2�i�d����M�y������k��~L& rI.���/�B,�"�p�WsS���5�=W����9��f.��U�O��JV\r���X?Y-$ ��-����IG�H����9�y�^�S��
�>@y��:�Ӏi֐����m�;n�@��<ޏFTxN9�`7/�!����@m��]�S����rM�� �,�����M��X�!ë́���оn�{PF�#��<�Yz����aQ��Ut/�ek���s��1)0�SΑ���C��<�@����~�r�,��\��P� ��|�x@�67PxAD`p!�&;����ΐ���?1���F���IH �ٺ�
,Y�t?+&W��Z�k�bn5����	�R�h,"s��
��\l
.p�P%x.m5���MQ
�b�,X���!lH.��.����GoqBcNNq��}�_pyI��N��I�YRH٬Gj4�2�'�����*l`Xu1��F6��ُyJ]��~�d���ImE�,�\�"�2�J�ُW�C���Ǔރ'��P/� >]�Lh��N�f�h�<pC�2�l�C�>����^
��L��SSзz�
��ӱ��l�Y��oY��UT�^��.z���$)��|L#7��@�u�l��r��u�;B����������ڧ�� �d!�I.k.��C�����ȑ�&@��~��_p]J�h,:�4�I���\��V7�-(+A'X�i���Y2���s��ƌ{y���R�.�P��s�Ā	�qeHl��[��]�ͨ`���b�j rt��6�e��<,�|�Z�eZ������i=�-3���x^�70RmJA�_�"9%��&�KWY�~�i�4	�_|Tz���Y��g�)G��.��K� �c�tU�vEmUeP����A��I#j���iih+�Խ��e��&n-!�,������6�,O���e�t���yˋ��~!6k����7W�7w2�NV&M�f0hː{�]\-��k��m�k�6�����l�n|t2�8y|�h�[Ѷ1��`��ڥ�U3�q9T��gpk���l��(#�,`1zsE^)P����O�׮�j�`6�E&I6��]�-�|k��8:�G$���E�uA���K�{Ɋ^��bO�����=�A{
ʑˏ �)z�ɝ�Đ��/x\�Gp):P�}�W`b�,׺˂��_Tv��WOe!`�^)\2�kA���iy�*ɥS��ǜ#[��[�F9�O�"��x�+_��%�F"���+
��:���iX^{a@�4Β�Tc1�����T��	�`��Q3��}�˘�	�}�������j]pRc��A֝]�]�,�NXƉD�f3	����Q�X�ŏ&�ϥ1CVo�z�ĊQ�Ua���&��x�%��]SoP��!�jc�1�=�):r�AQ����qAt	e�y�:��h��2(�R�`E�?���o��r% o����$�L�* q���K��=4b|`s�3� ��񫲆��2�B��3)�"�62����ۄ*�T�ˀ���k�P-j�/Hv��c�56�eE0q{9�L=�uA]F�jhu����L�WjY+b��]�E�$��c?8��8JG�:�Dئ0��?`p%��.>��Um|YN�A�������H����]E�/�Wʑ�q�	�y.�r�����\燹K
��Ɗk�݋wǶԶ.�َ��²�u��u���'�R/5Z_���y�������N��ޫ�ޠ|~~�16x ��}6�U�:�/#v��DT�h;2�AF�IFi2�<�T���G�څ�^�"��T�nL�r��`v][6iMK����h?O�k�P��Vn�Y�sWY���[�E��0��k��y�s�-{Ͻ}��_q`Q��빸d���i��'�ʣш9Z�c'��_�O�?��8`S���4�N�H��>�lڳ±*女�9uPcZ�y���2��b�_F��_[��-/�Wq����oF�A��z'�C�yp�k���1[ja���F<�`<a��i�(a0�;����z��W���6���l�],��lp���
�Zw��#뒣�şpY������>�疼{��Ժ羴໬����`f��5�=zSoP�wI��G���
��H�E�$�l��y��:u1w�j$1#�Φ�e��w}_��ѱ�wb �W��v䊁�������Π]�R�[�Xǟ}�ޠ0��[q��q����gF�a.y?=V����A~t�^s�n�LV����jp��1{�N9r�rltE��|�f���$�A����U6�q��)oh�_G����sFgǼL_^}｣�=�V߽ ��t��
!M)�
L��޻v��7(�N���=99��|�#�+��+t��-Ve�"cSq{+J��Mi
?Bʯ&�����}�^�Sp�8��C�"�E7����XGi:�Ԥ��q���DI�B����{�2 �c��x�����O�ӕ�ܲ�-����;MGt��]�u�!�S�g��I>�7����;����^���=g}��ܩg��1�O��	�xi`�~n�M�)5�Үy^���]��
]5l\`�H���O�r��h[��E|�W�<08����,|�`L]��O�l����:�����.T���@�A5P?�}��`���8�3�O�3OsD�2l��!��@�e�_���H�i�����6V���F�A�pEϋ�^�?��?���$�q�U�P���������������:�;3���^��4�'�A�稭�~�P���,h����UǏ�`+���☮���o�����/�+��R���*�q�#�<B���N��G� �o�Ϳ��~��4�O�D���Ô�x�~��_��7���H�]˳2�l4�@t��V�nW��P7���7���_�\4�Ce����o�%��c�=�q LZR�dsD�ݕ�:ȨP��� �E��<��@t��VT5x�n$��CUPi ^ƫ���\��|衇腟����s69�lz���=��Fv�5�V4�@���5��A�~��&�{Tu��Ï�ƍ���۷���M6����g�C��J* ��t:�r}�@4жik:e^�;@W�Pe�.?T�~�{��\3��w��3e#:�Z��lVk �On�m�3h���_h+:euqw�#t��n��L�M$�!H��3��/�忤g�y���|�3�����K|[[�����y ��3��?��W��h���Gi�7(�aw��U֌�����;~����'���}�c��}�>���;���_~�e�� @��o������Av<�Ǟ~�NO��<<#;z���7�
�4��F�AYz�\1v�8�PQ<�����O��?�^PU@�|������}�ԧ>E~�������}�k_��N�~���[�������D���Ƅ�}Sh���_h+������K/����~��_�5>޼y��@ª��sVi����?�C����=�g~��o���G�����O|���!:9x��~���_��щW�F��m�x.4�@{D�A^�Xյ�����8�' � n�q/��g�}���կ���E梿��/�c=L������	���+g���7����R�>z���~�ޠ�8`� � b����3����͜1v�}�+_��9����1?��g����DO<�:-<��z�~t���Mʃ;]��#+�;�q���~����X�'�t�PG|���~�����BF����-U "�Y_�!�]��տ�">t���ޏ�7_|�~����֏�2������?���a��@t��V�ȇMP3 t��'�j�ԃ���@
��[g#rEN�pL��-ʎ�tpxL?y��{�`��;����,���,�Ͽ���h��&���"��MC����r�j�H�}���W��tP��u�_��/�+�g)2�F���b��(��Q�r�F&��ɘΦ�4/G����Gc�α�/��b?w���!q��R��	N6�l.Ɯ�/g|)���2W٦�c����&�&�:��V@Y�)ke4�fۏ�}ё�s:~��>-�_G&/����7�x�}��W����d�Y|�}Sf'4���!E�@=�̩q�4Q�Vqd�	�(��k�1�IEպ�ౕ} �4j'S����!p�ԃ0�$�������;=��6�A]��<, ~Y,|C�2�eF��z���Y�U�e�2�e��ٜ ͠�K��!��f$An�Nn=󈺨������e:�M����Χ���ɈfyN��[�E�G>I�}��+�t���y�.�ٟ/]����h�{C������g,۞ࡕ��fT��b�a:Ǯ�3������C�����wx)�LҐ�3p�֯\S(�i�Ktv����;���c��?{�'T�1��r��\s1��p@�z`���ʟ�'�dL�h��g�����s
9������oY�n�����I��
x[��B�d��2BB� �;��A6�"���������?��`(L)����4���r3e���w��`
Y���`��R�A���~e��	!�}�%��cM>=�R�jpЁ�ܧ8:[1���C7���c7�r���/\�-�S:=�M�~�s�O򎿧���$��;h�fT&����L���%�@���cÞ��*�& ["9?p�%{Ē�ɝ��߆1��\󽤭ľ@% � e�?��S�

��4PhQ�\�K��s�=(��錊����}�9zۛ�Nw��M(����]�Py��HbT����%�/�_9�*l�jN��;���3K�n��NP�W�x���!z���ȧƾ�|�;���������?���+\�3��1̹�U�����In�����K't;���!�!�ݣIƍ\��@���Z@V�ʀ��
؎F)M�AG���<��윾��o��r���$`�p8��]v?q�1���PD�����Ou�v�J����X=�U��s��GoL�;���Ȍ��C�=�<�z��'h��\bC���K�`Q~~BV��)�'������f^*%�a�?�X�
��1�Gρּ{��@p��}�{;y�[�r���=�J;g7Wz��8���~l���L��.�b~�NΧ�{ ?e~<���Oy��R��
�L����q4;�C��_��;�d9Ki���íkA<P;�������3t����78���-��d���܋�;J�	M�1�>�My����?ћ��q�%)���}H�:�V�4�@�/�E�d�BNY�1����7��忥�|��t�����o;�JkK�	O�Tu�4�v��O�2�Z �5�r
�v��%C�Nٟ�5���O�B���ӛ��v?	�Cʒ	%^.�#�URl��'����ߩ�N���{a
b^�)n�Y���X2���+��y�n>z����{�Q���B7��C4 Hu�q�jl,Y��[$EQ���t�;��kd���*wÎ�����~�z��s˧w)��E�M��v�h��J�Imp���\Aӻ�ӭtNw^�!}�/�H7�`��S�8�4CL��S�:@��9_>�΁p���ƿe��88r;�[F|�{'�Qs���t�tN?���h��;����4��4�c���V�Uo���{�����Іc^X�+x��Ǧ"��޳�_�g��r'o�c�ܠ���I{�%�@�F�oa̋#��٫���JVu�t����n1,<gl~��814Ǝ�����	����}(9���1ݤ��9�t��lF�]X���Ǻ.���7���)y����mѪv��7m�m��LY�lk7�^�Й�}�cW�����Q�s��=���\���rN���	�����o��?�7�<P�8�������5�ʼ�`�Ѕ'�������M���PM�Cf��SY��8���Aن #��ײ��(�;4&��#���ͱ�:+�<yXv�� ���V!�Ɋ�(�r�1��y<t��1I��p�IP�X�\�wp�Z��,vZf�9����rb|�Yr��ǿ�cf:���Av O#*f����B�����&�+�o4F�n�׿�/uD�Y��B���}�e9G}���l�cŔ~�L8�X�w���������/�n��9I���#�䊹���.\�;������s�\��Ɯ���y�2� .���G��x�.::nGqP�B�ɻDʍN�D�3:�:NN�G��3�����ґ����gS_~���S�����(����~��ſ����|��)W��F�U�?�( ���Aلm����7��d4��|ͷ���+�����y6��l��#�M3�wϧ<�)���pD;��](x�4ʓ\�X�g4�ώm�O�@�	��<_���p�g�3��ݑIo��)\Y�u�����y��>�\��\#������,��?;����I7J�
�z�k�,������m�/Ʌ�	�cy��PF���|*��3�ߤ�#��H����s'|�l���e
`���S�˟������p�\,����(��W�?�Q����/Ty؛`��2����\��[d�����k.���w�:-�1Ϗ!�1��|J�甏3Kw_x����oџ��G�ݗ薟c�ӻ�{Fn2��ߓ	S@��WJ�R�\�~�W�>���y��l�6�/O%i@!��7۰[҄�.�#�ґ?y���w>J���³?`�E���3�Gq�y�ˉX�%���pe����JyY���ޅg�¤�*��%i��3n���sT(���<�u:;?!�
���(-~�E�^�������%��1�=t�����4��08�������Tje�1"`B�$�:w�ګǀm�?��O�ҋqhG�G ̰����t#�:�{��@\��>��E�����-�2D	m*Ʌ�,Q������<���U��s���:�>�ƔمT%K�cd���FTMc� P��Ԏ������������Qz�:������>G��3z���������� %�y`h�G���!S�~G�������S��"]}/O���.��Vc�K�������Ss#��S^���O������/W��ȓt�w����o�1߉�Ι{U)��U�\z�e2�@� �;��C��Dm�O�C���닢�҃^��[:%A����c�����P`a��_��b�ė+����B}���hY�]hْ?��7&�l�䴻$���`o�́�Aߡ�T����QǺ<��K��t�E���p��D}�TR5Uy@�R�E}G�n�c��ۻycl��HlF[鄨���q�M ��Qu''��h��s:�R���Ɲ;49?����/џ�ѿ�Iq�x�%<G;����l�1�q2�|�9�U�zB�|�9�^
�1�0`1�4Yj�NG��"�8N����<�M��c.�Wp�6c߸�F~�~硥_��;�Wߠ�{�?P�X6�I�{�s�E�)�A��!�����E�Y�F�KP��e���K>!�yn	m��f�0G�fŜ��t�E}���Ɉ}�u���q�s����T=j��* g�"r����>J$���e8��'1<j�./;�E��軋�SoЃ�X%CY, ��EN&,!�/�N �B���᳏4e܇�RKX��Sr��=l����"�'�_DQ��T�ޒV/�B`�;�$q_f�o��Tp�FoH����-]0R���s��:�s����Ώ~D/|������:=������~��-��ˮ�
Gc��2{� ��j�g�%d����>��**\_��yXDAYT��i���܋UBD*=�".����z�s������>���y���?��͈&~��C���R t>C��U
c/m}��
+E�}DB�?\'I(�̗�p�Xu>c=��;��IH��;�.Ց�Pxߑ�����̋���BF�_&�粦wL�s���V��Fy�Q�f�C3����<Q.�����O5fr��()�\|y:�
Y<!����"-��lg�t`����<�б���������{`?�~=��k�ɖ60Q�\'ss?��e�r���h�ssGՖ�-�^b�V��nBFG���j���D]�T��O)��J����}���_�B�O_�G=Cc�s���!izP�9�\�2�=?�aȼİo�*�E3mxpȪ;���_~�����וF_NY�je����@��%g�F��=ǅUߤ���������z�>�޷�y'��G�ǯݥ?�O_���M:x�a:M*���Frf%�>�KY��S�z�sJ��p1WR�5�S~�����"�{�����~�CV�����?��3����i�\�֑JD(&'�hμ��%����I���$�2�*���f����|<(�D�r��W^y�n�TТNpN�Lۤ5Π{t[ eX����I���ii<)Ӣ�}�DIL��ʼ�tvvB���~��R��݂�jR��l&.� ��{�Kg36"k���n�ʳ�� ���w�V�[pcuʷuC��ʅ�%�b���b	͉�xvr��q�r��?����o}�毿B?���t�������^�U�&�t����$�:����ă�T:��*P�0�/U���8l~�w~�>���.���10�QKT#�ɔ��[8yj�H"U_�7~�*�o���d����3���;���������7���z�[�G�&V����_���QuȘ�hG��Ї胿������X|��(�֞�P0z饗�K��6��/�z��`F9�e퍾��@���i�����N�򰒺@h�o����/�d,�-ꢡ3�������(�j��_��fG�\@�ѢN迏~���ѿ��}]nj]�] ��X��vA_��'?�?�O_`W��ث ���!b��s]}�Q��g?K�������5N��
�{�W�_�ǵ�T�=�Wjc5U�ظR��<2�߽}�+?}��_���EOM���G�x��:D����IA�QFSD�;���+��ұxwI�>��/���"U몒�r}|S�/�;0@�������-�U��b�'����z��8^�����G��h�W�|.*g3g��dt4{������_��s�������N���"H2~nA�����P�a|�Q^|�E���>F��δ�Zk'��L�{��Tm]x.�/���扰tu0=��EBK���j�1�������s��?���7�JiG�����2I�vo�_���C)��d/����B��δ	��̲׶�X7m����~�ӟ�/��Iz�1�\��ajT}���'pɎ&�}�O���{B��?�H�]�f�����_���6�9}]��*E���7}�������8��C_��ބԴ��s=K�l��,�G�RJo<N��i�O�g�1�O���s�����ޅY�Fi�1�+#6v�����~����5V2��7�x���58u�ɋ���N��a�� s�ް=1��u4?���6���o~����/�f�K��.ը���#V�"a���*�m?H����([HP��� (`�eJ�tJ�)��袊�H��*��%)����zɗ�)M����JP������Ϙ�����T�QI�25�2'�X����5_뻾����:�3 ��9�'��ZX�!Π�0̠ �#��G�<��oy9��NF����OO���]�bM��ps�!ϡ��$�M%S2�uH��S��$�s����霎��;�u�s?)�tӜ�#YN��|�����ӹף��W�尸[����*
��R�X�7��|P��$e��ټ�AF���D�����UoO6��x1�Ν;=]�A9��j,�L�ȧ��m|���
t�WL������7���h�s�B&،K.��`�DP�/r�쑠aKA*n��p�]1����^RR6g�Z��+=ȶ@����}�Z�'%zŗ��#P�'�X/K"T�$|'V�V�yA�s���hO݀a�����������[cs�H�pz�:VI����^j��q�����M�AZ|�nQb>������B��Ee���S\�\BBB���v��5�zR�4x�Dv�r2Q,���r0��<ۉ�i���@�����c*�����9��O�����D�=��e�q�v ��S�}2����Z�\5xU�QuB�nL����Z�Yd*�U�)t��*g�4�<˺2t��N73Y�	��S8���*�X�1�p���W9�_x�w�i$O����~��_h���ঐ�e�bؖjx�T�?2X�AF8����}�ˉ� k̂�m�(���`��(��O~l�RG��!	�;sDV�e��R���DT/�@���u�k���~��㩿a�{.������ܷg��|�[�y�=w�*����1��˙�~H}yli�q�g�p���h�{�=��������6��=x��b�R-����A}�~˕�����*�����-3h�cč�����dbI%��ŎR��Ǿ�k�x������ac�/��Ue���9	� ^��2̹����7������T��m��P yVe��<?��J�S���\[ZJ����8L�T s�y�$c�e~�Zp��ƣR���#��� �OV��w����̜������S�+|�q��!)o� đƎ�"���]�^ЧU���T/.��;��{ʻ%�?$a	�xQ� �4J�$ $�^���d`�m�o~�a�;1��21�C�e�@X�?Y�nV:x��<�'�+��M�;���#��c�g�7�r�ϟ�Q{fR�����g�'��B'1��%����RC��k?�ġ�eAy A���b�H���&|�r�h��mu��m��G)X�Bɜ1ڿ�x��|��ݺ�6>�X&��:1c_�1Ym���'l΅��ӹɢ�
�F#Nj=�8bp�7�@����1)�,uΜC:�C��pOi#�H#���:��ꋚ՜SM%Z�[���UNYzQz~��ޭ�tk�I4́�A�q$[�%�].�������X��Ds�n�ܹ%>� 7��g�N���Q��#�%/�N��k�W�c4�A�םX������ز><ԟ��Q�_7΅��1'X�)�MK ��8�j�@)w]ɫ�^'����A�wa�D��ƿ�������2�sL��Ŀ#��^i6ta!SoXi%j���\0�����pTI:z�i(޶��"cI��a#����V1G�8�nC���D�2H�;��=����u(�` ������E�F'c�Wu���i#D�E�,�@��>:3���}WV��>�|��bQU�_��y8���qFsw�RH���Dv���3#��l&�)��Q�2~=�E���pʜ	̍����'����c����K�\#%�A��UT�庒�9c�9g�D�8 д�8�WLU��C�� ܽ��k&方S��WVr��w13���@o�������X�9f��dthHl�����Wj��eVFzF�?n�E�uf��E1{�)�g�Tx���.�O�����&�Ve�)��0OX[2�	���Py'�%]/7�Ѷ	�B~�xA�O!K�*�b���D8�>�%6�]�H�T\(��1��F��[_���Z��R��ڌu̥ܿ�ؼQ:(P�1�Z��O�3�<�K��$�Y�c�]����bV�ݏ��q�r8���^|D9� _\�N4���L�z0\����%���!5�]��Җ�t�S=�si8n�ɦ�e���杲ta�lQV]΢���b#g���}�Cߖ�K�t�Vڣ,#Β�o��������'OJ臜�v3�1="&�͜�S�����̯��8b��{����_?�U��'�3���|]����b.R�=��5@��E�wEu�{�)�4���>d#k�ń�Uo�qK�T��a.y~C��CPv��Iq���/M�H�����0��~WR?�md��c%:p\�I#��ЛX�U}�T[莵�Ļ�&7�&��O�3�Ã�Rѥ1��0 ��YT��@��~I,�%bW���8[���zbtʦ�w+�//� �1`
df��yp���_v�7�����z1/9F�
q�لu���r����4�G��-l6�d�Ϙc7�׍'4bé1@��g�S���H���8��?>�WF�*���+1��R��b��p�	���Y�&h�#��fS��mC�]�d�V�A"n�,�s��ȸfN_�6l�v\G]����U��^#�b����J(V���`ӑ��0������:�gL��c?�E�9D=�L�f�*"�3�*��2�LT�˲�к.��f����A�V)�ݕ��Q�8ğ�\ڰ�mP�	m6��Y��>��G!C�Wqc�t09�Spق�<#�{�V�o��`(�����6k,2Yj�i���z0��>�9��w*[bq^��>J+��;���q�v|Էx�Q�4x?��(g�~���X��a�i�$,/r�����E�u]����t{�l�?|l�����^V��#�#����d���l��~�+��e�'��T��m\�	D�6��rW�{v�Ø���������<b#��3	E�A�A�ۋ�n�G�`Ŕ��WQ��ziai/i�}�J��>�QW���]߷E�s�,�� �K����E�B�[�(Ӻx�:8c�C|4IWL�{I@��c�Q��]���R�Y���q��č����]�u��ͅ> ����ZV����p��(�j�P�9���j�Բ�w�n�~P̄�����w��������F��(��O7K\��xo�Nju��d�y���V����j d� 2H9����T�y�]%�s��ʨ�1���aL,�po��
�Vs9ƀ���}��wW�w(�jl��\\MyY�0-�!	�;b�x�sDI���}��Po����9�cB%�,Q�(ӂ��o�w�������BWV�NJ���D�ԵKNE#����s�&�1� ���v�jN5���A��uP&��P?p���/�
 ��8 �0�g�]B�9��]��%�K�H�^(S�xj8QO s[���l��8lf��!Y8��mlQ����ͪzj{�x�t^��PUV:��\l����.���c��QJ�6G?P�6�c�R'
:�!�V���1g�	 ��ׄ�z�&�j_�3|+��c�6с��!<�������i������s9|�Y���G}���]4(�r�
|Kx\+�@���Z�w��Q�bU�]��(�rƪGaܼђr65�u��͐(���v��e��G�o�6�1���)���G߿��ﭢ�q9ʼ��Ī�C��/��ǝ��Z��f:��֎��J��TI���\F��@���*���u���P7���&�Td�}�wE��x≥[؛m�[n#�ר�9^{�5��� �"͌҉	��+X�D���:�mQ��Q������5a��b5�c������q+^�ڪ�k��.|�b���`|օG˹ix}����>�.��xl�������F��i�}qC�{z��gY����˸ĭ�.�F<�_~��\����ėA��kR�/&��?�qԟ�ٟm �*:Aĕ�z�)�g������}��w�[�o[�A�� �!�8Ip�?�s?G���.�:���������~��^���������E]�P�}@��ɂ�6�	�y��鳟�,}�ߤ���X%�.c�E�G�ȧF7eJtQW��Ha�
(u����u���Վ�s�Χ������;�����6�՝�Ɔ��w�wy��umd]��ꋨ+�v�pT-����j�Ţ�.
:����ơ� (���H:����-[�s������0Oj՟邵n�� ���駟�7�����g��?��?�/(�$,M����>����,�q	��b/�������0`�\��H߳�+���� C{!Y���E^�u���cu���U	i����<��zǜ��T�|����w���&��c�����U��N?��+�V�C�ӛS;	���AqT=��#��~W�����a����e�o�ю�3z�n�8tg<�ѱr�A����M�������D`��T��\�z������j�kYc��>�uR�ҁ�:�:88�O��ՄV�t��/�7��M���?������ɭ��hC���z�&^�$�Y:�Q��	�L�VkCcf&q;*�����K�D�<�}��_��NEb��	��鄆���g��&�1��u{�;�����:�"��16�8����]����g>����o|�ˡ� ��V-b}I%\�+m�j,��.�w��+c���9`ݷ��6���n.�ʹ誊kjB���EM/�'�#{����L(]�tr�3&�#^ ��M}I9!�k�^}�U��~��?�Z�Ĵ�ϖ�ׇA�������}�˄v����2R��J)ڿ꾄:}��`����X�YV�Uu���h7 =���;���}�T9Q����u��b�*.��.<�}�{}��>Y��r��P�[�Cc�Z��7����w���	�uW]����m)��<�� �*"����8E� FE �:%8E�����c$J�h�� �E�̃P���C-my(�>m�}�g��9�w׳�9�ܻ�������9�{��~��-��q�0c��,'vW䜆�ŲV���x��ݹ�%ݮ���sł�YC'�!7���9�Yw�;��rkؓR�g�!���GOr�˹�D[��8�]ѻ�����لE��AVzЃ����7�'"�AwL�0�p���zr�]t ��c����U����[M�O�.<�-.�j]���z�	�g=�.pFfıM!��Tm\.}�4�y�Q�zT��)��#�M�Qv�:ǲ��^�i���ﮎ���SҌvgM�E]�����ko.Xt"��ay��}�|�'c!)kvP��������2�!d��$ݽ�
i{TI���=L����$¶��+!�6L?O%�z�����1�:����O~򓋇<�!Su�!�g�m[I=JG�GZ��-��c��;�_~��6�H��u�f̛@���g�==,��~�(\ͺD�b�ܪ�J�.��b�Sc�(�h�o#%��=VKM�zU��'��(����8oa���uh?���/���s}'�����A�Y6En�5?Ѥ���W}��=GS)+J���IC�T1���zֳ�j�k_���;ѩD��2f��y�җ����\�����2kKwj�NI� p���,6HY�kF���F	ZG�~�I���Q��p�Q����O�����m��{Pv�z1J�r�<�>��g��¬���Yg�U�[���hG��H�T�a�I�O|���L���%�6۬��ÅcfE�C��;z�h�}|���Km�=�0aĝ��e7~U�����ǜ���^�29�K۔%(�UNUo?!ON�7��{�d'Dt�Up���?��?\I����g+�jo�JcD}/�8���͊�@�/�^,����tL�V�aX���՛��&�j�]tߨ�r?��(�<�(���M�@�T��%��G�v�	��ВX��㗾��i��%����ߏ}�c+'����$a����<����6-6
/�`����/1Q��.���֛$�e�Ŭ�kRs1U0j����k�[�9[�tG�Q�Վ���ф a)�5�Ǌ��+�v����LTs�<ND'j�?�+��4��9�3MvD�nw����p{�6�6���B�Fm�{�`�<�%�|lOT�׉Z�<DBv�C��pO�X��f��q$��]w�j��{&.b�����HX�Aܰd9ڶ-��0����ɚ桩^����ɨ��/�����\	��q�F��1��h*kZ�e�sL�	��6���W�bl�,�u�`�}3��V!q1ָ��$TJ�9� �1%P�$���%nJ�V��  :ܰ(��c�d�~�\���DZ���a���\���D%	1���Dɍ� ����~U��f�I��F���.&����F�������o}������q�����ĉ��	�6�#�h���&QF�N5��m���=�ܪ�W\qeIl�U�_�3�n�����ǫ㭪vܮ���w�[q�Ӿ�xӛ���T�g���pқ�����O�GPm� ��i[�����ʻ��yr��(�k�ȶ,�ُxdq�#w(n������7O4Bߎ�cs��s�Т�����5zF}��-�V��ާ�W\|��U��IB �~�u���LY�����C��JZ�M]�R͌r�29�ic�>M�S9V��۩�4�W�F�S��^���q��O+���*�4�P�K�b��o֍Z�9���G>��^xa�&���A��3A�N,�zgc�4&9"{��?x�@���+!fL
D59J�kUf1�M��"�`� ޖg鳟�l��-%u��>�4C$�����& ����}�F�Vi;)R�'��֚���'H�� �7kֈ�r���,��Vxf񠝸�����=�����K/�����ߛ��c�#��Y��4%@��B2�wԷʢv��1D�+�%�t�p�E��>��=D���/�ğ:D�X��yڐ�k
b�R>��E-+j5j�
`j��O̒��8yI�����:!���yÍ#H�ЈT�q����D��2w��vU�k��7��H"A�b��3�ָW���S�O��1,J�6�p�șU�.���+����%	3C%EN�c�����ʄ�&����09��fʥd��"9ۇ���mK�'%�HH���wT��.;�R'��,����@��$�����A�����v���k��J{馡X�گr�5�q]�2c�ږ$��8�0�`_v.��A�:T���юl�a�񗆹��M��w>x�H�M161�E_Sj^�X&帕8\;i����ô!�I	�ﲢ���o�X@H�@��H�<M�D�@=�6��eL�ib�^�V�n=A�+�&D�������t�A���h �����H�-ǒ�d�����l)�Hú���5�VUK������z�����D�b��/|a�-y��I�{`5��v��Z]6T��[��al���>q\�މ��Ci�6�=��K���/N7��hϺ�^"�YJrM�s��3��D�}�Sr�����I��h�t�_��:�Җ>��˫9n�D��*���	)������y�[�R�ɟ�IE�J|q�_IrH�z���u��[��F�>J�Nck��lfa�R/�4M�z�N�a���G*�8RC�8��	b9�(�����L	Oɴ����7K`���y�U_i$@`�"M�Z<�)�]S�"�B;�R�N��qO$~%K��u1���q�~Q�/R۲`�����q�uV7���t�鷛�y�n�(Nm���)0[���iM�9�5t
#��4
7˒Z�@�>��~5[s��qo���{.���׊'�p�7�馛�q���~q�8W��嶌�����K�C�t$����� a��K.��pP����%sD{W)�D�M���Tn�
a1`�uL��4�@O|��"MU�F	���UڎMg�yi;�!�O|�S3CJP����3�,������m���B����]�c7z�״�rꩧTR)	��6��f�8���3�qZ�T��w�����6h�2}J��w�=F�D������-�H��j�1ߋ�b�J���#��[m錏x�}@_���1`[�x�ue!������ԟ��K�)86��o�Ħl殘��g�,q��G	��xG�K��KS�D�L�ΈiW�A�̱뽣��`�4����7M�g���C���EB2yX�n���0N=�V/�F�6��{���Rخ��8d���\�H�1�k�Z2ߚn�G��^�	�VgJӅ���[�`�o��x*����f��&m�G�=.�G��ר	�vp�N;SrF��^���F!_Mփ�ML3qQ�5c��0F��[�,�����u7#��D{S�o|��邑�U 1��|#!ׇ���!")�O��'3�rv%A�^����=K�� ~�#��a�(	��K�ہ宫8�ViSF�����O���f���o���y����Nw���M8i����&�]�ȭ��T�_�6[^s7�8y#�+�.�����ݺg3
�>������f�U��r�>Ԍ�PW��Z�o�s7�ߗ�}��<Rm�X��G���*�T�Z��6�t��B@]�;߹�!��0Mm:��N���kh�bzٸ��I�i�s!��[�e���j1�][=�Sr��QK�?���i��M��S�4��Rӂ��<������~L��. ��v����2��{��{�����T��T	;��'p0�^�<��U+�����8�{1��M�����v�Y��G��%�몁�{ݽ�)��$��$�	�Q}�2�����YO%ym{R3.�|B��z�Ue��-��������;V���:�6�zV��$Sc�����J��EY��}Ǚ��J�iJ�Q�x��g�|g7�9��DW��Sdh����DDk��ţ��m���B��2"� F�J��j1v?�x���O6Sp�3�f�RM+ԏ�`lGH��7ٓ���e,��T]��6;��Oې��M&�R ���F����Mp��h~~�=�@1^4�����Ԑ�R�S��4�^S����~�����C͠uB׿�'!n1똃��!1�aoQ�a'��a�������T�-�v�Rt��z:��D��"�x���z�aWQ �1�Jv�����HTQR�c@�lg��j1殨�P<vv��ϏV���촽�-��:/m�6�`jj�p����ƅr�rQ�S1�vt:����e[�!w�n{Vr1ݦd��U��XVX�dzu�����U��:��0u��!;@�L��t���� �T�[��q]VW���R:��C<y�D���N�oT϶S}?��G�o耭�c�g'�΄�Ȭw�䚐�n!�M�X�9��<8��fm�����Ȋ$�����g��׈��d$�Hʎ�y�&�^�Ef��sKվ���UK��۷N��ɹ_�;��/�������F�.�����t�Z#@v˽w��n�w��ݾ߮�o��>P`Ȥ�?l5�h�`;%	Αn!!�����L�����9��n���<Ux�k��	�`���8F1�5����{�wj7�4��(EU4!~IJ�2Z��L�#1Kf���E4E�������U��Y�h�"����m�\��#Ozval�c똪�MmbsoB�:�k��(�79��E�r�X��w\��c�A$F�mҩ��v�V�L�cj:���-��[���d���t�����#�?�=���L��zf,���)#6b�r)^��WUʦ������|z��l��1�"����C�iU��� �*	W�	vc������TJ�i�/�����կ��و�����|eS�)���O�2�L��.a���=�G�.�a~��1��5=X ��66��L�H��gL�Յ2�=��oQK��t�)G�e���Sŏ	���DS��M${��{h~����5��T�Nl�Tjg��cI#E\�x��2E��{�6��(�s}�՘��l.��|J%�X�h�W`�7����S���()+M@>H�������������a � >ڔ�c� ��o��oT�vu�������?01��_�����'[rO�C@���s����eS��f��ۆrA�J�i���À��N�"Jl�ț6F�0����(Z�f���`Y=�����`�;�H��}b��x��l9������ֽO,��g�Oc-����A�,�hv����"l0�;��f��,��\��ǐ�hs�,8fEL�g�=c��Kʴ+�ǡ5��Z��H����]Ʀ�Fڞ���?l�jW�|�C��(&������f��g?���ѣG����x�h��zH��������=�i�N@�G�ҁ%���#	��n2h�@M J4<CH�G2�;$�A# �$5Cx�8yR�0U��v�c��9 ���1���z/�3��d��,lfÀjpS��#�&�	PO�
�̢�:7M|�\)R�vT�C��?Q2��"!5I�q���tĸ���n���M�f[;�}�u���I:.h��F�8Ǜ�c�.� M\w<,�ZO&�aKb��t E;�v�谐$�D�RP�� 2����Ӄ+�M'NF�5�����Ϫ�!%�����(ј"��g��&	�z���C��sm�u �vGA,<|���SmAl��9mC�I��p�xr��BA�Ĥ���j��_��Ƞ@$��>�[�1�`�G�TrO��y�^�i�k����.FJ~���)q1o2��퇴�s4�F5I{в�o\TgI�L�#�c���M�Y��pm�lW���}M�]ME}��F�F�h��&�t�z����-\ptԫ1.�/�؊6��4���Av����1��8�����;�<(S�ǈއ`|�rA���J�nw��܃�K��/��]�D[��6�e�zxi�m۽��ﭾ놙(A���X%`��3�`�4�!�5��C^��^v٧������\'�9}R>w����'(����B��ӐG`&"�L��x�w�^���}����\s�x�����۝�Zm�=���kգcە�n�sv�{ɁqA�FD��n��f���_��*�S��*���kl���N���m�u����6k�g�C7�w����7Vu��@}�[����b�����cܭ��Y���[ӰK"A��ƀכ`n��x��^R��̲mkm����w�����}���;�+?�S�᛼���}��/�U�|l���X���JT>9���
�VWr��J��o`��GK�n�:���=6)mU�9;:#���<-[[�����BِzX4��FD�"��5$%�(��k����I�3�� �Hc�m��τ�f)9:��3lѢc?)y��c����5JR|b�7D��O�E�z�o��@]�^���w�Y�u|Q_5�Ǟ���b�a�Q���X�w���)��r]�V�����6u����<��kw-"���=��CtlW��7�4��W~燋���}�F�.��+�#\���>N�:�����ҷqk��BFP �jN8������� ���Q)};���
=�V��KH�@���*�Ɖ-�y_��u��;�=��I+�Rvȁd�H�n���TOQ���r@lq��=M$������~����D�Z��cJ�P�Hg�Z>�O!��2�qM����������ܕ�b�b�9,.@5q��\X�2�O�C��eѡMudZǶ��XE�#�y0�nD�����Ї�z���-����Vln�� b�lȟ��3���TzS[�F���R������{�����I�_�vK>�b|����G*�u7cݶ�g��F�>�%e��	��������G��c�����T�a�+�Ds����(AJ*�ҷ�wtp�N_3)��\�{�Lj�n���%Sc����t�v�ǚ �?���w��2y�S�ߋ�UQ�p`B#!Cq㋦ɝ�c�@bՔd_Yf�4+�ND�q�� C���A�GɖIN9	=D�vC��tщ�>���-��IK"�5�J'�p��k׋��s��=�r��Wuz�#1����M��o��g� Yc�����ZI�H�r$�f�ݚ��_��b�
��}���Y�߽���:�.�2�ؾ�\)�@��q��Z��MK�Ƿ܂���U������Q��^_dt���"%f_kSd2��C)Q�aT1rt0Ё�=y/�,J�Q��R���rY6����T��B���=ՋVy'�'�0��L���^ԝ�B�^&*�E|/���&H�Ҡ>����	mm�\ӆR`�K��9_M:`��,�&'}jL'�aQDd�����E��R&�� � �ww�fN��Q݌�`4��:W㢼�,#���5!"{pf�Y�9ȟ���H�Q7,X
)^��+��0���w1O��%�A?����X�}q\�!�i]����ǗQ7�bfѡ-h{����r3��H�F!d�Fu�덅��Xm�J���������ë�M	Yb�=�>��?��j�jʈ��B%`&��ä��@g���$�x$l���5kס�9u�AN�S~#M�����D����L���r�Y\H$��¦�	�L���J�{�hc��qׂ<�d�/�n�a�x^{
�%�q!�<��H��&�s㍻�Nm_>ǌ@������"�@���Ȃ����y����]�\�.��?.���d�fΣ�n��=��J؞�M֙E����Q@��]�Y��c�$�=�21�<W�E����qV.���ndHN<�5Z�2+$�%���]�5,,�^T���7VG$!��"k��,���@T�6)<R)�"��|_�߇��p1�y����2~ם��VL�1OLOL�ܜvs[< i�	�kF6�H@��)6M���˘k,kLz�$� ݳ��z�4c����!s���ژ��k*����~��ݙ������؎���Q�H"�w��ݧҽ�q�e`x$�ڛvv����䭳&/k��Ԥ,��c66f��"�n�\�$bFA9��=s�.qA���I��`w�mtr����Hʱ�19��/(��GW*;���%���{���������$s������Ĕ�Q��>/zы��?�����ۿ��� �H#����F�9�a7�=7���k�(tT�p�X�z	<���B[������N�`O��c���?����J�سi�w����=�ګi�Q�lc^]}��yv�zm6؞Fy %cW�����i���x�ӧ�3Y%7OS���LK-�vc,Sγ�~��d���;�n���<�[�LsL["!C��ǮIp7�K\Xg�۲d�FC�O������͒�q������x~�g,����1���@by�_X<��ϭ�]��� ?��F=�m�1?��3����<�J����r0ؑ��@&r�[N%)lz����X��/��4���W~�W��h�H_7!箪��g�8��L��4�h����,�Mj�"�.���w=-$^���`_��MF?p�m�51�j%q�p�
5���D)~�ѵS�!>��OT��cǮ�Hv��g��Z]��=��#ӱ)�k��DB.�Ʒq��:+$3����zj?����l��1w��uw���Iuh����R̠���7F,�;wc��_�a}��6��<E�}<�Ņ��e��#)�PUN&�Q H�����'U8Wd��� ��(q���ܤ�:��.[|HLq̺C��pL`�c$����m%�&�g����7��Z��\�n����Ƣ��o��*�#�朎���,�E�m�J�q���]`bM�}[gL%<1c��!�f�~XVR�����Ѩ� �^�w��E%%�X��4�E��g�~  ?-IDAT�c|{*O�%oc�m��W�!���Y��,m��w������qa��h4_���`Ơ�N2a���؆)I��$��IeNd��D&�2	!�}��gz�R�G�V9������`���P����"\��mv;�=������v�����v|�B���{�P���\8��#N���M���q��J�q#��������:i�v�5m�H�q��Q����s��C��iVBM:�\��,��h[�'D��^r*Y��ȋ�[ϛ����&D�U�1�M?mڧ�9/��g�5�ĝ�1�v�7��V�
	$c}�<�$��<͸�h�85t������	G�6*UJ$�G:)�QʊR��Q���@1�$j߃|�~o}�[+'#;���$��gߍ�6
��I�ŉ`�͈<�(\�ٛ���8������Q�3��go}B������4�j>< ?~Ϣ�I�.H�f���m2������ �c�v�25-9:��Z�Z�g��ڤ�+�尬�.B�y�Yj%"�&o�6Mm�{s'���W0:�H�h��8'I���)!D)!:;��F��^?��?^<��(^����y�k��N�{��Lh7�����;��;�:�����S5G5Q8(���{ڦ�]��Nm��0��b��,�=�?#%Q?�f�i�b�7ܭL��Iy ��M��j��A��P�7F�Ԟ��E]TՋ�E�4��FU������-B'ѥ�͔�������ڳ7��?��(!s�3�LL:ߡ/�7~~��k����ʯ^Q�1+���B��{~ڞe�T�84��P���6m3����i8���ŵ��B	:c/�F_��Jh1G���j(p*=�Ϭb�!�׿��SB1e�N<�,����;&�ˢ�+Ҙ�B3���)���fa��f�-�q�"az�T�����*q�0$c�LӅ& ۞k��'��� Q���YH�c<�ҥ�n��\\=.�kK��p�o�e�0��T{2�׌Q�]iwsjvPk��x}R��f}��}��h���iS�&��sM��/�Q�im�;��yP;�;_�:c'�r��k1r!ڊ�hu��]��[���HL�{n��<�r���_�e�����T��h_s��+�ЕZ�hК0�I;��$np�p0��Ii����Hx�H�A��U9�b�ǅ'�o�t����v�IjѣO���#+���s8�E$�Hp1��Z�Ș�O�j����{�#�n>�'Z����[NL�U_�uo�(�8�o�pl9�flt�,��@C'�	�+���pR�EjS�5��@v'Z4�K ��4}(!K��:��8aD��nV:��<�.f|�6fMѡ�*����.��p�;�ȏR��Yr���k�g�l�$.7�'n$�Y�:�&�8)��q�r��)�����	��J�{��s�:�R�z��l��9%�o�i�8�tS_wsj�u��>��C|���2�_QC��yakM�����^L�����牎�6yYn��f�$U
_����fk$�׉�3E��R���!�(Ii
������g�%J�������+��
0Z ����'��l*S����ߨ��B��6Ш�����.�b���[�T1�	m��&T�}M�ܧ�)��x��Ƒ��F$Žܲ1�q�u�]��/�D��vj.�q�u���;����lçs�?j���q<g���‐4ixH���9�z��xhg�*ytRh���c0~T�@�I>RB^�r(حo�-��Lʪ�1�$j�w)�:qM@w�����a���$�J^c��I.J�}�u]�?���22f����������h���taK���A���`ڈ'�j����2���iF&�eq`RN	Ss���<��S?�S����}�Y�M/y�K�Pz���?ӄ��I�BRGZ�ꑉ8#�[tb���kԄA���\�g@�l��ta�^��y�{�t��Q�O�+dM���׼���bDF����nщ��a� �؞�!fH�-Ā��J�!�}��&�'����|��C�2��L�ݠ��P&	A�H���{�_<M4�)Ő.�t�Y�M'q�
�w�D.ǧ2x�m���<2�v���c!)�昗 �95n5���l�S�Y�<	��ѣG�$ώ׊��Lq�M�����ĎLڇ�LF�2��BR�[���!	jKn��nuuļ��2�)��lSب��f
̌���u�BR����V	u�f��^J�1������T�YיGʖ��`��7C�6󮡌��5�BR6���졦\pA�K��&"N�?o�F��)p�4nY�9�3222�	�}�d��O}�S�s�9g�#Ԙ&~6�t�9I|���/��
�K�s�21QFFFFhm�0T�#r@<r��D;rJ��0�{ڻ=�ìi:��"##cݰ��Mi�
sCxl�N�G�6��;m��)���Q.#0(�y�3222�I٬nF9�pȳ��I��ąT:�i)� JؚPx�d�t0�~FFF�:�U��I��"%��H�EN�&̲SKК,b~es,��M�iaj�O��<����]j%�Z�rЅu�E��-��x��u�m��L�^ư���!`I�D��@n�A]:)�(L���Y%�����>M	������jQ����~��{{�ym�7i4�梲-�EBIW�����`^���a���"fb���`�Е$0�z�h������c����ӗ���.��.�֧+�_�{��7��(��[ ���r�G��L��F+֊ǹ�^S�t�u�~��3�"n2�C�<I*&�o���̳�b���Z�s1�X`��N4��ҕ�d�y�����y�tQh2�e��/$_.�_v�e�|�Еz=�~�i�$>��*�9D2�;!�8�o������B���	l��&�yRe��zjSn:k�׏����D�7UIY2���FN
����qP�h��g���h�L<�Ň��7�Y�l�JU&���8wվ�������_,"V}�&�Ӄ�r�t��u�KR����g�����UB���`"C3�"��]�=SzFu��6�A'��1�llv׎�&~���#�B�)Z%���(�v-M�~&��u��_ J��� �-�UH\��)-�Ծo,2_�:J8�n_��?��Jȑ��v�6��=<+�ŕ0����p�HZ��Q-�E�wA�,��4��d��rc�I��f5�lS&���/w�y�i�Hm{1
�r��<��<�u��c�moOZ��Am��X<~��7�&:�b�aT��pU�t!�O6�������1��Hc{��s��y�SB�^�T ��H�H����(*:�C]��f�><��)��2����Y�N@8���b9�|��)�( ��ҿ6�(=v!)/Bzsh�h��IS��9΢���UtGDm�v澞��ڃc�����������ו#�bhcs����E���:���]ѕZ�@���>1o�������d�\��#�_��Xk%��e�bRG"R�K�&/�G��:�����
Ik�r܋E�{z����$>����_l�U-��ej��Nrߋ���BRv"��()!M��o4�]=rʕ�A'(_<FjȈ�������E��]�+�ؒh�0+7P�_���R�*I��n]q$��:V�=<:��4WD)y��K�K�?�6д�%�p�*���C4N�6~�E}"U	��9��XI>:5 �#J�qr(aQ�Y(�r��{D۱��y|�w����'�B��,������hۏ&��M&���K�U�/.�#��9��?c�h}'"N�����߫��&�E׷|�M�:!�M��q��T�>�e�$A�Z@D*!�5������pUڀ�׌�C-̲ESFZO�Kcɛ�cQM51̐�0��/�p�*�=��S�u�{/|���\��"U՛5��;��;�����U"u�t��UٚlÚ1D����Q�\�����`M�?3�D�2�M_7�c�a��y���|mDF4ediy�XH��O��x��.w)~�G~de�1��(}����*'�A%ɔ�����Hre���S��G����C��RBn�,WQ7������s���g�_�=WQ/˘��C���%f�E�x���2O��v8��sr�=�g�pc�p�X���Bə2"�@�� U�lW���D1z�P3l�q�b:�M6}�Oyi�Hj~'B�YR��w��ՔMH�چR4����o�a}����Qg8f�Dbn��>m涆�4>1�1��رc�@<r���yf��U8��A��aN|T�	Y�&��MΠ�hc��J��h��#�3b���I�߬C��*��C����ȣ�v��hb1$0��:���#I�����xEE�Ox��4����%��}�͠FB!SNH&�W����_��_��aEO	9>�����I��PRd��ݖ��	`��S�չg�0*��)�N6Y�1���M�~Glld)�OT�$��18���K/-^��O�ӫ�!n�A�yߤ�(!��feg�S�O���%�\R����o��*'�"���9%�u ,��T��k��$!���R3]���R-'Ν����r�}���xLCשN댭T���g�yf%1�����JBHAw��]+�4��@ۭ�Ѥr�{ܣ��=�'��aa�+I��Fs�:I����:��]N�CIbMvi��&Rr$�؇C���-b}����:�0uaL#�|��ѣA��E��k��s���n�� �7�=y�\*�Ʋ��I�y��_��q1w�I떆�}�'��(��󭬋�Ӵqǹ�R|?�_l��#�K�ɇT�$c&�7��$�YDJ�� �k��fzf�;#)�
�ޣ�t�f�����O�����[�tamB��և����}�p��-�"iD�@�ƱG��!b�hx>�G9(R��E����,��*�aD�t��27�cŉ�����S�
�[��&�.c�ز�#9�$�J��W?J�y�C4/x�x��ۢ��u2X�8��Le����{��^�
�
�U�SoS>O$,���Fa���:s<�2��m���;�kߦn���  8.�/ڑߋ[콗1���k���m����G?hwn�V�1%��7��Ź���6�T�o�+�f�LF?hu��A�q�ёd�t.�H���禶���w�cq��߽�|�o���)�]���J">$h���\ ���O�.��x�&|�9
2��@�0V�1��cP�%"��8 ��w�s��~�r�i�D��*��Z�I=8 �g#�(#��X�}���`��@�����/nH�C���:l,$�&{粘u��b�1yL*�@2�������Nw�Ӕ|!jl�D}0	�cpB�LLb���G	�8� 7I�g'[J��.�y�c�6d��̴̘�v���	]��A��&�Tbv*��x�3*����ԉ�D�0k}��_޳ﰴ�Y�����_x�W��7}�7��=�3%d	�.��������w�_�uJ5���lG��$�tDT'�|���$r��W\Q�C?�iO+��ۿ���Q�v'�Ă$�������⋫����q��б�ZA����L��_�B�'=�8��F;#�cT{���j1T-�[�[*�=(/䄚������8y�S�Z�O�2�&枠.8��cU0��I�J�('(�w�wW}H}u��׾6�O��.��ñ3��<���%���E�ډ%���1��������x�#*b�.UVm��u�nw�[��?�"�~��ӄ���p�!��������6Brz�s�S-jLp�)�y��Y��K;I�H_H���6����CZ31�c��;9)3m�/$f:C�|&1��aבv�a�����~��p�S��2�C2J�����S]��J��H=;�G�6��t���bx0��=Z��E/*�w��M��a2��x:|��M�R*�Y�<<u]�ՠf2~�K_*~�g������J%���?_��m�	 �yC�g�\ԫ�F���X��꫋�=�y����3����:�]�x߃<�a(a�&<�\���g��~自zП����x��+�M��\�I���F&ߕ�����N��;��r����c?�c�}�{��������y�{*���M+7�EJ~�CRٕ/�����2GR�C�.XV�p�ƕW^Y�T=���+�{�׎�D3iJ�����a"��e���he��N����ɀ<O/�V=Y��D,HhC������g?���}��%_�����\���-1�l�y��DR��j��4�hH�{�êh��[������	dV.$9$&$"�HL�ư���2�l�拈H&m	�:��?������W�RR�C��<&Ƅwۼ�c�x=����r�{߻�!�����m����3��u�}�S�\8lb�\�!N=4��؇)#�g����ƅG'wt��A6E[��(�g�\ϐ-�� &�'����>���Q��>���+&�7�o�	���}9nW���6L��M�4NT�OT]�����7�}���;m��$���~Im�1��*��8���X��O�t�<�Ҝ�E�@k��Ml/Ǳu��;,\��
-*f�KI�r�@�����9B�M�50Q��ɑ���́T
NM�
R�kV�}F7�))w��h��y��)�	�`�Q�w���l8��H��\�L�\�1�Wix���<�)�w~�wVڇ�nR�׌�b|�a�qq�9�T`�}ڍ��e 	��Tf��@�NK47�D�D[�:��2�s�]�(-��) �����,*7�H|qz���%�����!J1M���ԧ*[+m�b�T�Т��T:rB�X��/�3�_�zֳ��%��n���
�;�by�|D[ %��5��F�*c}лM9��c%�(φp`�p:�n�Y��z��~�C:��+���-�#�Mߘ*����=�A���h�E� ��c)���'b�Һ�o��o�L*�pPI~(�%�C�,Y���BU5���������h&gLiL��ݩ]�I�;l��/��&O2��"N�e��>�F�m=:&!d�B����ߍA�$��F�{nwGB�~Q3�&�6H�~����=V")G�����~����7���G?��Ņ^Xm!�"���1� N�N�1��tax�Yg�5���M�q��g���"���M�ї���&�����%e�:�,���������4ӌ��V���%b �[��
���c�X=�� a������?����̤4V3&M���Y,¬����%c�7F5~��ʹIR]%iͫc���$B:#�j{���VEZ�f��¸����2κ&�H������$fC�<%�P$#���$���ꆍ�e/{Y�7��:����å��<g�Xb/���.L:����WT���C�s����D^�B̀ҿ����D��"4i:�Iz���7i����AɀĄ��w��"�����lʔGɈ�$e��G>R�$���~�t(�8pSG��0��a!���
�{���Dc�b�`<���h�!/U{#���ԩM?��7}'���ǲDg��N\���2��]��O���n���O���f�����q��/^߅yBN��z��5�9�?cٱlAZƩ�6�o��o�&�y `�8�Pc� �)`Ou0���-��>CB������(�&��mZ���t�Y�X����֚�&[uF�XYB�y��׽�ڹ��?��U�7UW�6��c�x�c[m&xի^U��d��a3�C��B����864�W��e��*�,'^��:`VY�n�u��:c%����"�~�7sq�e���[�U�{ق��`zI	��9����.�Ȝ�:?�ȍ�h{�Q�XD>�>�g%�O��hKMM �T�����g�5]Xbb��F&�>���#"v*vdL������.^��T۰���g����ZEa�&�R&�۱�7���y���\&��u鄎6d�3t4�W����$�U�i�XWS�"�ɺ�_Ƃ���U��e7��5)(�qs��e"5̳���D�3?�3�9�'!6e>Ä�)C@�������J	9.0�ߴ�3�Cu]	�)$R�d������VfS��s�\t�R/�@�����o~�_��_+��GV$�T�t}�TN�̛��#s��u���¬�'�Q.<�V�yQ�3n���@�n�l�æ��7���}1Hg��q��<����׋���߭�0c�#i#Yc�~��X���wnT�H#0�y��RTL�K\GS�,��i�f�u2;����n/_'��|ች��l,2�HR����A�|�'EFbf{��������������q��I��������J'<l��	 暈����4�U�Q�E-�~tg������E��^M�{ɧ��D��nY-O�v��Ǿ`�2~u*36=u����x�È>�%񧾌xBM��yQT}���3cōg��3M�!��Aw���!	E���EL�γ�$E:�t+����Lr�'��ْ=�w��}���`��^C%�5PS����1Mƍ[G�*�ܤ����G�i|H

�/����������&b��b��ma_����1�'47���Ϲ��V����J�J~q���
��Q�r�|IHG��	^�s�4y�0����$K&jr�ZD:x�Х>1�)'aEi*��R	0��E�҉��7It}����F��&����m;X?I<Jb��Y�?s�>�����&2�:�(�4-�Q��}5�!b%�;�`�+��>���!����s�>��'|<�'�6C��n<��пT���O��R�ϲ3I��#��.>1�~:)CH��{��~J�Ji��&f0�	�S;�,��/4��".�qA�u�{��֫A{�2�x��1�LF�1+ɧ��as��}n}V]�t<��*�D�Q��UH�P8�¡gnf��n@$jm����l"�Âu��U� sb̺���B����B���©fO8�d�j{�,��g �G4���#�%4�j}"]p"�̒�W����e���Ѡ�)��}��=��(��}y":l�{�cz%6e;�FLNH����L8�c�
	��d�{�\m��ؕ��Tvf^�!�2�2�f!:Y�]ωL=���,MΓ(u 't�"�4=y�����cJ��~�T�J�������@��.��]tR�aK�
sFSa�ď����W���Jw��w�,�k��������
W����S��x����?��U���/����'?YhRt��í�4*��IN�����x��Xdr�������_>MR�ZRq��	2Ϯ�7f�M��;�Aj����(G3Hm�M����BsD*!˕J��~1�u4�4y��t�j!J��~l�T��-��iݘ.�q�{T�.�HY��ұAlP�g�>,�$���AӅ�ܓ���|����Ozq饗V��*x�رJEa�$�=���>��*[��3��o��o�P:�BIl�GƉ�n<p��f$Ij��˦}9jG1�$��pi��*7��Ԫ�1�
����h��Ak��{΁���*D�����Ӥ�x�B�m��Rö-�vղm��(�K�J�\b"VbSv�;��@RV=!����GC2��؆݊� �q1[����-.��iȜ� ~�!qM?�ª�:7�����^g?���(�v�4-��Q���~7��"�7&z�;L,����:J�m뗖�IL%Iʥ"�Kܝ�ob��c,��yOK�����dۅ)���>QJ�p>���YN�Äڲ<�L9����T 鸰��m?J�QPL�h�Z%VF�6��3�:��8c��;�/X�������:L�~��+bv�bG�3���z�Y�e�淩��	���羪�)��{�2��>�ދ��1]�l3׉�5=�,%�2�u�-�N�p�(�up����DI�Ѧ_�WTߋ��4�C43)ܡ�7�05��I���q��@�T ڗ������_مȗ�9�l��ڐ0Y`[�\�Y"�ԣ�H���CF�}YUz�$�l����&R�6�Yv�Yej�~/�ѩ���A�/�'�U�V���߄��c$�h�����tf�5���ѩ��!ڑ��l�1�"�6����hzz'eӁ�jFCy��?��?UN?�xxS��L���#��|����,���ѣ��N��Z'˺��R��(�3��y8�5W�(�Y:%�y$%8�Pu2����m+E���:%.%0�qcȬ8�e���N��jZ�ʼM�{�k?��c�2Hc�%�h��}	���6I� �^�蝔c�&���O$"_��E
fЦ�3�	H�{�ê�ؠƑ�]��J6R�Ҩ��a����kJ����=g��2剓Ή5�e�7M��R�*}��wQ�TRg���Ƨ��M��"��B�@���m�p�s(��lC��Muh�c��g�3`n蝔w2�M)S���ig_�K6��n����6��tڂ6l`p~	+�+���GH��{]I�l�U/��5�+��Ҵ�$�Fj�ep|r?Lr颳RnBj��[�㽆()FD��l�լ�ұ^q��ud�����JH� :��cA�������)Eh���X��h�v�����U]w�61ɐv�-�@����q�tt�t9����}�'�"�e$�Yr4W�uZ���$�X?�������ٷ�$�J�1A��?D{j���[�H�MB���l� �?��0�;)�pF�������?��xv'O��u	�$D�!�3�����!nA�} J�M�߉�~�����uy�W���j�H`�8�I���@ݢ��^k����͊D����I	DGe$߈8�b��1=Ksh�;�[]��!��y]HU����4��kĸV`�rTa�$2��б��7���Y�ש9a'�����r֔�����wCЬ_SY�ĉ_����J�m�%e	YGv4���k+�G;i$��� [C'��Ti�]|=K:���UckVǯJ�����U�[��
�&c�t�h�}P�*��Ȋ���ޑ�g-N��,�c�
=_qpᴽ���Q����:&����zd�[��YQB��۪�"�g�"�d����a����m-����&������T7�HZ]޳�Qnʆ˷���d/�X�޺ϟ1b)��A�I�1R	�����H*] .Q��^�pЅ�)4�E蠄���K�m2����{49�"9ļ�dGn�L���V:�����m�����+H�}�
�D�X�L<���x��wPD���H��~�E�$F����b���TF��V��8��[�VҾq�A��n���ϔ�b�p���>:���z*)�sXG���.M3"J�iv�&te>q!�=�	3q��~".RMW*�s�o��<<l�;���;j��t]�$�4g�1A�A��ERl��栛sb��vrǤ��A:�#/�"�6bb�7����&�TZ�R}�y8�QnHa��d��u�W^W>ߺ�;��Ef���u1yG'�g��N�n�uP��2m��"I6MP6�t��'̽��l�q�O_�~�s��昃�]����qB�	�jî~�)8J�濈�ڢ�3�v�{YO�V�g��a�g<G�I�����m���Sv��v�l�.�����r�Z�S��=���<��+r�s��?-Q�YuQx��|�g��5�~�wˁ�����]r�R�^�^|�wC�f�'ҺX�6�Ni����{���͒@XO-��̷/?�qF�����.��=��P��!���2��=:��u�y���}���Rj4�p�K��{]H�M���|�T�4}��ֆp�|U�E�wޞ{5���hk�}$g���A2�:�����וｭ|����X������ɼD��d�;�������7��pC�<�l��<Ky�yRb��yͣ����yP~��>�����4�ݲ�s�sy�)���ߘ����o������{�ۉߏ����/�i�Ӷ^���k��`�;v�Ne'?�|��π�8����tR�����%.vY��:�x�s�[����>��W�hn��Lr�B��
m�%�z�N!-$dN�y��_�Z9H��AA](�ݡJ_��fѮF�����>�Ƭ�����|�_���?���k����&��˗*�7�WJ:g̬�f��*=߇�����Ri�/	2�0$�L�ߦjnސ���#K���%��O�f�ͬ�mC�/�n4���̄��Ȥ�f����D9iOW�eˮɃ���@���r��a��bɱ-��ܦ����<��9F����W���l���g���,>mC=���.q��XKdR^O��|\\N��!��2!=�]"ZV�� c��	�����+��;ܩ|�w�| xF�`�J����C�����9����Y��RR��_�rbF�|�ox�g=e4"����p_/'������t3�1��)z �"Ҋ�<���(��@&\�s<��>U��������������w��'��ǔ����3էI���1Ⴁdۆ��$$w:���e�S+HC��_ӑi6��X���J�����{+E&��ś��O�$�&/�Z���]\m6` �����}LA��T�tQ��c�C�3��'�2_,	�#������������;���f�aQ��'�x����ڄ�i��-�'��zfi[5��N����.�~��淓��o*2�������tI4�\�<�|>͘W�LLm�� q+e)q�~I7����r⿳��������e�	Ic�@����	�I���+�U�d};�?ˡ}�z�I���.�EM�Z�+��a�vU��~:0����������=mUz�)�)2)�1��)�xl�ث�kC�κyRiBrW����|���3�/��7Hk�.��墶�?�|�[>�.�/w'�|Fdm�E1�sO���-�1%:ڃz")Kz�vz,�S�jq���k�=�N��1<�O�o�|NᏔ��_y߇�e;#��h�a
�����������.����p����%~jB��F�{��r~OQ�2T>��|ܧ|�k��Ix�|ܡ�.j��U���;y�B�V�J�A=O'�t$k�%D�e�|w�.?\�~|�e��X��ޑIy�QN��	���&�G<$�����J��� �5��QX�2�3��=�ǃ�����qvqx��_-�--�*�ʯ)v�ފt�a�ߛ�m ѳ��(��&k}����шL��O���)'������n����6��4n�< �/�u �㽼.����jq�|Q��������U�����}��N�$oH�vEGX��9c�Ȥ��@��x�xT��	�ă���z�'!w�)�������������~�U��|��|\S�{U�ᐼ�����%(����"w�������O�p���|�R��hI,��ݵ�{!�_|�)�����1G��3�X:3]��yn�)rǭ9��?~����uaw%!_R�D�?S>>^��7��G�C�$�SR.��"c-�Iy('`���X>d\^Զ�>����x1��!��>�M��^S�JU�/j�����2٩w ��>�_������T���p�1-з)dRpu�sX	�wq|��k����b���$�9��W'#��"��P�q�]ǥ6)�� -�B�e�]���u��A��N��82)� %�Vu����-�$����z���ĉCي�9�rB���Ȥ<L$����Ö�!�k�������ڡlE'g�e�!2)� ����]��̎�R�c']_����ѣC�9O;������B&����D_�a�5�$�[a�Hz!�,)�/2)�f$0_�%��y&#���G���ml�]���_v*���␱��G���M��%�@�dm�%C����9c�L�#��g�I���Iy6I�ʞ�=�E'#�$dRn���锔�'1��q�G_��"��8@$A���1�4s7nnn^����G��!�dR�؃L�� [�GgS��*��Ͽ�cǗ
R��C�6�9w�m��ǁ�%�b6e@ZMv,vM�CAj�7��/2)�;]۔$i�q���;Im`(۽3�L��@��ր$-v+�꼼�����f��C鿌%�Iy@��T�)����<I��n��>R���2�D&�q Iy�۬�|m�)OЇ&�IyM�Iy�`�Jʷ�R��{��`Hyr�bFF�L�#A��pF� ��׺�������/vr���"��8@�E��Au}���݊��r�upr�DgD������G ������k�o��p�ĉ�I������;@&�5E&��k�iu�r���~83�&�5E&���T���:��{��`�y���d���"��x0�IX�'�ܾ�k��W�y>���"���5)%�E19@���1C"e����q�Ȥ<��^s�5]��`$�~��u��|0������<�rF�L���F�1�:�R��qWC1杒�ư�3K ��xЩ����=$���u����֤~]Kʃ�_�rȤ< ՎYRf�X�����3$�L�rȤ<tN�Ű}�]o#:'�l�X_dRl�z�]q����x㍣u�M��њg2�C&�q`c{{{0$�� �!�רm��!��x0$��c�[v�e�A&�Yڤ31琸�)2)gǏ��;%�!E�L"%:%�}��Ȥ�1C��p�`�Az�v��dRΘ��Lj���L�;E�Y���!�r�,)�s�Ő0!�NI4۔���ǁ�'��&5R�hI� ���2�@&�FL��\RX�v677��"�B&呠�h�!�/��%�k:K ��x�5ifR��6������o�Ȥ<�]��C�_�)gTȤ<t2�1��:�N(2ie�����ђr�Ɏ���"��80v�Ũ�xw���Iy�csŐ����ТK�Ƙ�UF�L��@�!�D�}`���XSdR�hG0���%�l����ǁ�O��������3!gDdRΘ���蚸6�]2��d2)�]�N(�OCZt�0�d�)2)�9���&���"�rF#�����Em0�rO;3���ǁν�c�$76Ʊc1�մ���G&�� ��%�1~G������ǁQoCc��9�s�ر"#dR�n�u��YRΨ�Iy<�$3i�^��h�L��@!qCKh3v��y&c9dRF;	'ө�a`��y���Ȥ��Ȥ<���FR>��ӷo��Ʊ�L6_dTȤ<��|ѹ$�1��K�߀�Ќ"��8��3�T�]���Z�;%����2�@&�q`��m�����EgԤ<�E5c	dRvFNZ��1������XSdR��c&-�vs1^��Q��2)� 8����1�2R�-Ÿ�%�
��G����NIk`q��۔7�2�uv�����G�l�C��v�����v�um���t�!��x0�8ޱo��T�͒��"��xеd;$Iy�螴�D�ԭS�6���"�rF#7�ѵ:>��Q�S��`��X_dR:��677EZ%�vJZ��i���5���!�r�,��:�$f��|����E&�F�]�/��\w�u�|�1E&�Fl[s现b@; '������Ȥ�ш�����V�C�EQC�A�I9�B&�Fl�;���3}h�|��Ȥ<t�iuJ2CZt&�L�2)g4bgx�}Ǽ��m�SdRFMZ]c`۬7������佦Ȥ�ш�m� ]o�T�2�f�L��A�����S�lSΈȤ�1�!�b䎾>�3�Ԥ-�Iy$�z�����ǜ�t-)gR^SdR	��l�H'`��
�1rI�(�|�Ԛ"��H��qIt�u�!-:-�k�v0��X��ǃNO{����].]/:C:�u�sʐ�/c	dR	�I�))L����Ԯ�= ��{H���2)�夾��K�|�tI�;_�@��/2)gTȤ<��|��KiR�ұ&�=$I�ȑ#�ǎ봽7���-2)����7��Uhՠ$�dNtx���ٔi�N�O��h�L�#AIZ��J~j�ؤF�디�$)����uy��K ��HPNj$��H�֤����$w6����TR.�摵E&�`{{�rgD3�8��I�l�!�m=�E"��Iy$(I����!б�MtZ���y}�Iy$ ����c'��P.bc�ʖ��[SdR	JBfvE48DZH}]�̐$��ۺ�<����F����Ӻ$ҁ��FY�����I��,�_$�T��%�Iy$(%��:�#I�<��[��L^�!�}ں�|�C�_���ф���\�4�T(5�!�}��i4H���3V�!̌�'_g�5�I��8��$�u�ŐB�2���f�>1!���IyH6�S��6�T��S�[&ь
��G�R��K�t��.wJ׎��qzf��+�7R����Y o��e���d,��� �[�S�    IEND�B`�PK
     B"BY<��G�4  �4  /   images/e4b09d94-725a-4fc8-8861-adc4f6b1a3b4.png�PNG

   IHDR   d   �   �{#   	pHYs  �  ��+  4�IDATx��}y�&Wu�U��u��^��ۦ�`l�݆�ŁL�0�B� �H���Q%�3�(�A���H�(3�$8	؀�M��������^��{���-Uw���{�n�WU_�ׯ�!�O���}Uu�:���{o�j�]]M�>�"M���g���&.=2~U�ꎰ�'�Zk��Z�&e�Pٚ��f��a���A+�	bs]��x@�HE�r�
4�՘'��������wm)S�=s��q�	��:@%�fE�'�B1����;q���v�H�xJ�� PQ7�ヅ�}�y��wGOѢ)��{g�7^wA-<�&��g���������~����Z	ƷF����o���Q���L?��+Ma�t������-����="`0P�M�aʆ���5U�H���z����H
ڦ�V`�M�v�_A��#S1�����p�3�|�j��gU���}�hm��&�k/��?��'�~���=�k�I/��`\��Eͫ�V� �{l��wX�CN1�A&Z4s�,�JH�o  4m-����'[�+�  \d�jO��� �-����0��IZ>�h��6j��uf&h�4 �����k��ժa>!Ts��h|��k�|��.��g�h?������v�H��"�7�4}���=������g�6HAG�d��Urh��@��r�R����o�Ő0:������\��{���PW����w��%���Qo���Ί �tRϠ�� "����w�뽗}����BS����}q�q矼c}�F=��4���BD�m��As�2���Z���i5���Aj�&��Hy��Y)g~eEM�,myT[L��� ��X9�r�QXq����nY[]�gx�i��*�ڪ"�:C�,(�������������ZY\&�����]F�0��l_�� �ж�:bD���o��TV� ��";Rb"���N��~Z]o9Z�}g#A��B����bJډ���nax��m�K�y�J��Q�P�
[���x�J	�����YE�3�r�mK�hZ�)���L���?�"�-r$}a;�7K�4�Z�\H��W��ZOE1�0:X2�^�S�b�0
L�l]j}@jÙ�Y�al[d˲��;��o��UZ҉1T��F��FsP3P)w��j�YE[)ѓ��AXR��bM��1�6�4��JG佻��o[�3��!c
Pg�$�<K� 1�@�Vg�({e��\~� |r�&j6�Y� �Q16�IƅZ���TFQ>�ڄ�E��a���q�:^ D�hb��X�������2��X��:3�p�ԍ>�ܽ��1Ѥ�1����tk�3��G�X���N|�����E���a��-��L�C�ˮ��6J�WSd�1iE���E��QW� ��mLh���9���f �v�$�Z�L+ׁ�=1sM��J�&�=��Ǉ�'rWT�\�������>E����U�>A�ڧ��� n����j ����-�V�ޯ�@P�NT�!�*��1���?��ğpqc�Fi ���(R��R!�-�\��E��h�G�'z�Ҧ�&[mYw���<���sl10�]�ϣbjt4�m�Frs2
���LK',Q<����8u�N�ʀ�jyn���ǢH���ƷL�h�ҩ�Ӗͦ���׶��:�L���ީ�X4�sh�D���0�w�41�Ʌ����W`�^.;������d�S{fҸL�WNB-��O.Rn���jM+�C�7u���fj���E� �WZݤGP�lpφCw,`Α�,X�T� �2�Wg�M8����r���)�E�<��MOr5�mJ�����΀"J\�,�G�	��g򠔢���%��#����u�Cԙ��4�[o���^]�s0u������Z�p�pV�a����Y(	z
�����6t�5+eE��/�ܭ��J���Zy�n��?$#t��Ubd�Ӵ�iS�	�\�v�BQc�I��F�%j�ܳ�@��Ǌ��k��i��V����øGn�l��^�A:j({�j+� pw� ӰS�2>f��D&Z�I5�����ʢ%2VXg�$�MON(�<�����ھ�&7Og\k�����ODu�r=�u���]��*gUa�Tqik1Q˛uH<p{e��v&Ne��>*���kߥr�dY�L�u��zGu\s(��ӷ���,��R�yxz��G�$@fgs�/�t�nh�.�ğ�h�������8�b-����!r:����gx併�o\w�ul�A^�ĊJ_D�����7R�K$��}u:37�������D�����1���� p��'���V��^����_�.�4�p��g��H�W�`0�(����j��67a6��J9� ��<�}����ͽ�W����:�Z��ōr��	��RkQe��T%5Ew���."m�����׮����sV�c� d$� �Ĉ�86x�����`��0Ty���CY��>�R8����᎛��UR�gF*��5į,�]��+��G��`y)H�����lFC�Ψ�!�� ��%<�c�u�_HH�,Ԡ�h4��� ��v��*��V%r׺���T��G͛�.���Ze%��\UeU�%{9KV'kѷIn�h�UZYB,��1G�E{毕A�-�XM�j68�~�N�,;x����/Q�عJ%}*jn��|S<(���#Q�I��ݶ�q���h�5ErR�5u�L�:Mi���6�[C����כ_�h��� Y[ӹ=�f=�V!��T�(�}�ƻ=v�0��+#3l��2���������nGg�ң���Jjsjh�[���[Z;�9�BIwy�N<b����*�PE[.�� ^�oVk����St������;xϱ��]��T3t�'V#`Df0�<�з��f#�ymM�i�Xq�F�!�hܴ�z�G�A9ŕ�8��p�B��{�}#�Kn��/HB��p8�uF�H����[*[q�{p� �a� q�0Hor7m�Ͱ+��
m'%3��pS�.d���MT��PL�>7�T�3�+�vE�1�A�*Q���ܬ�&JF��_T2͓��'�h��S�n%$S��xZqoC.U&N�^j�9;��N��N��:fPOݳߕJ�`�s���Vj'��Zy�Wɲ)�]����\��BO��Dns~GBt��O���j���$i1hѱ ᬼ_dWS�I��ڢ�	�ɍ@�)�yr�ǅB7�3RG^��L�*�#B���(!�;��i���큛U�0Lڮ����!\-�dێ7X)��o^��ɛ�$k����eۓN'#G@��w#��ί���ۤ�Dr�u�'�������Ad����F� �r�6�݆AR��"Ô��SH`E�2ڢ��T]���� h�YCg{%\a#����7݄�߈��֍禂����<��Z��_I�W`O�n�����ҋiqb3E�.��f�Ӳ�!��8kЖKf)�"喻�gv�#���;BXޘ�[�\`Gj�~���øb�~J�Yaә��f�IC9�X��bj��E�ZC,3Hfv�4��r�0��l�����	�]�_~��P��az��:x� �q�bԗ��;v�M7�L��̨{rz���Mƅ�ҫʉ��f<�IRL�ٕ�X�n���ł�,�b�ΰ9�NVMeV�h�w������k�R�a�g�e�J�n����k"|������]x���ٹ����:~�8��G?�_|��%�1^���[��S��\r�e{����ǂJI2Ӕ`,�KtB�VKp��O��X��U&�7g��ϸ:Ņ}�n�g�%��\��W&/���0 #��'�-���{�(�`��y�fz�;�A?����"�A �.��"z����#�v�[����9K/?�L�<��Ų�g��&F�#!�uZ]R�;Nʍ��;8�XZ�j6���o�	�{N�8A�����?�)�v�m,��x≌��h���7��_|����w��Z��;ۙ�xU�s|���B����л��.��;n��f�)����<I� ��+����l��T��;����M��P���o}+���t��Q�ꪫ�?��0A��1����:���=�;��
Q��	=�CV�	d%r���_Me��_TQ�j�L��ה�<�;Xi���_O��ַX=�,�k������x���Y�C5f��7I�Ta��{u��K;��^�;t��x��nJ���/�k�.V�J���477�% b
h����F�	ȚsU
.�!�k�j
����p�Z��gA4���p�p��:��E��N�!Zc=N��HJ*���X�'"���̧�d���ß*���t:L���j6S��%�/�&�A5X y@�`e��R=^���ak��=�r/Rf� $1д4o��Gv�߹ڼI��OZ���A��l�O+��Sl�:m�g�e<u�v�r�笜Z!fI��ƦǨ1�t�w*px��~L'_~�+�\���'��`w�p0Jb�$�$�ࡥ�%�΅^�A7�p��Qj"� �S��h����a��!��EZ8t��?q��8�y�����~�Kٜ���xdΐ9t\�d�1�'f3!
qA��#'�;�L�� �k��uh�m�QQk�,�v���	L���W�{��<2>����.//S���o�kC�����
m۶��q��x���qx���#T�a��.d�`d�<3�B��*'��Fn9���8���\L�j �]es!���8�#킅A�"JW/����F4�0ڥ��T���I%�yY�,,��}��f�sF��A8-�}�k�СC�Џ��n���'M�L��Q�H�W��{�U|���r!�'���m��A�D�6$��颖�z����ʾ��駟�F C����pZn��z�P�t�7�*'��I��){���5x������u�Eb}I�Ʉ0.꛰[*>��Vr� ��ss�>p�@�����>�(��pZ�����3���]C��[���ƌ��)~��C*3��
,���ZUy*XRy����
���\�>k�Ad��}qp�=��O��g�e@5����{�X��h/b.�T�C��s�����X?�F�hcS�Fm�v�����]���kA�g����0ڠC�
Yꁖ��(%���,��}����Z�l��]g-��廾��ļ��7�m�ݞCx��J�?dgP0���|���?�E�����~z衇X��"���?�0=���t��W��B�;m�x��F`�/�\�%G,G��Ж�N�d�dY�v/�M,�(�5��.Gh�wlz�KH,�V�.I�G��]��iv�&6���P6�(��7ӝb�6�$*c[g,�YOӇ�㴸�d�����W�g����'����5�:q�$=���5�y��u4{�k)n52kKA��̒Gc�z�l%�ɮ�k�}|�E+��5ӟ�T��)�;f�R�&�]����y;�5��_)�2�O�]S�����w�I��Reۋ`�n�4�����i�>�Hia��\� N�=���� ��~c�W��e\�~o8W��=�HK@��D2�2��NE ��~nn�ZF
MH��
*��C�)��ˁ��t�\f���䇩̸1QqW���D&kH�
�*z�/��s~D��wS|mV�'��Z�u�gj��JV ��?����h����;eb/1�K�R��,f����{���u$�OTbfA�E�Ŭzz0��NQ��  ٙ�`��:a��l��-H1**Wz��?:z��z�Z���D�[,��k�۸�P!1�N֨䎕z侐ȑ��.3[׵ꫬj	b�я�k�Okr�K����x����]Svq�Y}�=�մ�ڼ�=Q��3gg�(��R���݂Љ��� ,����f�o��\���3��.������v�wd�=�mŒ�1���O����ˊѡ-R��&O�6Ϟ:z�VN,!��-�i��as|5��`J�� �`��� �8��6G�5����5�ͫ*))�]�or�~K��u��e��8h�*0E��S%�*��]�*~��n`&�����V(Ri8�@�">��VJ�J�@��hI�,��qm�H��p��))V�Gn�΅/����-Ȯ��Q-'�z+��l�E� ���bN�t�eq���Ҝ�R�*;hI��Ujb	�tߟ��^v}H^d.wJ�V*8ð�f/��P�@q`q�FP~O�#lL�Hً�
�f�Y��
Z�wM�X+��hم)�?gHlU������:����%#���.ri���#��<^
{*NPc�E��#��ն�rvl;Ad��y�V�M�hH�O�V�N�7@pm�c�0>�Ԙ[c�*gٌ�nMK�X`f��Z�ޓ	s-C楫*v&u�աa������l6� i�b�8N�3}�$F�r�ʑ���T�7���.&_��W޵�˲��,~F?_�v��.�g�&k��� �!��9p�Lm��̽:�qN�[;#�^��CI���L�ڤ�	�aa	/X�w���)��dN���,�o�P���ew#���; ���v���&�;e�_���1�'I�Ϸ2�킖�y��p��J��	
�/�b����̹'�T�y�s����y�v�|,�z�6d��J��zCW"���8��R	5	��(�͈�D9�"Ʌ`�*������f����I�����>\�s��"@�$��@��wOPD�mr}b ¬�E�cC�پ^�C� �DUC^|�4@���+)�b^��#�[X��
=�a�y|�M�n�(�rI6@-Et��1�ݾ�-�8$2��gg
������W����|��u%A�ə)�>�u7��'N�±�6��u
�On���Lz:��r
��W�S�K�q7�L;����W�sk�����Sa� 0N�V��nntO-��Я������S+�=�	��HL��E�ܱ9��z����Vz�(���)n ���
�m��4դZ	@��K���%)q�X�l���q���,c��w�k���Y.�00��Z��ľ9n�B���Jx>VOd�N� *#�����[y=�)�d��$���'M�&�Ƿ+Mi�^��}�� ��)K���NWoMe���z�b���Y7/v톳JF�*�:�{�"�|�gj\HBƪ0�tm�|@�mFW�����ʱ��4$�Y5��Ȫ圤�Zʿ}z=�f岢��b�-����d/��sԮ�M���1�0���dh���?��3�YS6�q���փ�`��U%��Am���N�ƍ�2�H��	4�MM��$��[.�߰�p֔D��U���M�|B��J�ûb$$��Lv	2;:S��R�)�xqr�4-�@�>��L$�%s2�Ƅ��)c�����
@	$�c�&�<~� hj��l����g��B�$�ew�!^i;}Ѷ�yl�J�
#8��잵3��D����lp��43��#������R�yKs��}�|�5��@~�=�O7����U#���~(;�q����>݈�`�>X��Q�Ա��%��,R�Q��IC[�<v	������nM�-�{��
����rY�%-_@YA�o+���"�C�Z9T.�I6qԼҋ|�|�xz�y���l´�y���x���UW$����EU��c:wS��՟�&�ǹ��[B��N�Z�j��u��C��`�[��[�^=B&� OO]G/��ڨ��$_��zO�IFl��G��be:|M��~�uU��y'��Q��Cᐆ�H��������܍������������_DQ�W2t�t>{=c��̭ӄQ�^��̷m+��\�.���g�����A�󴼴L3� ��JX;�
E�`��o�&s��Ç������~����^��y�Aa̤�
E�o�>��7��;�a�]��K�_�B�+vQ��(͹ڭ_���ӱ��hk�A�:Řu?{�Y��W4Fn�����:����f�Y�,5{�g/���ǁ�/-sm�S�BZ��Pv?���$��!� O�Bd�'��y���G۷o�[�v���F��K�Z7����k+P��m��S4�-Q;�.<*�$�}7�e�����+��ҀV&w�տ�?h�뉒���^6r���qf�Θ8���݋K_n��!z��LMU?x���e��~;�d-+TӅ%y���M��P��S�AZn�������!���x��@��wY��|v�J�%�/���VqҴNf���	~iOOF��)(�����g��:��>�)�z[��#��{��^z���;�d7E�zHMݥ%Z����i��Nzve��p�\P~�X9,��\S�8$��[!�rY��^�<H�P��3}��q�"��Y%v��d�n1r{!*���+]�=�$[`��K�WJ���Ot��oS��9V�C���{� ��ƌ�5T�}
1�x�Ez��?H�����|�G4��9_H<:�����޽{���>�ؼ�{�|�ڭ����mRi��9�>�!�d�%\�������*�9��1C��A�x�{�3�����xÙ}�����?p=U�A[�w줏|�#�LH\����+�p,��!)V���;�@����}����3����*���]�aa�;eJ���ԃ}���q��/S���iylʔ��T�t{��=o���/f�k�CǞ���ߣ�3NT�Dd�ݕ���v�jl��*6����t���L]���)���?��!���
���#3�|���㯣^اF3��/���8Ql��Q]�������{�m�~�Zz�)CP�����u-��q��~+�)��^�J#ׅQ�����X��M)AŦcSX>0Ώ�J�|Lݐf�,噵�9�mq�U�o��)ÑD-D��%rxU�q�xØ����Z��<;i~,�����Dj�AC;i�zV�)2B���!�y���F�c��ήU���sނ���z��^�mfӳgkԄL͈�bGkl��7�M8��pę)3��Qe�ж���cY�S6���D���"��v�s��͖���/$��:v-�Sr [����{v.]���h��#'�g��C�u���-�|ڌ�e�<y�� �/��"]wݵ#����n�JSS�	b@�͛6�����@U���4�q#ڄ��k]�WzY�ؙ�.[l`LMM������ލ7�H�]v�m2�L���������C^z�%ަ��X��D���������x
�iirUvBk�[����Tf9�ٽ{/��n��uR���ulA�#��>:uj��(x��3[f���G^����.m����A5�!eggg��oz+�.m�[��o�ۿ�o������D�n�&&&�Z�3�6mⅨ�V����f�C ���[y�����R7�t�s��4��V�6��&��k�5�s�N��]����H���'����rD��ַ�Ņ�#�qH��_1�5�u%u�y{����;�s;����b+j��,b1�J�Ӆ���e��7�������ƙ�7�D"����� w��{_���'��t�:dF'��g�eFD>���4l��20zw��M�;f����0��ꫮ�cG��>�{_�����g����7Ļ��khrb�p�6���K���ZB"�s�%t��Q:~�8]w͵���e�-��Jr4fHo��&jc%�,⛦�[n�ٸ��ѭ�*w%�� kc�ٿ����'�|2#3�2�"j��-F�7�o�=����W^y�L��K ��&F0D�Ơh6[f�l;k�ā3u��~�'\a�1c
_��B6n���Tr .�}1����7�q-{\�?u�~���a&''�����{��~� !�' L����.�0�">� _�0#O�z&�^r���0p
α�@6����Y��	�HE)��c�c�f��h��M�MYI�����Z�w�/51�1D�eĒQ������� _��1�����1&&���\@/��'�1�[7f
�0^ 
�0G����?�J6�r���w���}��L�����\�5�oR&�R8>(�� �.�p��� �]>KK��E������E������h]�+��š2�	|:F�׿����b[8�b
��Qox�$}�_�g��9}@ʀ`0%} Q'�����aR��V6�����ݷo?s��ï��1H���\���?��!��R�֭xO1e';kֿLǎc�ˇ�'�X|����Cbe	g�e���ո��D�!�e�'�хp��Y�� ��ia
����s�џz�)>)�plʃX<� 0�)�|ꩧ��KD����O����YԂ+~�c�<�H߿���&�������-6dfgw������}��S,�ADL���KB	��#�<�\��!o!��L�F�@��f���
]P��7p�%���'���:X�9~��3p8 � ��1�
�u�iE�o��f���~�3H(��KL����'F1�����z��ޯ}�kə\�;���g�v��������ԧ>����%�Hǻ�����)}�K_���1����w��k�e����Bi@����>�v���3G��@��`����@���+3��	���>�HYp��g���{6H6�ca�ǐúR���!�1A�B6���S`_�{@ ����"�` �]��A /�{�E��ڂ��u�Q�Q��H(��lڃip� �F{�J����w�сlۨ��L��aų*�zBB% |����#X����SSS#�"߫��8�GD��U����h�krH���ndĚ�����)�=<{�h=�O�e��0Q 
.���A j�:�u�L��x�U&f�z�f?+��	��N�x�����~ױ��oA	�o9��<�?dN����R�)�| M�,������A���¡*C8���K��� s�$8�$qYx
J�V��'����Jw�
_�΀9[��AF��\V��_�ubgbN�tlq��c��Pn6ô��ix�ad���S���e��R�s����8ۊ~�C�	|���F���U���vl�c1í5@U�� ��D�G�A�$�?v6 C��c�/�Ed�b5�-�u D~Wv� M�N"A���G �����j�O���-:��LAB9����pe�߈aA߬���3VCD D RAL��[^� RQO>4R�)hR�l /���|��h�,���Q�uǈ�Q�$ g�mF���ˮ�#�,˒�ğ*+�w��*�`g���}��A$�\F�蘵��|��DE�	��L�!"���V�Ћ OIWEj����Ea~�i:�8�2x�+���>��0�@L�b�n��R���<�;��N&2��
"�^f=����l̽�G0����@Y?�R�����s�qp��pgF�� V���?Ρẋ`$B�6�)�����Q�oDv�P�
�(X���h��A�6DdƲ
 �@��������@g�S�pq6 s�}$����e��tC�@(��0߁h����X�
�ozӛ��65)���i�*�
Đ9|;��
/g*9/"���w~���/���X��I��� �jF!ʡ|Q��������&Q��FB%AD��s�c��|�G㗿��$�����_t�s(u�t���?�^�@k5dV#�27d���V~�S>��O�����&-A��R5�9v�OxZ�3�«[��}�����H�Hg�;��[�VM]�P�2��iW������u&�p����	'��/�@rӄ蒇PFZY"k�R���_=#���I��d@�!*~ D�;ZQV�`���ʰVy�U�Y�yD�"��	�@����v��窛�q�O|��!����C�Y	�UE�g%KQ��9,��_����L�ӽ�~;B�|v~@r����Od�����yN/���s2:��:**��xy��|��̶yT�C�	�T͙�:�X��{v1O>��>�@PQ���7����C����, :�qC#�|���D�0G��0N>t"����)��Q�r�eV�䐕žF��?4Uu�Qr���Ͳ�UP�h��n���'���Ea������cw*["��6Y�m�eɪ��;mdTk~(�0/;655�{����'��l��[����q����s+�� x�̌6�����e��R�r�-k�������lQ�3���S�%�oS�i<��c靈H������ �_l|��>q/�-�0��j�/��_<1��}|��y>���'��
8�ꚾ}�XF���.���y.��g��@��<���8P^3߾��{������� gF�}�ڣ���|�9d��<}�\������ ��7��C�s�<W�j�E;���;���|Q�50:���%bm�w����w�;�M��*���W��U:ۀ�03:�����H��:t臦�w����)������&��|����!���|�m>���Q�g�}o3C��䪈 v����͆�҆�c���E�׌�c���'�Ȕ�!���m��m�0�m�^��q���I���D�[߹6���4L�g;�+�!��X��ʾAPF� X��-�*"�����"�ԃ>�%�?�-��E��_c����#�K���É��o��!a_e::�=o�.!��G�]E>�_%[�bInlAR!��%#u�����o��e%P�i��Æ��iDW�qHTyΔ�ͺ��<�˯��A)A6J 6��h�@�B�Te�a�?�|�m۶g��۫�� 1������0`�)U��Jz�镢H��Rr_�SV�d�xPw�*�$�RR}<*���p���"���2
�*F�0�h��?�я�ϲXȆe���-e6��B�y�K%��dp�ߓ����n�����R�TYY�O�tЪuc��i��C�R�A��S�x�R����8�y����H�)��WWe�xbj��nJ���=��UY�ѫk^;k��!*=�SW!��]r����xl��*��Q	mN�!�2��M���e�!zT�͈>�Cܤ�y�x�z�r|��a�0O+9f�3�3�T�sO�;(#He,��2R�]^*��C~��F��+A*���P��r�<�UV����"YѲ�-��<m�(�:����O6z>T)B���)Y�؍;#�{�E@�(6Ȋk*�B�x5"w�����{�U{�xP�T�"o�gY�s�C�ܼ�Og���}cK@�P�$8y�Ω;("J\)e�T�nmI����å����:)T�H��!e6�w�ΥDל�T� ��5��0�,I�(q"x���}�0o�s��~W�Ժ"��qk4*�͇����j�σ9(�kH����"ιdk�7Rԇ���>SG��zs����h���\]';rD�/    IEND�B`�PK
     C"BY���+� +� /   images/c49304c6-1828-42f7-9c78-6513b79a7c1a.png�PNG

   IHDR  p  �   �#I   gAMA  ���a   	pHYs  �  ��+  ��IDATx��y�$�}����ꞙ���c��.��  HIH$hP4)Yv�r�Ö�2Ç�p�4�p8�v8"-G�RP�EC�dP$x�$	,.b��b{ �;gOwWe��|W�ˣ��kz��g>����|���˗��o�~��V                ��Q                8Tp                28                                �               �C               �!��               ��A�               p� �                8dp                28                                �               �C               �!��               ��A�               p� �                8dp                28                                �               �C               �!��               ��A�     7*�����"�����b��P*��s���*B��l�.         8     �FC�ʜ:����=s�/�}��/�j��(&��m����w���[o����D7����W����{�����_��u�V�Tu��^��λ�����/�r˩/��^         p� �     ��[}�����?��/|�{��ݹp�|n7��ZJU��x�ԩo��-o�������+��[�Ʋơ��x�s����g~��ֹ�vf���2��PJ�N&ř���������s�=�~��g��X         k��     n$��9s���/?�w���w~����[�B���\E!*S	!���������N7��׽�u�[�o�D�PU��o|����ß���{��VǬ�R8�F�|>��2�'�z�O�S���c?�©[N=To�         �68     ���Z+����_~���z��o�eg����8�b:��κD�׈٬<q�����s��=w���ӧO?[������/��3���{^���QJ�P��)�3��0r.*[��ۧ{������_�;��WZ���E         �Z �     �)�:{��K{��o��ݽ�z�ҭZI��*a����B�ey����g�~�5�O������e�8��o=���{�5R�R�,R>���� ������}���|�;���ں��ɛ_�:         X     p�P�={�%;;��#6��ްDQ^v�~�i�e)lU�*S�o}�����׼L��9q=�Q���sۙ3/�g�=%��J>_�v�S�<�2��8���l�y�ܙ��9s�e7�|˗�X�         X     p�Pl]ܺ���O9o)�3��lI8+"���R/QL
QV����g��fN��V��Enoo�~�ҥ{��6��R))���:��X�7"��1B�u����-��.�.�����R        pA�     7
j6�����(���@�(�m���0��8aJQo,'���M���&L\���l~rw�{�R����<	[���3GZ+�?�)]g������;�'�P��        `mp     ��BQU�1!�D9�/L�7��zU��
%+a��C*c�FY�"8�g�˟jn�WVj'��S��%�p���V	'�1Ҫ�4����`|	        pY0�     7
N��i��/HP�oJ��}�p�6���_�U5��g�s������*'��M�hBDK%!����`���j*_        \L�    ��B1/�UUM��2X�j2��N���λ���:+׻�G}�v�T�TIg��x�2>���o��zA�7Vb��FI[	]�.Z         �� �     �or�2�fiMa�u	��ۗ��N���(E	�B�+�N(n �0�U���QA�a��6,\�)�sZ��*��         �     �Q��:&�����h'6�Jj�Z����}J�#�`�����u/�p�F���"%Y'���!g��Y���ʹ5�	`l>n���        ����     n�5�T�ffXk����V��u�#�6��XAk-�0��T�D��q㲡�ϹJ���&��ϣ�O޽L���������        `p     ���u5�JKgaCz���D�2X�0�٠��Q���s&RXkoVI5�ż(
k� #�]�8C)�cq�V��'rq�         ��     �8��f��Sifs�ċD�6a�P���cu���67��Vi�
V\�X����ظ��S��M)�/��3����Y'��ʉ7*���
         �     �p�#&N�a���V��Dt���[H�l�e'ސ�9Q��\)��w��Y�ؚn��UY��e��(���伧��NŖ�[U�����G         W     p�c��i�y���\O����En�7��]�!�Q��V�z����8v���+���}��BϦ�b�אE���ܤxO*J{ц�J/(����(���nt���        `Mp     �u��֩�R�[�w�d㎍'��R��FتR!U����ZŖ��p��8YV���ƻ�1;R���׏��EJ9�ޢ��WYy�D���s�R�(�jR���pH�v<q�&y뭷n(�N�q]�?��R1        �>@�     �#�Z{Җ�K�>��7}�K_��3�������O����NQ*�C�)�5��R[�g�yq�B�����0��N>���g���7���7<x��_QߒRn��ʹΣ[ϝ;��3O?�گ|�o}���ړO=��n9�P���������J�G����Yۘ���q�m�}�?yӛ~��?�C���=���[n��	��w�<�         X	     p�����͞?�������#��o���o>��ͳ�mӶؔ�Զ�2B�`HC9S�]��Xa*+*-ť�+��O|�u��_{����]����~�����j�E)�9q4����_����ۿ��?�����k�=��]e9;!��)m�5V�*�p��Υ�u�k�l^���6������x�����'����}�{�m�k�g[         �Rp     ���4eu�c��������������������b^�eY�#6u!L��)���'��B���q�%��O�[fr��V1�ܧ^��߼뙯|�����~����W�I�8bXkO|���_�������c����޽y2)��V9��(��3É5�zC�N�[�pYbM}��N'��湴����'���O<��/<��W|����_��_��S�N=To�         �	     ���x�[O��'�����N���W��.��D������4Z��i7���LP��R'P��j������m)��ʉV��������>'.���_y�8��P��Qr��/mߟ�ɟ��=����o.T!e%���ʖ���_A�a�񿝋��Xo�ùYq;ʲ��������}�ЇĻ�������3�����         �=A�     �'����^9y���ni�;p����JZ���B�5�+�bCG*FTQ�!��'���Xa��U�n�[�䤜Ow?������W��=�K��Gkŉ��<����x��ٛT}F��]g�R�[��7TȋF�a�X# �f�lt4a\^+9��N�/m���?��[~�=?����旄��         A�     ��2'/<��WllomVR���ı�J��CI�
!e�]�x�F�⿣���o��C;�!�^W:�,���g�0�Ο|��o���}��~�m?}�s����Gnoo��я����Է�3����D(�dR:�c��[Hܦ�<��:o2'�7-�c��Ȣ��J�{{����������~����7M �         �     p�P�vo���_�3)��Z�M#E��P�^�!��C�-L(/�0^� �H�hA�����[�����s�RY[�b2۞���k/|��;~�gabK\��sg������a��(�DJ5�J+���n(g}D���r��<R^���~��d�����j��/�������^���d:�~W         �Bp     ���4;�ͭg��YZ+������I�2q)d��@A*��3��@��EN�`�D��lx��E���4���}ﶝ��{�x���#"�x�̙�Ξ;s��*�,nL���ċ\�R�B���ަ�1�����?D)�1VL&QV����s���C/��϶ON�Ӡ        �Qp     �uCUUE�;��NW`��^�1�	8������ʠ$�N� UTذ�l/��0���"�R�J�ʅ���vw7D�r�����j^mZk��7�r�ލJ$eG����8�D2��kg�����o��:�f1�a�	        �&�     ���X5��j��ն^t�@�x�	9��XD�"z �:�l$��A�og��[�p�%�[��%#Jg�CZ��h��0��'����RRV.;���?���;�Ig՜]4�!BX�s�v>N�>.��c�U��         �'8     ��Z#*-���Ѳ��V6�� :
�i$�)R4���I��]��`��TNȡ�?�:o���)˲���,�[��)���M�H+RV��z9�TY�[�ֶ�)�L�         8     ��AJ��Q�I�s"�F���g��5��5����FfjB�hy#���7>alXv&*#gN������*�R��y�ŝU�#6	9Tc]Ó�/Rv�.>?2�n[��]���*[:��         �'8     ����j���(+�4R��K4�a��!Z��$��$үd2"	+�BE��ܡ�Uٍ��Z㌋(/P�]�!R���"�-�:�wʛ��g�ĻR�8��:-         `Op     ����*STU��nH�$�:�N����`�� JF�6(:�`�"��&�
�U>��J�J�q�rp�a��Z�����B���$T���#f�i�-�2�o�ca����V�T8         ���     ���.Q:A�WXh����霪��ř�P���=J��s�ad�B%(����?+�>�>\%�)�#�Ӣ��p�\�d�Q�w������\Б�P�"� ��pc���        �C     \'Hk��fRU3c��X��J�ʈ�.�5�Z9����ڍ�&$h9��A�o��	������ة��ь�5Z����82Y�se�|���[	m�p�N���N����[.I�R�����%hZ�rT��r��x�L_         # �     �����5��V������ٕb6�ڂ�I
�0C��%jd�(���<l#HPƈ�X�ܺB���lD�[mg��0��6绻�yY��T��*�N%WT��DK�`�C5V:D�dA�Z�0e5��|.�!wf3]��D         �� �     �����O����������ܶa��+%�T9G*��%�xC	��%�`A"^��NDw 2Y��!\!�vC��Y�(+�)��̳��Nջ��C��]��<R��ę�޵�5���嬑���PLq�ƥJp��D&X-�gN���G6��
���Voo_�ekk��i!&u���        �C     e������s�ų?�����{��}��*!����*��Jz� N��nG|�D+AS`����dt���
��V:�j�+O�nol}��~���~���^�����O����ŵ��d��YU�˟}��w~�3�����m�:��E1�N�ш6�^�Y�h��ok�'_����弨8�$ƈ�,��d���O<�я}�o����sq:�~���{�CA�        �     E�(�&�={勏������}˹������Y�(��ZL�gi�I6��T�'Y���	�`��a���@��đ,S��vEO'b������ū?�_��z�����N��_{�o���'^r�g�@�"�!�6��{������/����_z��|�/��|�x1QB:�K�Ep?#m���.E6�mf��6"�/��RZN&���g�ųg����_��W���_����mo{��x�������x��Y��        ���     ��޾������_�����G�䍗�|�����M�/�ۘ���pR��ʉ1�b�(��҃�"D��S<^� E�ё�
�[ސ1�īA�P���j~���?��?�*}���;��η��?���~��Q��8��l~�G>�������;>��?�)g�O&��lV�w�T**�F�!e��"��r�)�X��e�D����Xf:٨�SO�{�����o���ߟ���y��O��G��C��?�������hpG               8ZXkO=���������?���'�`.�;y��Վ�b��pv7���p2��B���А����gE���p�7dc��.��A�V������ڊ�hav����x��|����~�����e�}D\}��,�������������}����JI]���e�lP����X�`mkyC$�G&�V:���!�vZ%+�6��g�=���/>����dZ����mss�[+         8     �h�u��k���׿_����6��N�(�H#�Dy�Rk�\x8Z�0��e��-�0��Ʋ�R*���O+g��}�Ue%�(��*!�\ݲ3;���'������O����_���7��E�;w�������g�s�0��:��(�u�(�u�I����F�NF��}J��-�Wъ�q�S���^�E>�5F���_��l6��ٽ�S>��'�x������vh&         npp     �QB���W^���_�1�4��JU8Q�SS(at�ܤ)�U��S��MH+O�׸�Fȑ-{"�Ve럺>�*|H[�EYZu���7?��?}�����8�җ>*���	��u�.�|�����Ɇ,��N&Q��)7Z��l4*!'�Ɇ��ˎD�β��y�����l>�����=w���>��7����^_?        pÃ�     �����[�N:sޓ���"��L��Z��s�`#y�ɠF\�D�gn�#�F�X��.C��!Ʃ� �8��^p��lUUR<�Խ�O<��/}醸�nT���OU3�1-6d-n�Ƌ7T�$"���ż�5�_����ֱ�!;���0�_�,ugɤ�-�X�w/m���W����lv�cǶnT        �     %�|6���('�h%�N���o忽܁(�ʀ$4h
���On�"�D��#��uh#�R��N��3�m����9?{�dhRv��(ȋ/�ܝ]�ι�5b�&B�sRZ(����|J����1�F �l,w$�F�h�1�z-��!�s(!6&S1/w��l6=w��-UU��|��         ��A�     G	e�xC����!��*Ż Q~9y<ɭH����
':�B��T�:X�i����E	��qYw\Sɲ�VX1FU�]'����"�wv6Mi
��?Z�����[g�s��l�Rt]��ζN,>�¾�:Y�����FY�,��f3]��>�T,�t        �     p������V'�PJX�ù�:�IB��hD��h-oсs� Fp��r}�"A<�|�Υ��ڙ�eU	Q����N�\�&r�;�Xc�TJz�JykAh]�x�K�-c���I+�Hw||�cK�q��p���J               8R([)����H�;� ��D���r�����c��B�u��lnDч]w)=rA��a�E�`��#1UЄ̍�������J�T^���u/nqCt�%T#�ȅ}A��:G�͊��F�2m���9�h�D���UU���         8     �H��:Yب?^���o����Hz�G��4R���l�Q�!��&��/Bp�@T,����V�[Q��H�h��\]��ҥ5�
�E�N礒q��y�M���D�$�F&�B�ur����I۰�         p     ���ؘ���-kx����N(�B4�$a�[|�t�n�]AC!d+DPxx�B��E^�P����mQ��DU�-�ð,�,[hg��	%�9��+c���G�<�KF�����v�1�)~/��u>Y�o         $p     ������8�0^�a���Ԅl� �h`��#�5�����H�/p���%El{;	�E�ɲ���P�	eY�����iPʶb;���̅Jnu#w�����&���ݱ�c��R�G        �     p�.=��'�����F+�Uf$#���ICn"�4��o�#�F!lO��1x	���\���}���q(8���X��j��D/u��l��Q��v[r�⾝K����{{CIQ'q��4fL         npp     ��C9� �MGp�"IF2� ��L@ ��pF��$o)=�I�����Ǧ�(�4T������J�eY�ʪ����%�^"���'F�&��E�:�Kk������ʅW*�3         xp     ���TF��[nRj�dH�dH��7��1��"�Ȭu$�Ar"�C�`Iæ�6�)�pÈx�ݷ�o�w�"D�
g"�0$
r>�-��$Z�i[EGȑ�O�D�m��l+I8K��&�[��]I��0��_��cU�~        pÃ�     �^#Q	�]�x-�RV�AX��fD�������&
<�1'=�ɯ�����)�G�1� �h���kE��HU;�֧����&T�U�pخEOf%���a�ޮU���Ζl�OǚG\�n}U�        �     p�����r.�3p!��A<�e�����"-�B]���x�dI���҆���LËA�����Y����N�`�ϼ5�Ӧ����E�P�LYJk�TE5������n ����?0&��-o����7�rU���        @     )*c�N��c���K��S��b��TG1���b��»Ri��3�hG{���ܦ$����[��lz8��ʆ�e�c��e����J��������u	Y����*�Ӥ��Չ^�W����X�H
�=���-y�B�dq#Xݨ�|
�.\Y:8         8     �h��-����DJc�\!�J(�+T��^C�*R^�!������ܢ4�hI�3�U��i�v2o��2&:�p�?�H�z��3'Q�3��S���*�T��S�*SIYQ�M8!Gs��1!G����l�%JZ�wɒ¶.S*�6��:}��              p�p
�ܔ(k�-
��.�t�.�siD����u2�Va��6�Y�P��	A�!� $��p��� �%FIQ���5���e���!��(c�.M�WeV8�v�M�⊎@Ctd(}W,i��w����W}��n         $p     ��B&aF���4 ��E����ܷ�����:D4�1D�J�Blcr���'~���$I�Vd����V*X��Oea�V=����Hk�L�RrAF9_���N�4�>})Ng��{����.���        �     -��U����Bǧ�R
��m4�5�����jEaCF$F��c±����5�txaGp���Z�T7�����Q+�/�����o2��u{�w��������lE         ��     �Vff���J�'Qi�lD���"�h�#
����v��*���"�ǔ��FH&h�^�a��C���uv@C����g�u�׎X�paMO��,w4f�$�'m��^E6:º<>�_ZQG��]&              1�CU*+�XBy!��F0T=�qj c���(��H��#,�x�A�`�X#�BLJ��(� Aà��#8ك[�*#�1N:���E��S��Q���)��\�yA�A��Zqy`�l��U"7�\̘��QI��I b���(e��t��T�D"        ��A�     G	e*����NTa�P�[X�E�i�x�"X���HRTw]�/���F��d��
�I�1A��
��8�����mq(1t��2J4��ݼ���#Y҈�kL�.}W*";wAc����               8J(a�n%A���X��hi9��ը/��#�dr�ұ�a�G˅��gE4L��yMq�#���5�b]B���Xr�gVW����U&���I�A�0#Z�H���@d(�h��$)i�,���        pm��     �N9!�5ҹ�p:'�pB�l�@���z���3��H_50t�2p��jxC���S$W*���D�����K� +����	l���RT:��J�ȴQ��^����zE�|m,��$��ҙ�X}�F:P0��t���        �     p�0�(*Yh#�Z~�F&dt�p���m�^K��&���+���'�T�.@��
�
��۝��`��&i�����ժ8a�=�9�M&����U^E!�A|:�/>�I���DZ�Fr�"�0"Y�0Q�њ�h��[�N}AL徕�L7J)Ո�        �     p�PZ*�!
;w��� �PAY �)�RE��T��o�CD�	�mn�\�+9���Tj*����5h�"�p,pxaDQ�Rkm���!��E*�qY�Z��
8d��4�$��/G���nU�Rg��������5231-&FJy"        �k��%����C6}    p�$����׏��a~a�����-k�	�4�:�»2����V2��������#���+脈�j�i<\|FJ1�?��bWm[l66?�x��<8l/�(���Fh/ؐYD��$��\��N��1+��eA��a�Q��\�b�EU�ʘj�^��j�Ee
   �O�j���+��pT�  ��+&��꺟�,���d{X��5��4��SC��\�����/�<_�
an�l,˻�c�rM�3��� Y�\�a_�ܨ�>�УϵZn�MW��<��~/��m���>��v/n�T��>f'�TQ{Q�>���_J_\`r����%uh"	r����6ڧ(���a�rYG>�Ӱ���f�[힬�F'����s�O��.�6�������Ϝ={�����Ԫ��DN�ъ0��#�H�w�R�V�����υ ��w͌1jk{��������[���t���^u�]qݺ\���r�}�ھk�M]6>9��*���Z�n�õ|���&W�]g��+��B]g��zn#.����׎|7G=���> ���A8\#;�?7����������;�;Ǫ��VU�msXg�78QVR���J%÷h&���3��_���6��'=�{��B�s�6K�H�΁���e�V��g쏸V�7i��(c�v�Z۞��'�?�2{��v�.��������������.*�{1܅{���e�T�b׫�F�#��3~g}���_�0��h{O��a7;r-�_+6��W�u�ؾX5�c�I���Qq�H���+��e��:n��
�А�]���<P���qv�M����~��B*_6���m���=˷R6�5��>{㋝���4F���܎�~v�+m˺���A��MJz�1���F����Ap�a[��O���b^�7y[��\m�� ��wd8�.t9)&�.&3������~����q;;6�yS�ɴ��u=��޲����̳^� �޶C����#��M^�D��2�Mȼ�iV���Ӵ�v\z����߾��O��g�>Le�)+]�J�x��(&B
�6���?i۱�r�%�����}W��e1�̦�b�}��_y�+���?�؛g���в���LHo�~b��ܷ�1f�#���Ŵ�#y�,��s��P��J��O���������mln���|�5V	o�Dɔ�	�1�O��o��m�Ֆ�������2UJg�퇑�°G]-����H�d�m�mʝOk�i"�*�88ݥ�
j��Y���SLP��l�a�M�4c�N��8��]���Z�UA��W/��]�����r�c�Xp���8�\�}�5�f�A��7x=ȹ�}3>���=xBe3j�*�x߈V��gϘ��P�j�5��$Dޕlʺ�ˢ�+:�[ۮ��r�^���k���ܒ?�l�uv���=���.����'�Y0g� �;F��5rNñ������胊f��]�[��B^ͥ����z���ZB�8Mcaی�cm7эn\?�i%�z�d�VUQ�B빮?u�q�{���|�}��lן��w  �2����C��ݳs�Γ-�Y��p�����۟z�~��O�З���W}�o�y�c��UY)7�[�JK��qa�^�K�IK���TD�Գ	�k����ݧ�"�߶?�%�a�mwxCm�t��
�;�x"M����XP�1�|�J��õs�b����l��[��pe�᝭ꨵ]�\o[fO�믲�Gs���}4̑���zeìP��t.ӭ����dV7,"Yt*���r����<ú�a���U������~�Qz�X�*�n���+X&�$<[
���ƽ�\����U��w��d��l�l��q��D������=�?����u�a�hS}��%�t�;�3��Z��^jp{Ծ~8Fw7�֬S^>d6���K�jG۸}���E�a�,g�����K�=M]a�b��2vp�ޱ/���a\������{�t'�\_�����隍���_����ֲ�鄆�����>3�jt0A��{�?b%���:1��olS��!���e��G5ì�Zۦ�=�?7WET�c�$Nqy⏞N�dՇ�/�Mw��_��^�|=&��B�1|=�퇫�B��q���C)e'�v{���gIB��q����fn}�F%�с�f]m��eiU����$*1~��{�֟��h�St��E���o��H����������������-�nUg�����g�T�������M7�
���z	�oTV;W'�__T]N&����r,=�V9��پ����cc:)�tI���ӤLh��,q䂎�}[��1VXv�\���(�P޵�Do]:������׿���\����eu�)��QT�����(>���<��-��Jg\��<�@�������_�����;F�H���E4b|����E}`'Z��	�䶊1fg�k�m3�/�M��2�V7�p�5�/��Uu�����vg<�~���ص�_Q�<C��F�Ն�p��m��EFX��:��N���b�V�Zeߢ�r�8��y$���Y��4��_F�iH�/����I�Ӈ5�p�a˲�AF�M��-n�o�C��*ñ�?t�K8�nX|=�Z��uA"R�ڷ�X1p/�����j<��c�<���h���;Hq�G!n#��}���&H��`s���$���*5Rew<���ʚ�S��x��d���W���6�g���ٻ��~�\�n�/�N�v��>�K�c\quw]�R1M�_�V�CT���+R�`a!DT�.�Ҷ�F��z��i�O���i��*i�i��
�[�7�]w�Zu���Ns��I_sO#�h`�����3�b%�t0:oQw���c�0�ʤ���M�n<�ʆ��q�_���|�m�.B�߾fke05�<�6#W{)U8��3��m��)���c3ݘ�O��y瞻�>�����W���߼��{��Oω ��0t_�m�$$q�&��M�-��L���ZM6� F�[��Yr�x��=�O���Y����k�~� ]�z/q�ɷ<9�gl��16pUg�W�S����[i�k���Y��s5vX���E�L����)���E��K��u#�X��~�I�H{����_��a�f�a����H6�i�dS�����:�:������ٽ�g����ڕ�Ϛ&:��u��WY*˱��i��6i�hu+��r2	cse���H���m��� ��(��8�U�w�+�v�Ϭn{�g��8�q���p�L8��w�~����������÷���wl���|>۬;��*�9(a�t�h�6��y|�;_H�"�0��!j�9&����l��{9�c �����Z�-a;2���#3^�hd�C�-���*ebQU�sP��AŽ�I�o�W�܏��`ݟ���F�.�g9����uy�_پ=j;o_���=�0��s���U�Uc���H��Ķ���}U`�3{��?؉������T�������!�h	�{�3ݺ ���̆"�a^�&{ߎj	^�,����3����~�s-�H��1fv�#���Q\�,,>�H������ц,���Wok���>wރE���\_��_���Nw^�lީ���v*��c� �i"II����T�����X׈�.?�h,���2�.���}��t�'>��q��Jf_�u{�M�U�;L)��:?��p�t�.�օЪ�G�C��d*7&9�t�A&vW��Wy8A�{�,��$�84�����!�f��s�Ᏺ��E)zc�86I3��	ci�G�b"6�*��'�緎?���+[	iJ'�i�[�"泉㤦l��l�����R�G�?��u	Vbcc�?!�z"���ŢTs�%���O��{�;�	6򸓀Ý�t�a��������^�x�[_UU8� ��U޸̋��W����d�4�H���6���h���c/��Gw*^� ÷	F�I�<���щ��l��/�}!��Q�2�:��9�c�$����룛ꢹǳ��[tV�nD�?VIu�?�V�⮁?��CPa�Z*Eׯ�F�u��p�qm�:��c���8h����=�]��5&_�A��]Vm�f���F�S�w�7&p��ׇ��8g��5S��}���C�����uz0;<�<L~_�T�B��쪬o�n���f����7ۣ�������[Y_3J��8K):���qޱ7~�<9:?->�@�al�®�n�1ŕ�J{������ �Y�v곴�������N���͟��e��؇�]7���+�C�$ڞAB|�2�"�����y��g�o��+�I<��p�Ο�7S�x�[�Kû�ߙ��~���Hs)A��t�mև��zD֗i,�8\4&6�J���4�N��26��c3Ѫ,���w�}ׅ�����N�t��(3��SJ[���ƹy��F����|��5^�]�Wd�u[À�0�$Nir�W �w̙D���i��_��@�3i����e��<�;N�����ˏ�v�v7��\'����&���;/\�0���N�lE��vN��Pc`/�"���{R�e�Z&��A�8ӘNY��I�&�M?�11��P�d|�_N	Mf���;�ߧ#�Ͷ�m��O����N\��X1�ItrE��pڇis�Sw��otħ����6]���6�v&Nq�7h:�X���z�&!�XPƞ�&��J�SO�"��(����XY.�.��"�_���5k��4�.̐�v��	����e�h������r�ϲ����n�e8}۽�MZ�eM��b�^pI��F�^��/}�N1�����퐄�Ny�TW)\��o
ټ͕�Y�(���Ux1N�u~�ֹ����V�_M�[Rq�`��W�$�ʗC&�L|�!��u�l�,��Ʀ�����qf�m���0-�tC�ï�����6N��٬���Е�?EQ��I1�L6��vǥ�^z��ӧO?�<v�K^�z�wE�sx9wr'���_��#�����꯾���5�ϝ���rjf�RU!7&Sa�8@���%Ԅ���O�$Y��d�u�~�؀l��Hq��AX;�<�g�c����� �sꋌ\��떫i_�.Y^�U�|��Y��\k���e��P��̒�ֹf�}��O`�B��]�f��=�J˟��o����]7�e�u����(�Q4�l��/���'\�鍤��<�Ha�$��ɟu����E�4H��X��
��l�D,��ފ|�H��	�����ĸ��~$�
��ԋf�У���w��,�g���I&��%��r߯[���*'�~�_힖ݟ���m�t釽Bd]�a��?M*I���#z���lGc~o�Ė��1={Uϝ�c�ُR.�b��s���Q��cS]�ɢ�o��L6&��Z�L�6����j>�(�q�e�����B+Q:� �(���P��1�B�'?�؅h_[m��l��PPeE�-6e��X�l�w�%Qxg���Ȼ�Jn�I=���-�c/�Ad��	���y�F|�,�H���&�ma�񽙔&7!�欼K9	�ݿ�|�D�Hq>\v��h�Hh��e�e6~[��0�}�P��ETk�	�fz$^����\~������U�T�m�r�1ㄒ*R)���;��U/��W�6�fU�jW��z�ZS����0�^B�2ec�3,	j����u���g��T?)����|Μ#�a�*�ܑT�ݜ��GY��y���X�<��P댓��`]����H':�A{UƎ?r���Mu����]w��1>g;�hG��c��t�kcz����#7+z/���W�{/�n�*6�O�����dݡ�:���#�� {Ʈ}^_�׻�k�������1]��?���=�!�v�U6�5r֝�Z�����*g?��d����U����W���~��n�2㬟�uǎ}���K��l���Y@.f�[���;�v��i��*cu����fE'\w.)���x��=ƈ���UU�2f?g�r�qESd��Bxg�~��gש�����u4��0~J��'��{�'�L��t>Uئ�I�L)ØC�e=l�����:�c��ս�(�D�2��7�б�'���.���A��.�RӖ�Ft�(=��Q��V#J������!z������S���R|k��T�FT����.�� $+��lA�Ҋr#Ҙ�$���ً+����w�HI��R}�NLv�:�^t��c���=�x���]�Oं�n�$�oD��N"Xu���_���<�lϭ���O�3T��C�rш�r��:"�t�J6/=t���6�b��{QA�m*|/	�(6+�2Z��\��=,ZP��V�#��At_��MI�soY�&ZہݣtMW��b�J�f��v)S��DMQ����#�{���������fATZ�ϭ��n
E�G�1e�t�h��[��b�j^��Ʒq�<����ꋤ�৹�݂�[�5ːN]��Ci�+�`�7e�id����K�r�����)SB��t�ӌJS��Tw�$0t�x��p�^U�׽Ʌ�y������%(��Xךm���cǷ�.ο���<��������{�_�u�ݟ�Z?/��F�w^��;O�����7?�G����η���ŭ��3R���M��s��R����w���� �oi�n&�R�:��x��H����:��Ҭf4"��|�����/Zg�����|Pb���De���h�
�,�
��p�؄ば�i�Ղ�5�-�sQI�����qy"�5��j���HV�~��Oؕ�l(���ߪy6~�%[�zQ˶q�_O����n�{m�RR�_��>k{�^�6ul۵��f�4�P��ۗq����N�pugy	��8������PJ.��^t�u*���Q��g�xB[zq�mk�WySq��Z����`W8��<�p�N�j��W�+��<�-N��˷�X�vi�EQf;+��P 4��XR5am��m���D'����Q�gun3���c�7�zi��EoL�	���XL;4��lR�.=d��8�f�x��y�9^�n��@>ۈ��w��ᆡ�iK�)��jN<<�2Eo�U�&��5�m���1U�\���NS�g痹lD���0��q��"�~|�盅�sEUYz�#�8��&��A�M���S�P��|r�3^*"�ܔ�n�c��J��&z�S��I��l�i�ګE��~��O�;�*Q�!'�ԟ����n�k�'t��������LW���̎�L�+����tF���_�}��m���%���O;�{$��b��r6q��M7_�Ɋ4��otL����&+���S�ޱ���c��N���?����*m�X�gV� ���.�˷e��H{+��p�U�#��x7]Z�dѽ7t��:���y7��-ݸb��Y!7�γ��62Gb?VD&�]c�|2�d�OXSh��>tw�hy��bA5�����;�Hׯ���mSw�q�0lV��nF�E�`US�{}aa���	fC}��EsM�c��������~��S6F���*QY%�h�P7��ӕ*�B�5ۭQc
k�7�gIrb����0�ӂ�,*W�p)�JL��i�����s���?RO��Ff���%.�_��v�Z�~n��ER�2�2e+�6��R�6{X�l��yf��[��{[~9�����<҃i���l[~G�q���
��iSjC�3���"��neY9QGU4I��Q��^>
i-�wx�'7�y�&	8�q��i/ә�c����eD�G�q�����
��MƇH�6���'�9�$�t_(�s��n�K놭w#V1��'+��C�x��M�
l+�h�OB�l�X���?���S޹��h�w7�,m���f=�Wt��vܜ���4.Y�:�r�B�L�a;�K׾�P6�JR�n���Y���"�Y���j�{o��ј2����鈙��6��B�o~]�>堼��sL[u��N׵wO�sm�k�/�m��5��W����G^�r�I��j���%�]�9��4���f��}�t�doy�~k�S�:7���<�i�r��'��.a���׾�p�u{��+M�)%�UL����ʄ�&����u3�kΞ?k�T��o?�������~�������{����U�[�9�^�uNVrӗ�����_�������+ϟ=s�lVN'��*&ZL
%6�� ��~���#�&^x�5H�m���+��f�h���N&#��I�hTپ+Y+�����RRc7HE���l���b�uň�I�n�g�c�Ĵ���U.����3_'�8cSyc1]��6���x��V�y�{iq�V9Vn�!�Y���%[�?��Vn:6i���H�j�x�{�:���Q�7�����ӱ����X2A1�u��tռ^r�֮wF��%��x[�J�I�*m������e�go���۽��h���;lo����㺵����%��_�2X���!�j��x<��.����`�UO�`�Uv�gi�-�ph߂IQ�y�0�;^bʎ-��V�<�Y�md���4w�Ҧ�=�V�2쵧4W� ],��ռa��^�sY����z,��L�(��0FEz{I��n�KU���n�1���;�tj6$�U>o��o)d�P�}��a2:m���m	�I"c��k�I7c��|�2����nel61�hR�?��������E����'6��e��Q�zI��p2*q/�[�pJ4s0/�&r��q�w�0��cu�̎��k�o��-7i}�2���Q�:=���e�y��#M�4��mD��&Mr�Z�BdaF���kaFӽ��`V�-?��m�*��G���&���J]�~��t�.gd2L�J�:��d�X�e�AA��gU�{˭��G<��2ܱ߇����[�����I�a�M���~��Lz�)���^4<b�V[b,��7vG���d���X���ۍ����4����˯��y��'�*u�^}������L}><��XW9֪T����,?���e�{i�h��g8&��j9=�K����W���X"X��US�?�U����x_خО�r/�cIl�ur�u�/�$�����ʞw6ռ��~]�D�6�}\_���r=ҧl�� !~��!�qU�/���֠�aT�	�6 �Tki/�K��K:ءmc��C�XQey�W�jY�"��M
�ϫ��Ϥ<�*Z/h2��о�`=}�5�g�x�t��]�@�{n�5�6��\h�TR���y���ME�^ވ���-���e��\� b�l�w!���&U6�k�U�� ����I5��>m���')�^�ȯK��h�=�����Av~^�y��6�c�����G�r��9�Q�}�}�>�w]��n�#9����]�<}e3	\���mX�.�����Dڲ��5�ɶ/C�{�#��2&����!C�Ҕ�a�6疷w��f�A�ݷ��u�fi��@s�d��ﭨ)��:�}�T^�yy�G*��M�y��l������˩Ȳ��_�u�<�i���\9P>�u�l��s�]�� �
Z:�l�����ɇ6����2�8�q����l���rƷ	��rV��_���:�v{{{�����˿�K���x������~�رc��%bo�pLϞ;����~�'���#����u�|�=�N��ɤ�:�Ӊ3�[���|!������ym�����&�a1V!�"θ<�a�U(�E�Վ���	����m�IO��ì�v92�Z�Na�Ȇ�5̋��}����V�_G�ai4.#M�pP�K�ج�A���x}LjY��>V���a��g����J���?���r�(�u����)�e�940����A��r���䀼
^���v��VlVoo;��+�~�Q���}��^�lF��ʕ�|��B�*V�6d3��՗�W���he6�\h�,�0���w'A��s��܉,���`]?M���7(����٘��ڀ���G�����:�c�&�HH+�/���"lu��݉������A�"�ͦ�h����fHcsm����yK9��j߮_��2{	F�8�dhrE�܊x�*�Ō�Bw���X��X��M^�m�	$��4~��9��ޛQҢ��N�zVi��uJ;���)ca�"˓�k��Y^��PbQ�4R7�o������{�^��kq�t?}��5��S�c3�i�3�2���q���{�=���C�+ͪ�qPe�J���.��ȸ0�ۛ���<j�s۳����*}�U���Z�f���Ϻ�Uڠ�<��b��\�9�a]}����g�cԜ�h;��|Lާ��;�W�Þ�����I��=�>�rt�7�v
%����Aݣ{�k܃6��c���*�z"�s�3V���Ʈp���,_�\�z]��e�j�G=�����u~>�}~��O�ꉲ�,�[���KSUi�~晧_�?���s'O�x�~��߮ÿ(��u��-���g����~�m;��7�结��cbRL�t���*�vfou!���'���1�U��J��C6�A��?I��Q�uu�j�A)��A-$F�GiB��oy�\c���
�dR������C��D�|�n>�i&��RiԽ�\w�9�{�A���W�?�;���ؗ˾�d��W,�e�;���A�����K���BH1^�|��j�m{��̵�peF��������ػ�������V.3�0K�TlsK��|�@�k��b�︴W$��p,�~����Pq8��X�k��\��^��s����C��������}�ŷ��[�N����)�#�Rg[���)�v�
���� ��N�u������Aul�y��w�Nԋ¶MK'�jVC������hR���yAK}�|�O��ڌ�N)�j�֋�m��C��`��R��{�b�e�u�^3�no�'rQ�y�Ac��4F������1,�P�����K�o)�y��g�H�!�eU�>H��w�M���4(��81O�~X4��B���'��)�� /S�]���8���K.�X�B�ο=��k�.n;�Bz۫o*��̥7x�x;S_����أq���ז�������m��˾o,�zd�y��� ����)�F_+s?�Q��i���`�m{y�ڸp���b�Z\vG�
���E��:��"��Go\o�n�+ܱ�S��Oa���e��.c�U�^��,��{��R��%4g4F���,���e��_��{��1Fw�2��]�X�x��0[5�V��ew6
Q�o;�o��,�g��J"W��#�a?�;(^"��V}�w�E�}����b/� ,�?�Y�A	V)��מ���r^���еZ���{1*>�22��R�1ZU����>��������{��~�'N���:����[�Q��~��7nm]��ҥ�ǎ��8�)�PuJ�"�N)��`'����8���S�P4���H�5�����Ϭ=/���u.�uc���^a�;�k�U*�l�/L_H�<���4���Ƅ\�f�Uv�A��inm�dO�;�_G!�;v3�i���٤.��k&�WIU��H枬���I�6��7�X^d���m������t�y�+'#��"ˑPF��b_4�����[���H\�Z�����F3�>v1R�e8�x+4�iQv��ظ���E.\�$?{�L2��c���/�+ɕ<�5�.�8
i\�5���g����X�kmw]31֯\c{ڈd�ԧ���;!.��Q������\�!Y���C�w�����m�SMٶYi���e�n�]�T������6�:ckr�d���m'�b�����T�����/��Q�P0[ʱ�9�h���,�j��?�I�T^�`W�k��r�/�e�g�F5Or���Z��c����?Aٽ���mwo]D65D�f/�?Ǝ�ԸE��,V-:�������A��knZ����m#:3��0��8�2+׽�Mv��0��!DǅJ�&��R�G��1r�~�U~�l}����6i�m�Nup??L<�1\~=�]$��I4��}~�GM���y(R��SNת��]U�F�Uѽ�#�e�o�
wC'����}�/:�?��K����]K��?�*�qϺ�r�k�����k9Z��k�U�6��պ��5�:ջ���7[g�k�)fy_Pƺ{��}�T߭��9P�PW,�Kn����m�������c����v����d�reI��2�2��[wx��=[&�i\�L��(3Q;QF�F[?�k���Im�/���DJl�����J=�wǺ5e�x@�8�p�Gppr��ߛu����������:sp��!�ǀ���޴ 	���kS\��Q�������ZZz�sp�@3���ƅ�-�*�n	�]gpTPKM�D������chM9hV�2��9�*�،0��{�a��b�_���I�&A��X�@<����"Z����/�ž�e����6�׮T�ӎAZ u��o9S<���K��]������ ��o0�U�V��:2.�dfE�vk�����������_���������o�X�)�gm��7������/�����;���p6�e�ŲX.�=>ef�L�yg�&Y8ӌd�o�a�T���E��" 7��1[O����4�u'q	�c??<�x�]�-�4��&=��3HQ�ó\F�� DG�;�5�� 9Fxe��XPR	�w�$*�F���|1'q>��Aza��ю�y��#��(m�G�s��6P��&6fd1�U;�����\<T�5�z����֯(����Hu��ea&%��$n�n]1z�rc��sGlk����|��!`&��<���3|Yi�������x�z���E`B��U�Ds�y`���+uW����<pS�����+$�}J�����y�"8o'u)*��d����Y5���]Gϻl�k�6�R���B�o,3���������M�p�ڑ�*�k �+i-�dX���fb��U�/ 5	�Y-�^p�:�$EӬ}->�3`����MC��^��F[���&h���n�N��э2Pp�T-�l��>�����PC�Eig�{͗Y]�+V$���S�t���M4~<M��������,w���^�_U
R��_��.^r-��T�։�]��*��/ھ�aΘ-�f�H���oSp��[ݷ���:�'A����2�(n��[�nݵ�����2C��|�/	盦�<o��zG3E~$?��Е��0t��½/�I�gz���3C�Ⱦx4z�����@��x��"�k�?H,���:sW��|���3B�%-.ۊWB�.$��!��n�Ibop�x��1e��C���<f�Y��|�u��1/��w�8��^�fM����j���&���^��>���Dՠ9 W��a���rq�N��L�ņ~����Ek�kh���1��!m���wȺE�E�sz�9X�/���]j�� �7���KŮ��Y�����r��a��`�ـ�,��lV�W+�)�\��>�������?������?������?/:Q�+��$����W��w��o������a1��`67�-k����GC6��L����W1-'Zc-8�)I<��1@,Xy���;�V���ʮ�@_W��ky�h���I���>JK�.�G��O���_m���	�%�G�y���H,��a:7���j,�vti����t��������^�~��hh�S�Cin�To?��]�{h{�R����1�ߥ��F�9^��;T����s�����ByO��}.őI�B�Pc���:Db^N�������e.^�k1^��)*�M�]ޔ�
�CM�Iυ�!:NMo�ǌ��)��B}S��m�O��.�P�>ۗ�'PH��:��Y���r����к��.�3���zw����>�q�4��]>���0��'�_RZl3�E�����`�J;}����)��Yi�A�����oAe7��.r����O��zF-8^yJO�hJ�/�sw�7l�6E�>)������vbt��;6�iv�p�2��b�(��l(�Z�Zz�t��BC&���{�(I���곦/�ڦl�Yו�(�r0��ɢ���	�w�7�5_��3]?@/�ץ˄��N��bt����E5^�#�z��춃��^���oˬ���ͼ-�w���Q�6Q�l��v�v�lG���"�C��nj���/��7��[/֒9��;���/���8�5fa����od��m�UDe��#˔�Ō�Z(��kc��48u?f�2䇥�O����)��{<ݸ'�����~����aM�E헵�j��m�����_>�9'>��EH*�ݹ�ˌT�vɯ	������}o���Sp�`?m5D6"�u�T�h��C1C�ʻ-�ꄸ�p�ݨ{1H���N�����̋��}�%��>4��/�����2�d�oצ�����V�m�Y�����/������ƿ�{�b�X����8���_�ɟ��_���>�6�r�����f�K�h��Ό�� @I��bC@�`|�Z^*C^Ƥ�`���o	�8�"
����gz�:{ˬ��v�����~o��2t���tB�j�wy��nʴ���C�y��[LSSy�/D�q5d|�ɳ;��'7j)=�>�/Cwk���gh;xp ��2 tǇ�#�E���S�����'R��d�LQty��n�~�\��!y��髎b:1�\ӗ>�ХK�S�ө�g$�O����'�8��c�����	��6��J�[�BP@�'�,5� \�tu� ��v�L��ڸkJk}Ji�rFu@�7����0�L��<"�t��C�~y�{����>HS�_��6�G<y��.tE=��t�Gja���M�l'Ġk;��x���<K5�i4;���i����b6�D��x���7�Lu|vJ��o�1�|)fc4s�P�J�sx$��¢���΀A>3㣼{�?E�|�P��jy0�D��_�c�����4_�N�V7�e�ѩƀ*/�S����vyұO.S\8�?��n>/��]��9q��G��N�����-⎷������H~�>/���{�� �2�84r���j:���B�P׏}�<��&�Ч�ct��ʔ��FHGk*${�$��ű�8ƌ�l۪]�X<�;�w��LIs(ՃmAׇ���y�}� �x3�,6����4�m����h|�Bퟦ~�5:/�J>M�w춳�I-�+����VM;����O�w/Cw����T>��d8쳯��c�Q�+Z�ܷ�:�h�oӑ�6�B���}�a��~a�>�k��|��s٪�"R�X}��� 
0F?��[a,��M�-�mޜ<��ԏq;��v�����ļ���3sX�����,;������޷������_���-[k��Jุ�|��g��^m�)��f0�-`��!3s��4�0t��c��?�ƚx���X1�:CG���~l����4�~M�&P�<��@"5��u�m�KA��oS�M�!�,g�J���m����x[��>���O� v�n��`�B�����~��i2��f���\t�$�;~�R�_h�"�!~H�|�VM�t���me(c�ѥ�N��®�+���>� �|0����S���5="Ɏ��y)e������[j��=�Qv����`����SpIuw�������z����8&~L��R�Lu�ۥvG �hW	m��¢�-��FC�B��"�Z;���y��BP�}]��bϷe��U(	p��Z�(Ls?�f�W���ƺ|�wP�A�&���[Z����]� ������Y�f���&T��p�c�d۳��м-��?B���q6�l�ڼ	tW���:� �	�>�|��0dW�tФ��/cx���X��y��=$�Sa��y2\�4O��}lX��������vH�KwA�����.�x����uuD�~:�T>O�c�����%;���s$T޹�C�Ʋa9��i��ߤx�P��q�\J�ǈ�X��Hm�P?��:4o����QHf$z���k��)��ٔC�m����>��"���m�.��m<�3g�	>C�x~���*'�.����.J+Ze��m�D\�ۗ/�?NX�ŕ�����Yο���������O�����_���Oʢoq-���Փ���Ĺ=S%\�ּ�I�?̋���J�H˾�e�0�&mn�Ύn���4Щ��i��Z���@�b���s�x?�}X���AƋ�I	P��o>���D�!�m��4i�C&.��9�p���Oj-�.�^�Q�ڡѬ���zG��X_��e��s�$������Շ6��vm��Eo��'�=��g����^�����mD���K�;6O��o���η\B�*4��)���3�&褐�����E������y��mV��E�]��f6����g�2So��@ǥ���;���̝Sb�����-P7��]�62��T>6~}��ǈ � .�R�n[�lVNqȜ~�bP;:>FS���$�q�>�eSi��j�	���M����5���6���-j��(�z��8���`zy�/2�r6�{�L�!{�?/�[9[�װ�lj]��y�"�z9B�nWi|��/�?h_Vtj}�T[?�y��}Ry�'�w�vJϥؐ1?"4ߦ�����lO�Wcގ��w�~�G�z�[��4�_��8�1�v,��!i<����&��۾}����)�1���T�v���ژiz�㕮is�1cF��!}��<�~��7��(�]�B��KjC�/�ڥ�����A�kp���C�P\>O4	�-�{�M�M��A�Ch9��ug��xW������Cl,�>��ƯI�Ƅ�z<o�qtj���mȹ4^Q�cF���vK��f~�e۸�g�6hGȠUN��%���w���Z� ��P�EV�Wc����������������괼�`���vsxysy�E�'�Y��*fBv�:��5��P薲Z /�#S@rԥI�os+��ϛ�����<�g�u�ie8�1���Vi<y��)��-}^��4/�'Z;�~	9Y)c/���M�ͨ��k��3����>'=��$>�՟Ҏ�v���hLmG�=cȔ�1��Ƈ�BM�R�&�W�9���ϔgv>�o��	ƃ�6��񂤻5^�vM��@�t�&;X��fm�:��k��!:���]e*E�s�l����8x�k��o��0��e�7�;�����E�~����]@^,�X.JG`Y�.�/�a��qû$E�&��z|��K��氭7V�U���laS��E�ܵ#/��㰋<Ks��˴.�û�)�M�Y�}�(�h�>lS�_Nd���4;:�͎j�Rs��x�TF�YC��8N�?�����?�INFP��D�m�v����������r	V��_)k�K��c*�3��y�녏��O�r�V�_�7�.����V��뭓A��q����r2h� :�|�
�[w�����g��8�W�a%<)�+/#�/=���:�k)�H�'5n��h2�n{�!x4{����S��8$�"E>e��)�<�EI�9~�V��缞1�,�G�(S)���b��/�N���4��c�9^z�ޓ�1��%ސ��SZ;��h�uh<bc����{�vh~"׹):��'�5O=����O�u_���ͪ�I'h��B��+w���ݞ3᳃И���(�sM����qnt��=�I24ARdj_�鼇6~!��t5�Ξ�pjq*�>�9ޥ�A��1���>~��z��o��m^7��?�|��n�f3u�z%p����/+
[�V��F�'��$��)��:�V���V�V�Do��FC��P]�>x4�%x�A����4��k��P�4�UÝZFj+��O;B�����Rr�Sx:e�	9y!<�2�h����R�J��~ܧL��vPBG
�}�k��j8�t��m�u���	n���q�/M�b:G��R��]�[����P}��L��s�Թ3��$�kmv��\�?��e�d���<7.1�.���Y�E_��e38::�G��G�Xfn �=^�8��[��`i;2�{FѼ�\/q׼u����f�p}}]�]��6�6�v���0��0���w���ѱ+m}��O�1ME��_�M����1$�|J�IM�B�$��!&j�	�k�Q0��`ց�]0�*�fy�4:88���GpxxP���P��F�;q��ys�x�cR����x9�Hˉ=c�./.���ܸĩ(l2�l����F�9/��~4��>�[�_S��>��35"�^�L�,k��?��}��a��[q<�>�e4ۧ/τh�C�H�a̿���m�c�RB���݆��_%�#d�h���4�L���S�?���B�G��iW���#��Ԗ�n�ڑ�;E/��!H�o?'�����+�`[y"[
��Oʯ�4�������	���������n����Xh}��X¡�I*p�G�_�+�.�>I�Ƅ]}��u�M�}�9�!c~ ���h�(�g�������3��YmG�c_�+˘��ˣ�jubc� l+�
z%p��^6w}Q����A8s�GW���I%9j!ЌK����3O�RO}�ݱzwy~H�!�?Tg�#7�>���!��Ǹ���.���76/���/}`�]�l�?]��6��	n�5�ֱCt�]��@�ņ�},ݹ�n�>C�� Y���o�o6���n����������z[�-��3��uQ@�`�� w b��3�i���c������puu����Wnw<N���� ���i(h�ۤA��s�c~���_��Ks�%�G���SW 8���ʡ��D!#\�P���;�XvIHf�������a)cp�<*�d*���1�xQ��l�����ϢJ�2D�J���E�]��Ks��������֫5\�2v}u�l�[���ʃD�E�R�B@���[��{,�e�ѷޱ��]�-2���1���_�3�����0��K^S@���ů�c�?c�N_N��}���1^�Zj�}�c,=<��.Ls����B8-#��R����vj��%�e��B��������4?:�7�e���K�J���XΘ0�m4����_�yJk�����C|�[�!\Ɂ��6�d_�pdWWW��Q�^	�]sc�>��\�� |7��m(֐]'4�M0�>Aj�����x�2���&�X�>���jL�=��b�	&�`�	$��.�f�K��o�?~��<y���e���=�a�v�;`��bn��ǫX�칆t��	2�^S;�g�{vk�����)\_�������QV�%������|[���MvH��o���w�h	w]�/k�}>_���q)cO��h�:̬��݅&�'�dȿ�Y�{a�@���U�W��B�2u�U�&�TG�̳�8xt��V�7pvv�v��*1��ͳk�R��2˷7(���%֟c�1�.�`�	&�`�	&�;h���6�6��=d�a9��5)�O�i�� J���^����v�_�ÄT���Z�٥_��% ��)=��Hԧ�R�̾�-n�e�>�O)뀒LI	�P�A,	��O}��$$�Δ>	�y�M�p<u9r!�ǆ�|P�os}}���|��O�����?��U���D�"�`8�L�	�B�9Uq����3T��.��Pco<|� 9)L0�ܮ�Qk�Jsz��*o�ۅᣣG���c8>>��b�۷�m��s�J�k��#cG,`���yƯ$CF�9+�U�vݰ`�O�,�n��>���`yp '�Wp~~�v�(H}M_����P4���1�s������zN�/�d!v���8��%�������9<<�gϞ���ߡ�d��f��'V�gr��`�K1�6(y�|۝8�G�%kd�[R� �ٺ������cq[�5V��$�eپ�1_��d�GGp��>~��v��:PT�ش�j��U-���@㷾~�X�|�	&�`�	&���}H����Ɣ�.�]�˯��xȋ��o_�O�2�k�z�����g)�7b>l(i��D��W���i�c��|3�N)a��pp�tQ�ig-���u)�I�-a�B��B>���)�\-yCK4�W�ӭ�	�7�&>.T��Fv'�}8�*X��ϒ�u7�����gOq�-�;�#��pCp��	&�`�	&�`dLתCe�9ۯ�{ֈ?8X��/���S���v ���-�.���-Ȳ�����$��.��5���]1l҇]���[�6U=����1��\��]����?���6�*��՚����Q>{�\�d���fG\�N]�Rf;�k͡j}/L���a
�I�q�H���ٝ��$�K��w�kN�x�y���)��8?,��ٳgprr
���Yכ���ɀ�//��-m���I�K�(�a�Z����(��Y�$��	�A��r��Ţ��ÅK̚�#[J��嶥TY�|��ޱǕ:<�X�e>+�]�]9�`��|x������,��0XᏂ��}�	&�`�	&�`�O�Ej�A�V�%鳸�#ǥ%��h�x��b/:���c�����7^Ӟ�	��o��;�Q��.�GwՓ�(%�sѯ���I�3�)���{��}��~"��VN�ԯ<@��m�V�B,y%ַ|>�Oi�>����1���d*֯�����9���g��"�~��yQ�W��y���!I�8��S�P^���9��o�Z��f��ܧ�C�q�7[>f�9����.�@��<�GJc���)|���?��������3#�QȝC��BD�bP)fHLp�AS1��@�~��)��}hI�P}�	>}H��	&�`��� �54��+�~)7БX,�pzzO�>���CW~�^�gj�>so�{'b�ٖ+X�Vn� [�.$o7k��}2���;��])2���9fՑ-Kwl�|>�=f.i�=n�ɫ�y�[�-�r���C�����>��͍K���D4۪O��gH_J��������Z,�G%�-�n�E���6_�!�p���X���tJm2���ӓ8~t���'A�ċZFJ��,�W'l2�����֫u-c�����Q��.��%-5,E����J)��-���\,ay0/�~Q~.\R���]�V�δ�������ѣGp����Jz��S�6��x��P��~����d��a7�]�B�
)�ծx&�h�	>��|L0����M[�A�]*]K]\�ʧ<��iZceBq|�H�G$�6�Hj_,�=�φ�OSi�f�����$�,�b�kJ}�Pz>�Ե��o�m��^��y�&-���kw�{�{��x�_K�P��䈘��8S���!�	��b�~��X<D*��5�׶�s��HQ��8�;~� �@C�,�\���#|�m�T ���Z��o#*R&�	&�0�L0�� ��/�u\�vY���ÃCx��9<yr
�<�g���ެ�3s̮7��7����=\\����ecw͛*X���mN?��.<�����qpp ��G.�����Y���m�y�i��?Ϟ=�7o��۷o�vl\=�V�m$t��#9:2����=<0�k�l�����g�@�TPծ,]����uڱ��[W�Kt*��'�'�J{�6l���=V�ì����;ٜ}8s;���ܸ�
 ��>�x0�j^+谅J�]������N�� =:*��,�.�;��Y�3��<99����Ǖ;V���a�i����<)p���0�_��O��;��L�>�|�J �%L}�آfla�?�R6R[%�;e�>�d�z��-䦔���ph�Tg���m�9u�_���Z�i� R_�.FK0t�Z��O}�j���S4^��+S����9M�P8.΃�l�t��ī�Lq>�% �:(~�F����N7R� �5��8B:&�G�Sj'OB�ʄ���C�s��0�"q��acH�tC��~>(.`ܥi@ə���BFS!�_�D��K�#���6}Jꏱ�E��R�:v���3��	&��A�5˻���V�����������[�����8==����[����f`�Uv��`~ߝ}����������jN��v��h/�7P�_��B��Z�}�|~Ǎ"���k��^���,�s8>~O���ё���b��q��os �<{�������s_�j
h�:� �r�֩��z0`����!;�0��l�M(��>�Z�fu��`��ҡT���W_�b6wt��k����EdJv�r_�����s�ws��$�6~��f1a��ڀ�5��le��*�����K�4���S'k>٤�3 �b�۶-�K�#����%�\]]�{X�Ӡ���%v�i-�_����l�]��!�Y�g�	v��<|��Sm�L�y�e��?t��#����UC	|��>/��P�/�=����3Z}Z��F��8�Ĳ�"���G�՟��g�#Z�]�C�$�B����%@���Y3�ڠ�F��u))a#$�!�Z��i��i�ǥH�NuGH�hm���1��MT���7ۡ(�$d}�P�^_Eu�����)kC��I�`�	&�`�	&��!�f+��%�Įla�r�u��ɱǕ���1/^��GGGn�ؾE��.�9k���z�g~'�˫�ֹ�ym�g�b���>A=�.Cڀ��2vg��T;�#$�6+wlûw�������/�]5��v'���'O����ׯ_���Z�.<� �Gh]h�{�F����-x�>N��ܳi�ʞ�?���@{��|�p����^���\�ac!�M�U6���(��.e�Ç3�X��9��	P�=�e��C���\o�=M`�9����6ϫ㐪�����]�?8z?y�vY.���e��K�dŶ��'pP��~����J�䵬��eȪ��ry���R�L0�L0���d� -������!u��M�b��*������W������v�Q_���cjB���'�"b͜��v۾��CZr�)%��=z��i ��m�C++�l���'��P�$�R�B�c��u^��r�g�֘n�'xh %��cY)N#���w7ҭ�����Pҕ�+��+����_l	�ט��f���/����dp�����3�:����gA2^Bti�4�{H[5���q;p�9v]L0�P��F�\���"C���9h�zC��`�Jx��;�����wm���7�Y�����}���+��wĊ�YU�v�-(*'�Z	�w(�s�i��;���N_�u�2��nq���%m�n��'O����]`��7l�Dl
w�ʗ_~�9>���:������&*�}_]knEG�%qܯ#Tn�������8��7�1-j��_�QCv�g%>nw�Y��.�j�K�Ì/�����>�o��-0)�%�4)����$V5rN���J+�&#�a٬z��G��AX���������ɓ�ۆݑ|�ʡ=&fS��r��o�����[�+�Y;h&Ji0�=6��s]�W8��>�z,�p�	&�`�	&�`����}�PBڳt�/"�2v����C��""]��l�Ը���H��1�_��q� eA�>ٍ}��I{1�ң@H��>�%���2���74A�H}�% �������`���5�h!}��?1z�y��L��h�<�ƀ�q2�mu=�z���t��2�!!����6�p﹅#���P�S�>���C��o���G�h��}'g���c�=��)qg�	&�`����{.�U��)̃?Ƙz�֚����~��[��v~���� ���ŗ�����[����0��gd�ʈyK�"/Ą��ƀ�(U�)�E�pai���rg?�˗/���S��.)e��I)9�M9�N/�x�|x���p�^W��C���S��|�
/��b�&��1�����m}|�f���={O�?�Ң�q�F��Ѽ���k'gv�|����I�v���:�MM��Gb�'��T�y3���8�F�X�W���o�)������ɉ�f�Y��V%��-q}���~�>����|��ފ�v8O��0�6L0�L0��*�7�-�]T� ��)oǣ��]Pbgg�"?^���JS��4�����>����`0�$xL0�}ʻ|����mc}������s�4g������7��G�)}�%�I�!e�>C��K@k���f�p`����Y����P���%Ho��3R�}�b����P>�`�	&��au<ݧ�Q#/�9<{�^�x�7l���f�F�����-޽}�v��`�$��Իn�����Mi�������E�����Ii�9H���G�زv����+x������b^���9%� ����1����O�������	Ci�0�|jb�#d�����.|7���Q(�v���a���=� �志��=.�;�gߨ��d�`0�������GX��u�4/�.���7��Θ�+�C3ڟm�7�؋��nw���?���ͳgO�����V�U�G��W_��V�>�A�((�	K��2,��ӰkL0�L0�|
0V�[z97��=�_��Ҥi�NiqNN����
N������w{AYK	����Ч��gR�� ����!�k)��!>�����o�k���^�1�:B	"��}���K�� O
����D��'2�9�=4��֎s�^ l�[D�9�P��/i ��1����&ke��)�hh�0�9z?E	�k�̽гl���3����I�BJr	��3d�J�C�McO���;oW��$���@��6���wYd�L0������������/���6k�C�=Nen!��V�5���-�}��'H�]6r��40��P�D�b�E��9p�}굧�zU��HPЁ<l�j���e�<�LJ�1o޼������/����%�K�Gn�z�[���y�����~��[D�����P�`0�5;U�"V�;d��D:v�9l�Le?s�7�㽜�������[G�T|��U����ÃC�����{��;��O���`Q򠕧���N���D٬:���T�MD���Y�kڄ%}�΢~Ci��V� os�߿������7pv����+8:z����bemfw����/)6���(&��g��v�Ԡ>6�;�:��<җ�nI#v�V&��	��c�k>F<Ct@��ɷ�}u�����R����G�>���ġ&�`�1A[�t�m��U���<�.��2&Y�w�����N�tR^Z{��`�8��&]9�8�%x��ں�v/�W��O����31@��]�0~�vO�w���B�tT����u�GU�~�4UrT�`|C��i}�qb})Y7������B��-)�D�l���/-����AiKY�?4#Q�S6�k}�k�$�.�{,�aL��
�
̆�L~�TJ?߾Q�z�N"C�<�g�	&��>��K��1��~�p<�ötD?{/^�(��ܢ�f���E��ݝ��`��?�����[kԙ��sL��j��c棭�ۤ�-Z�y��a�>
;!��^w�i�?�G���gt��<^b;U��d��_�Ӂ�Ǫ�_�_��_�e~Ϟ>���(V�\�jK��x�䴼������W��\����B�݃�5�9Q_�����u���������$��Q�����
��+>�+�wI%/,�i�s��{t�M���o,�����û�������`%�&9�0��E���thv�)�ϩ/4���M������)�,��O��*Ϟ>������3جV�\/\RǗ_���]F2|C��3��Q��O��n���'Ә�\+j���]�M��$���I�sR���D
	7�/�V�/볠�o7�C�g��?:��ZI.�$���ƄP
��.O0��ZLjZ��M�E�Iz�Wj�+��(ަ�P��~��n{&^�|A�����T�_~�4}>$1"T6�����5B�;���e��Hqhm��,���o�Aa�܁�"3.���>�`s���@ n'�ѧC�>�6�;�.D_���~j��B,��w������X��P0�� %����^����zur�'�`��taz����s1�`���o���O��گW+W����ݳ��߾�g�a�Z׋��#k�WMВ8�o�0��;cl�����-���`��l�%��b���l���%��r��m�}�w)�G��]ʸ���mެ7��-\|���^����c�����lO�<�U���o��f�i���#�C^	و����j�$��s�}n�MiЄ�
8*��믿v���6����� ��9\]\���}�WW%n</#��v�D�p @�WRC
C6f�W<e>��D�����������3x����>�l�(�)w�^V.���/�ݻ���緰^]�	��	&NI��vG�u2W��	R�ox0K+��u�f\�>�]�K��8<�yM�X�@��D!���ݰoY���!�)LpA[������G݆$��̸o����,�!��m&���6�����L�o�s�d���5�_�uI뼘� I=�Ҙ1��+�%��5ccH"I}݌�b�!/�y��m�OH��Z㻝~��{boŞ�/�rXG��
$��3���z�6i��Pf�DGj�B�T�6f���&�Xp2�)��g��ؽ�p��8L�Lp���=�`ȱ���e�?V����&w;أ�r>����o������h�T����������s9�6/쾃n��ֳ]�.Q����s�/��߁���_���ǰ������S��?�C���w)i]k�đ����<��n��Ri��Ïo���%|��Wp����
puu]'����	�߾k��j��Oi!�iF�����KǦ��$ c�5���c�,�f3x��������9�6I(��c�KY;�����o����i�>�$'xQQ�#iL�F5�f�ÍM��>(��"�����r�&��o6���;���W��]����`�][���˗ϡ(u�O?�8��|[�
������3�'���ᴲ�/@�)���;)4k~D�M�=!��~�1�~����ǁ������B<���;�NJ�p�&�`�1���$_��\��#���ر�|s�o}렠�{)85[�a�w}`���)���=���M��L�������^F�r�TuM�ɡ6��;S�3��_��=�:6�}�Pq[z`�I�uz)�ٕCy��v�wq��0-��	��f�oؔ�Y��B�3��x5cOjz_
�r)�NSG�0eg~G���h��}�0�kY�3hYiL��� h(�.}J�I����?|Z:�C�Ap�u�I��?ܶ�E�M2rwп�9ۚ��i�{��9|��K7wl7אo�p�X²�����[T��6a�.�����A�ST��_h�sK��]�ď"/�ܭ}|���}�G����	�yV/R���O�������#��^�b1�m��l�d�����F��n�����.���ߗ׾�'O����%��X.�/�,�/�Çe�jN�}����l�����w��m�M�dP;s���s����4��)��p!�M�O����gϜ,mJ�;�X>;(��&o؝7�)P��$c�����N��Ed[���U�BQ�g�e�\�N�x����[����٭6r�����GGpxp����f����|���ޟ��Z}�U�L���%�N�|���7�����y�9��K�_D�+��XO
H:1����m���4��=�;4�h��0����zwBq�1�ޔ�^�m�Z(P�_�|�	>G���|̸��K�yv�H�q�x��
㵝��`�v��;e'7I^���@��}"�Վ�i0�>�O�|�&i�p/����/+�Yj4�9S�}��¦9:%8��J��|V�������dED��$y���<���7c�~ N���y�O�:�c-z�d\��
+�&<Hk�]/P� ֶ] )�')�P|�,�L���
��_h&��7�L�����w�1���qw ͯcѧ�.�����*�Ɓ_��a[��!8��$�f;���1���%�l����a�����.᷿����T�Y�G��b�V}�rx£Pp��j��o��������u�_����!��������%��3�n�}�lɾ��v�≥�r��.��~*����ɩ{�&pl�-=�/�����`}���T;+Ѕ�V}�,�0��_r��2񭩢͋�����X�2:�,<o���i�_y����?�7��(��G�pR��Ǐ�7�DF��c�$ j����d���JKT;蘚'�/����!��,0�~������W�r�3Y=��7�������ܔ�f��"ʫ�VӅ��S�����h]����S�mQ%�wM����L��[�)	�m���L{F듇g/�$������HeBq�1�~�����|�	>e@�6��O��^4���p����}B���n�U	��0�0�:\襉i�&Ѐ���'} -	��˜������4��Ni���^��̬ 3b��
��ܓQ��@�u�l |@4�ȑ
)�0�`�3���@��S���%Opޑ����JJ��R��.)��Lq�`��}A�z_��XROJ�\:�*������ӫ�lj���+S�AI�'9�� ���_��qa_��@*�k����h7�Ƃ&kH�i��I�ŗ��ѣ#����������C�����~��#��%|T��Q�SH�5S5���Uuz�&�v�ؔ�v�p��׿������~����������?��ptt������#�mST[p������k� rT��l���>f�<::�W����֫��vג�iؖt�ͬ��$x`���A��M����;�ݝK���H~ʇ��+���36[2v\-㖙q<��/����əM�9Z,���<�����.��Yc�j���gw��/x�0Y�O[�;\"�#��mPʟ����i"K� R�Qb���G�����o��e���`���u9������c���r�~����;�T�4@hhh�@�{��4��_�%��Md�`$�f��О�x�/��s��}B���i+���8�x0�~�u�!�+=Ӈ���P������7B�yػ�L0AL��ܶ~�uZ���}>d�y���`�>�I�r�s�XbD�>��~�O�����q#�d�)����?�~���/m����;W��!8`��I>9ǃe8��Z�͝ȪϪ> �:/}w��Sཔ@�ݿ�1�X�-�{BoiuH�Eiq�?
�jeB4��2I	����kܧ���{�#�>8���V���AJ�I���!-@M0����Pݡ�:B0���$IB��Mn�-%P�z���)<y���q�H1nQy�\�۟߸�UYV�E�:��`����eVM9���9��j7�_��̾�-{t��������_��D��I Ŭp4�ʼ�<��:H����>��-���K�/n7���K8>=�W��p;����O.yö�T-H�`��F�Md��ɻ�?ڢ���rKTE~����>��!l�X'��">a�~}��)|��l6X��n�	+c��w�~W�C���}[���,_v�h�D�P��֡��F����o�ٖ2�3��/_����ᴆb��ϟ�:�u)�`B����A�':-$��q��vװ���+�Zl#�G��O}&T.�I���1��5L��Gy�l�!t����d!�WN��6�O0��	}c/!<�mǕ���)�A�wߧ�b-A #�>7��ÐO�B(���K)�ŀ�EiIP�1�:9��]pJ}/A�x�����w>Gh˶�M�+���}|�&���$������ŷU�g��܅&�I�wM(�2�ֱ���=� ����)w�e��8 ����S�J���|N���a��,9�MrFs��u���1��?�o>���gOa�Z����K\�;a��������Yi��E�F�O�h��$!"�X��S�����|1��ӓ�\�p������ƿ�{�\,�ޙ���zA�T�%�E|땾��3�ge��g޽{�%���K���]|?8Z��/���X���h(��>'�?/��u\4�c�_n��x{0ܟٽ-�nL�Y��/�p�n�ʮ��|>��?�gg����*�v����hșo�x	ŏ0����/����x������Gw����X.ps�r;��r���3x��/Lk���Nj��r����(ZR��n�E�!��1�[�H�ׇ
}�ǆ�'�2��h���������J'����|sW>���N�֧S��>A�$�۳7����.?�AjRn������>\q<��eCr��d�!�!c���S�IzIML��ϡ������8%��e�?,=6v�<�qo����a
S��a����K4(Fˌ�F��sHƫ������a�kT8�/B�E(;�6�И�y�K
��vl�崺5a+k:����s�*�|$������D��1��L���������C^/��L� l��t��[�%h˥�r�jl����6�wB���ݚN�'�4��s����F9�M�+���,���}��x�$gp�Fk�ߴ�#�5������z��Ϙ�������[wԃ�1�&&�[�K�%��F�~�����­]���S�*lϼ|�%�l���>�w�(�M7WU=�2�2�Ё�87�����񣒾%l�(n.��*_}�5��/��M�L\���n�g���I���dá��ٝK�mq^gH�����y�����/Ak���i�N%(�!,C�ǂ��/_£�G.yc�Z�k����9�}����%o�ID�3v���G}*>BJ_���E�"_��|��D������"��j6���{88�d3�@e`�]������]���g���15�M�E;mj��;�B0�K��M�绁����H�/}q����oI� )~��e3�lz;"Uǥ�r���n��u[�}�1!gZ��8R�9��?��CS���yZz�6��!5�I�3�?���l��;7�K�p�	���&H�3�8l8�s[�G_O���K�KT������m�k��w�}��.�}<��Ǩ�S�q���Q�G�G��k�xM06첦�׶�\7�|�P�F�eh48�ڧ�qJ$p�8���Q��R�Щ��C
t��'z�L:�6<� �j̥ڊ�P�k�EHS�Ź����s��^���Z9�1��u�y])�Ҷc���〦�i�՗�)����
���e�7��P��tuD����`}���i�~��v;�~	�o���Ix�&Ct�,��T��~�Lx���5�+9��:Ne���۸��p@�BנG�Ǳ��o�n�����!|��װY簾ٸĈ�G��.������ٙ#�&o�6e����+���tJ�{�!ڮy���V���y�����vn����t������g���/6����_��_CVҸ�l��ZC�0���S���������W�V-2W߫���3��O{����ݓ%�m����&o�/l��O8��zo��eM��oQ=�4[�}{<ы/��-7�ꈢ�Cx��~��X��d�����D�N2�s��E�[��I��m;�����#��ۃ�2)6"�][<����s��o�u�(,���
V�,���_|������K�]�������{"}��]�*�]�F����nB�9��]��]ˎ}|>:_#����qmYeH�M&���q@���B��m��}ԝ�+*���k/��b�>�I>v��⊒�z׃cq�������{�L<�W�c���`H�pm�����A�����,�,R��=~m����ڵ�Cm�ϙW����-���5�h��&6�._�k���T~H}�����9-��,7˫W��	�&.���m ����%4tq<u�V
�p�T�� �<|K<E��2�"Xb�X�B,������@_����oP����N�w�쏕y{� e�f��I�k)�.hk��_�^�$l�;/W����]�����=ה�Wm����]���2�a��>wi���D*�7�R���k��;�M�ᑐ�~�����&d/�ԃ�h2��"��)���|�����`����� ���������bO��߰E�§'d��5vK��&�v`6�^�l��s6�UǛ5-��/�����D:O�����./.��/ʾ[��3������ŋ����\�_B�om�H��%��E�t�A�TGk���v����hڟ��A�Ⱥ��`�q�z�vB�Y�OB
��$
X���W_�c,��Wk8::r|��O?��'�][,ni���#�k+@w��veм����lP���	)`s�����?���_��w�1��z����5�<��_|���K��Ó��F�t ��Ϸ��"M�r�����f|��Zn�c�Ao?x5Ab� E˵y��|��m���R�veJ�T�O�ǊJ��šRbo��xo_-NOh|�Oy���mӿP�ol����)�����<����K|�s�X<L[�}����%}|�����s:i���T�����~쓂��ˤ�}v��Ħ'L�������"ro�;�!8>g^�=��x�Ơ$<w�kP)~�u�;�J������4�W��T���qq:h�&� 
��R�K�R��T�1l(@����R0|a-4iwq�渚�f��7�.F�m���>��P��w�s�χ!��<6��ij@|�ؤ��e�N��9~�P䎾61҉�>K�z�����0���Fg��x���0�1f��c��t�$L1��5�����������.j����� ��H��=��z�.��7�h������)��ܸ&�YK8?;�7o�0��g3�6
Y���j
�����k�.�5���ة�`+>G�q�����y�I*1e����ǧ0�-�{k���ٮay�t}yu~��1-�-��
��3�)���dW#&��]�l?�.j��'�=F�Q�`�p�(��a����p�<��s'k�'l���������dgHB����)�Lik��_O��$�~��ل�gO������m���<=��o�z[^��P���T�Xj��ȝfr<a\xo�m��ewt���`,�0R�ͺ�v"����2�����.����0f������K�I���cq|���V�F>�-���C��)4N��r�����lL�{����[��,��B~|�7%:n���:��ݘ�O��s��t�8�w	C�VR�z�	�@�G�=~-%��6u�F+B,	T��'Vp|�n�N�!m]-�=�
`���Bv8B�E����^�ӳ��v/��!�ۿ�@���s|�� ���@+�ԏ�-?�B�t�6D#��^N���1M�4�Q�t?�:��i�cJ��wASj F�8hB�1��D�4f1� ��O�MZ�]����s�φ���F�1 ������\��/�㆚�ל�B<�:n1���7��)�_�1ڥ���M��� �P�xGm*_�.���lf�����'ppp ����5��. �޾��M�ÀG�;B�L;�N��#vq���Jlߨw��#�k��+b��YC�C��3����޽{��]��zS�i�wO�>��~����&����ǒ�2���#��+����{���W�ڻ�� -߭��+�T?K�G����pxx�N����$)[�� S�Ǜ�?A^^�ǥ�f����1!6��nP�I�	U��xm>\�����o�����^o�\��hn���cDu��c�<��Ѷ%B�m��e��_9�ơm��u�<�_����;1�)�G��*'�a�L�}�P*��?D�:P�#��h��Pƛ��[�	�����y����Ƹ�I���C�(�m�}n���k���Ri�E�R�4~�ߧ��i�J��V7����Oֵ�v_WN�c�'j;��T?9E�h>�L0��7�v��;���X~*h��kC� %�{_*��%p6�[�þ�b��}�&�i��ؒ�/��y4c6d��g%��)��*�;}Nb\�@�m��	m���P�D��Rm��:�8�po@
F��V��a�����R�)x�>�'��O(-Z�aWz���)~ׂ �xku�R����!<Tg5ך{���4签�����}��'�$��A;�|�	�WXzѴ/�|�Gݚ|����:�2�=���>o�y���k�h�fi}��r��G��j��od�K�8��>�}t�{V%Zzb�Nk%6HC���|J��v�A_�t��1_��V}�M�I�K�x9�a���؝����>\�j�uD��>|t�����UW]wE�>������Yڵ�]@����>n�o��7$ pw��}��0�nݴ\u�z&s	v����k��a˹�WW.q�&nd��PZCK�_�i��6:9�[�m�M�i!{����h���;??w;q����VO��9<{����#l��EC[�����g���琤�鄐od�����c�,������Z[*��O*� �_g����5<)����in�k[��A�%�v���_�Le[�}�!��v~��}�����N��gx�z$]_9��1��J�D�4��s���K0T�Ry��[H���M���!U�R������lC~-$�!��l�H�%�t`]@g%=����M�A���Δlz��X}�O��.���n������4
c��4�Jt�k)eBύiӦ�WCp�6��}(�9?Ǟu���;X&4�<zVWi,Z<f���XB���ߐ���̯s[����DM��7�Ɋ,3ѭ��%pj�������,/�-���3CK�
�.�y
sk�����?�}���8��-��f�u���sz��''Ψ�¼�����Ul���~mw��ɨ)!��o��{����ៈ��L�gW���o�KFĀˍ��@޻�
9|�;� �9����t�()(2��QR��5.5�y]R�V/�∿�ş�%r[WgO=���2��?z}8`�`�-����H�6�g7p��	A���_�Wz�;J�xq�y�ZZ��RmMp�tv*\�J8S#MOH��t�L����E�tgu����}yZ��}�8��)�sج�~n��`V����{��Q��::�3�Mh;�G�;6��*ӾM�nWCӶ�V��UN�^Q�m[�g�A�w�0�J�6e�g��̕q�nlɪh�oml��qY�;� \]\����W�`c�~�Jt��������wۺm�چI�T7Ĝ��dj-=+�C?��C�z���~��|�q��݁����;�z.d�Q{_jK��j�?ǖ"O��ږ�䃼d���C����?�X�η���W�
b?s��x�O@y=�2�G�Ub���1B|D<F�Gj�|���<�W����p|���/�{ɢ�M�0_����K��`�����8t�<�/�|궍`�ƣ�t����)���oC~�D3�[��WLֵχ�����'�ʉf/��Z�H��3Zy͖����vݘ@u�D�f��q��_�>�,�)>��T��	�I���SA�#d�r�����ޢ��5���=<>�}�w@�}��5$�@����z\o�>�[�ߗ�vJq��~�j����/͑�9$�_BuS^Ҟ�b)�*K����_C�ޮ���kb�C�+TN�_��M����
v�m�\�b���A�<��K�/Bt�hIi�f/IOJ�N���ؘ��!���p��Bs��1��XH�4!�N�}����>u�h���!VW�~N�w4��.�N��L�Z+�خb�鬵�h�^
ѯAhL5���NNი���gp��ָX���;�XF�=��P1ͿkQ�,�?��y��1�\���P�^�w��H8~����Τ�YS�K���~���r7��mw	ԩ����� ��d���%Or)&�����}��]�� �z����Y��L�a�t��[�ű`I
��Kx��������o�e;TW���� ��x���^���l�E)�̷)<��UH>d����Q��>�F*�>ts�"��4_�丏������8z	'�g�}���ia�X��>l n�Y;���p}s?~��Y�YΉ���hh��}Pݓc3�I��s|[���@ ��F�xsܸ�������W5��h�}b��k�1�����z���_�{��1��r{�Tu*�m���[�#ΐӝ�X��I1����\�^����o�wA~�htK�C
`2���������ae�Yty���x��]Z;��m-[�]@9ͫ*�Vum۩��D����\]ݸ�Tf�*Q���ٳgpQ��v����&�M��ۘߤz%�:����c7;-R����C n�ǐ�,�q4�A��pH���9V|^
��]ڼ��!W;��њ����6p?��i��El��=ڍQ�b1����'��6��"�s[(.�����B_�ӈ��"����U}u�d�I�km	�>��M��^����Ը�X��}p���+�H��"��80T�=Bi���)�5�k݆�%��X9)�d_Z�<�
|ަ����	kg�.��f�He8�R{�Bh���m
C�L�CS��[_
�>Ϩq��/�Ծ�w�~��e9o�O�h5,�N� |���iv���oI��yM�[��H��t�&���}$p�׵��1��ŀ	sð�AU�m0����D&Ry���]`w���[�VMS�نf^/uT�r6�����C���[1��uo���i,�3�f~�\�݉16Jʹ����I|)��S�ƌ]n����T\��>�0�E�A�P�@�#0VX>6���%~M�!K��� ��qT���c�������C!�����~.ڸw���N��ԏ�Õ@�X�	��c�ȇ'��L��:�<$]�}.���o�ѱ��5�C��~�s.��X�Wr.��K�b������V77�MKܕ���wpyy	����g�U�˴l�ƶ���.����.�ozVT�2�z��}�A{(�{ ��w�PwNv�}h��36c��ˑ5�8f���.�_^^����z�IQ��ѣ#׷�5�"�w�2R�@��s'��*{\.��)�,����ю5�X�TW^��]{�۳����<�:>���dwlq�U���w(g3Gc6�Z��Q����Eܗ��&���g��
�-�|�� $��e�"]]��U]3pS���+89=t�3���Mc������is|R���t�d�y�ni��9s�����
�>��<}�pi~�Ŗ�}�q�%n�O�}�LZ׉tw&Jwc�8,��;{*vĕﴅ�[�� i�R�F��C1
�y-�����a^>DS�͐>��_��]|�ɯo��������bp	��NE�6��	�<�>/��6g��ג��4���>�=7ħ꫓%����1�3nO
1YJG�G�e�. �wN���}��]��a_��O� �&�C��Ɨ��۵t߭}_�QI�8��o����ٳ) ����^�*����J��'����'������pK~��#H;MI�hs:B��L��+m��]n���dX�1c��/��!Y��r]��|�]�P�h����C�~MR�����cC��ݵQ����љJcS_�f�C����^zc����l�u�8���90�>4�-ee��_��o�I�@r���5d�4e�:ڪ+j�c�|A�+x_5�=���Vglr�2�j ���Ж(�Ս�Z�
A��D��J��S�)���xH�XY�S���ӷ^q(�$_U�X��*�
��9B�h��X
��w��N谛�0U�x\r,��p�6ߥ�ZF�2Ou�t�@����D��7�1ƀh�#�9��b�jz�6x#V�4���)^���vRP�-���O��9=�]OR1.��ɓ'��g[f��;���
0�ς�10����������\^3�O
q�z^�t��&ѳҏ�>l�=d������-B�U�G��S[�(Zo��x���M�x��-|u�e����gϟ���MYfS�g�*'�2� &�)r��Gz�x4��?�ݽ^@k�~�ƥ��;u㼎������<>>��������f��w��U	v�>��|��� 'i5[�y-;�8���c����t��b��I^�P�詥<�uIQ!0u�����kj�xl����<}z�������'O���ō;��'la�~غ<��Ѧ#�41�z5��i-�h �1���~L�4�t�EynK��%{��;}}l͡�i4�-���bv ���m�ᕆ�ُ�v�/ئ��Y���}jvrUv��m��"ɿ_��OA�����B�R����C�v�۫ݱi,:�eCtIm�2�K}}�XPy�;�)c�:'�6����yQҙ!�$Yݧ �[�r�ˇ��t.��2'��WT���I����C�6�C�T_ C�9�/J��K}�"$G���Oۋ��#�-��.� ���R}��R����i����4�7/V+z��F��(0������@�d������(��H�s��k_��~Z�S�^��c~�~}���m<*��׎|җ�N�O����C�U�Z�rܭr6�^��L\7I�sHy~����I}���p���Y������	��#T
l2�j*n�5�3Z7�:>>ň���]gcAȰ����~ܺꀗ��Ȼ�>uE��B,9m\Ռ���P��F���O�/b���6h��:Y�{]�8����~�7�>�++���[�%��Y�q�*%Z����Y}���#2�$�1�{)o8h�2���q�u��$:8.�������ӌ��ܝkv�B�t( ы�Bo�ǌA��?u"�tv�c$�_�Fyg�ށ�"�H���M�H58�8i|,5}�b,h��<q�+�)}�أ��:xD�QZ&NV�ԏ��`	��Lx������pr���1\�^Km����2�~���x񺧿2,k��,�B"�k9��ڶ[��A�\k�tx||۵=֡�_�],p����`�y$���6�©4�a���֦�5��f��S�FV�������E^�R�z�b��YQ�`sw�"Z:�Jx�~�Z��V;��qe][Gs�i��R5L��,=�jl28��NOO����ڿe�ӧO��7p}�u;�x��Ӌư�_�� n�:B65�_�7�Ð�����4|)t�N4��-]����2����6� <~n�DK�C��3��R�b>���������I���f�0�Sly˷�����b~H��5?��e��y[�.|VW�j�)�
��@$�j�k�����-Y��� ��{=_a}M�GW�^0�W;��#\����?���덟���M��-W5I��6{�?�n�;~�R���w'��A�{����vħ��)4��r��#>�+��Po��ޖ]�]R���{�]�Ec
/�9�}x�>/�,����k?+��5��<S���L��B�œ1���5���J4J>�f�q����9/6w����ߕ�P�|��}����3�ߤ����F^�|��:�-H�N�^n� ��k���v��8ͱ��V�}��&���)�	�M�����$���K%�,ٱ�����qh�I�>M\'=�86P� ���}��ꟾ�W���#�!�Mqq�qLZ�BH���C�N��S����> ��'�O�)�Bt�95�kS�`mC�Ӏ�P���TU�-k��?�+=P�����֝��z������tն,i�{����P�Lw����mW�C�2)|��B�7���@���hy=X�UEF��o �d�p�9WjWH�;� *>�e��v%��j�����%�F�kب��/��`�n����È��oƄ�}��r��'N��8n�jG:Ըp���pe�92����O'P_�/M $'�;u���&	a��"9�"=��1���T��'S&0����"(�y��g[�7�ς�(�j�J��4�i�}���t��E���s��N�F[������5^�;C�/��M�/K�l��5c����F�����4�s:ekc1>'H	�:M��j�?`��h�h�}�<G����$ӱ2��W����C�/�ʨV7�}���U���q�����V����u������Y���z��]��[<��~��&L�g3����Y;�e�Թi�a�P-�z��N��s|��H���v�kS�/L�*[~6	#�YIT��!�����ض��ik����*lC��n!�;��v.Z���M���[ןU?�&�D��;B��[��x"6@�Gw�g\����6�l0�A������I�ā�N�W-�-���a[�������/���=H��<;z��b�2���s#з)�9�����}�Xr;�aў��]�pI٭�c����q�,���A�sV��z������	�c�����;:z�7k��M8����Ϛ���MueK���O��6aL!���lɧ�m�v2N�ŀ=.�|�
�1�s�x����:4��.�xM��9~,�R=��f��-�N_#������E�O�a�a��3�W�2i�;a�OD��~�Fg���ʛ����4Vc�Q�6Iv)���+O+������o��3)���H�gH���6!�:s?d��>��G矔q�~K�4�!�pj��t ��":�L}J�
v��c#z�H-�w� �8�.� �n��Md�l�����$����˳dҲ!�?�8(��[���+���[�P=��^�� ��[��9�hVu�[�@�N� mA?�3�\��o�-H#-S�K�ר�ʏ��П�i!���x�'4��>�xU�#�4���%��Q$�o�~����i��)T�Ch�K�o��	o�t��O�5�:��2�$��t�ԖN&o /�z��rzC�0�;)�-6�c���^�t�I����0�_�%pD�Az���a'��[�@��Ծ��������gM�� � �^��|̠ײ��s� P�-M�)�*��hT���Yi'����BwT�ه����+�����2�7��T�T�t��f�h��5�?�2Es���B���	�_C
Q*��X*oȸ�=\�+Z�Z�+��ޭ#d��(�n���� R&����E�� ���N}ּ�:�RV���g���p�Z�]����@���gȱ��FV����F
1:5#�r�Ai�������ϰ\���*��5�$��UaY�������Ql�.3��DY�.�z��z3K"����fl�j���Ƣh��*�lr'�a��n���
Гd�
&ux��p�en'f[��3Ȫݗd��������ox���y��]^]��T��m�]D^f�K�h�/�(�Qh{���`��L~F((�ʝ>f?;z��ہ��}#d��R_p#b| �.���k��V�%��v�j�,�.���O{,Ѽ䏳�s���j������ѕ�������_O�}ߟ������Ͻ� x+�:Z��|C}tfcCl�d��0)Ђv��/�`vzz��VGd>Q������t(ܚ�B�1���+�u �Ύ5�'&e1%�g��I�5d�]D���@�TFڝ0%�H���>�j�y4�Sq�'����s��|g}�Rh�e�����xr�����W�Ew��U�����X��Kk���פ=۪��A��!��͒�Kh^�6�J>F�����i)q����=>ٷ��[����%���~���o��9�m�TV�Iq�X�Nï��*�1����!G�eR���R'2 '(����=Ƃ�Ⱦt�dg��)6����奝¤� �R�v�l	�F�����gH�~��I�K���}��-�*��V�(���+�r�a�`Ҏ`�~0�c�����.���\ˮ<@�����_����>�u�5�^�^����4mC�^��_<�����D�BSeU�{R���A�Y��5��v����gZ�I:��{�i�W��ɞf#Ӿa��)b��fo���>�Si�ts��[#}w�h�� ��g��ЕIp�N�(��~K�(���kàQ�����lum�p�v�=$ �@r�R�c)A~�+q�����,���*װT�g�|1!���k��-�hSy6��2-x�XUc|SY���l����s#�|cc\��{���Tt�͝@
R}2�������9�����1�7�h��g9m�xH��d�HD,�¯��F���[���Ҥѡ��ǚo۴�9/�����i.H�B�W��'�h�w�>�u��;e>"�R�~�ז>�ͷ��m���S=��"7�s���[���4�"��|�GR�����r�Wb�阁����]*t>��!*�3g����gs888pG���/`�Z�j�3������İ$S|���>���|K ��X��9���W�GkH�<�VT� l�9{��Uu��-G?aG�e;�_�-+�Lu��z������o�B�m���[�o�%\H�{���t��`��%�?eE��8�-�x@'E[����hO w�ôlQ'��+����hA�Ol�VP���G����f�8�U��P�<������$�d��Y��Isܱӳ�u� F���Rq�~\u����9�r<�]�/���Ņ��d�(e
6������j�:NgcUc[%�q�t=��I۫���������7#�T<1��I䫬�_@�T�պet�%�SAcs����!�e(��a��3����x�ku��b��"���%�uN�lu���)\�o�BQc*��t�Um1�	��{�p�v9B?:k�pp�HF�7jm�y�ގ��d�ct�R\����I�(� �»û�ޕ�W�O��6H�j1�?�K+��N��b0��ַ.M��@+-������������]<���z�^#��r��DWS�r5f?ι��M������B�Hϧ�)�ϔ>�$l(�K�^���i�3?tl:��[u �l�oX��ܽ{���q�����s4�F�gdlK��F�,�`��	��@\�@a������4ec Q��<*�B�IURE��!�E �D��oK�e�F���F�H��{�c�ʷ����k}��{�3W��9w��=ֳ�ݫW�.�J}������V�m����KǗ\k�m[=��O��|u|/��vz�A���;�~C]�I�wX"��c-�Cb�t���©ޙs�5�d�z^c���M�z/nY���Y�t����Cm�w���Z������߃a�c��{��9�t��&W$01C�J�}��!�f�lh���ެX; >�^�(�g�a2Ú�7�p��N���HM�֘�z�w׌O�vJ���%�K�	6���z[J?B�����kB�)�ə������~VZtά�Yq`�)����. �F�P��$�gЯ������3=�cM������isXaB={`0�gy�*���z�e?�q��x�W"�=��߄���Rn�a��v^��Eה �_��X�ZۥD�YI�o����xׁ�5����w�V�^~:&���Sm� o2�������$��g�0ƅ7͖�,tp����#��r�64R���x=Ku�_�>,嘣�nB_�W9��}J����;�=?�nY��銵iiUq(��R�q#� ���cP�/�;u����E�3d7F��Kݒ��(��^��˞�x�9�`Jȋ�q�u����Q�e3f�*�A�_�N=��ZF�"׎�9������9��v�Q�urzJ�ggt��]j1�b���#a��辔�~a4��?��w�zz��h���ak\��;�@���+����Ϻv��e�����,�1���E���=yf�����V�`�`5gEɾ�p�s�'g�3��~+W�&}`�,�serLRǂ���q:'��q�o��%��iƓq7�i	����\iZ�cJ2o�<i��iM�Bq�n��}^�[0962c�en��J[�Y(�������v�r�sz\tY!���W�^��4@8�|n8#����d?�ǒ�5�š�:�cp˗b�w=�g����1`>����p��y���8��g}����ւt{�^�}SC���b�l��F�5�$�Q�U�/y��@� ��Vu��@���L�/�O�7d���(.R8n�\03����rP��5��l�����_�_?T�ut��g� �K?:Vθ��E��niz[�ב�U��b)S�Z[Rm_�j�r�|:Q�ت]�yZiگ� �#
2@�춰="������u�>;v�liT��������d�C�c��J�ý��C��k���ғy�=B��s���'���������w�6�>�L&U+~)��!�cCԯ�oYVnȽ!����s?(Wǃۆ�_��+���G�����F�>��8��>6A��}��8�������p�x3Tz[������.��k2P������W����R�è,��.��}�pD*x� �����T�@��OOǢm�?m�`:��!�>V&]���{�T����wO�?V˵8RgO3R�3mK!�	�@hL�x� \��x�t� l>�4`�B�9��g+�Tj	�#��)��Q"�FZ�  ��)�2t��n6cv�&{Xw��N�L���ފ�Y
)"M��F�b`��.���^�^
뢍�$+��l}�;��u��W4z�g	���	4-��%9��v���I��n��1�NV�flY(eđ��w&i���:�w��Z(�C����[�Ȋ�`љͧ�jf&�ߋ���F}�e R'vI�.7�;^7�k^"EJ6�~ }P���S�L�0V�o�'���Y��FZA!*����^e�4�<��@�j���F��%����K��+�~(-���@��8ϔlg�8���e�4$�]�#`��1N�wb���.�u\��Jؠlku�t�fM+B�����tV�}J�z'������IH��$6j	m��C-�ol�Z%�n����&�S̗
�X;����1V��-�����5��3�6�Ҷ���!�E[��X���s|�ҙ��
�r)�qchhZ�{���I����6��q7����ݎ���瞫d�hT�_�F�@'���N3�L&��a�B�-tz�G���n~u�sWg:���%~��aL���ؗ�/�x�+*G����X�*s3m:<������5��8(!�dF����ҋ}1�)q�滛�w�=okBIq�����̴�&oD-�q��đSFp�(㐯YS�*�����kQ�e�����J����(�U�X���ʵ���k��Y^�xǸR	j�*~�}��"�[�ӓ-m���9�{����₟k����:<e����`e�o��T>7z���*�Wk�liL��B`~�Mu��~m2Ř\`?H)}�<ȼ�V�'�^�Ӄ������������u�p�t�IǺv\d�O��7���9T6�elх0�^[��u�kQǩfX,Z��s�f�����ʛCG	r?�/s�4���=9��j|���)R2\Ļc�Oc&x��ׄy�C�u��R�J���Q��@�0�Я9�Gy�����n����S��2w�yѡ|^�Z��<=O9���?b��H2n1�2�����%+��5XE�2�KU��}�W�By9�o��wǔ�M,��t��������d����v�0��4d�>&��,��)�+{3
f���wЩ�Ȕ��e6��V�H�e����u���<����O�Έǽ�����(�~��v�k���n�!}�����!��>�+�����1��2~ۗe�#Ʈ��(f�l�����;���֑^��e�|�K8��E~_f�z�����4��D	��l���$%p��zZ֖ct�c�@Y��cۊzB��P��ջ�o-���ֶS�tJ]� ��7�c��\��c����������Xs����0QKD'KI|T��ڏ���Y��+��.��#��"�Ǳ���'�8��C�.7��v\)�ߝn���wb?����i`�ÑC��}׫OO����u�.a�9��8�����7�yk�7C0%8o#[��0�s7����T��`20����c�F�#�λ�c�\������unZt�C������2�q�kph��M��G�c��Y:>�7����m�qeY��EǕ5��'X��uL�Gv��G<��Fj����R�H��^��ar�w����U���k3R&_Ec�*�D�T0�C0�ƱR'*40!��К�����e�f�0𧊈j���l���V&�s�y�b�ayʭ!�~���~��刕�c5�#������ܐ��E\s�OX�	��Շ����X�$�8X���}��c0��HQ?�u^�ޖ	���05��d�^��sj�8��/�^<VHƛ��";��*�Q��2��Ni���d�1�9�z�X=uDl�#��C'���m����{~�)Fk}vxm��
���/ǡ٢�m߯�T��f�o��Z��m
��1�x�BV2���i�U���甊8^��&�� �OG:@�����?����5%ֱf8݇=�j_�w�E��"�$��|N��u[Q�o�x}�_�����f|��aP�ed#z9��X��j�$�q���}21�e�uRT�JG�՝��rm���%\�<��ˋ�]�Wt�)�h����
v�'�;[�l�5��1��g��cHR�i���[����v�O��Ws��d�v+8_B�ڵ��>�N����	�E��K�p�w���cMu�d5�L>�W�|sX��[�|̙2��&�튙���c���a���\�rS�Z�g͠�T�������<�PF���ߠ�r�hc�Y��v��R�e�o�A�n��'<��:��"�����0�Sd�~E9�����Bpk�1�v�Q�;\�֒�0����p����z��uZQ/���׫��D��=�f/��'�W}}m��eɢ�*��G�La\q��5yϫ��lDGh�LZ� 9�|6�䨷��T��:!͜e4!<������*�1hE��t�j.ІA��I�g�>��dD~�߃����@-�bl������d}}�~�� 9��0��XD�</:*Z��q7���s�U�kv�RC�u���;�+9���<��f������?V�9�̍�v��S�V���kr�j)f��`���J_#�7��c�����k��nɓ��zm����E��.�8h�b��R�s݌mM�Z�m����Y�}��C׺}��L�l�V���rл�r[g�3�'���u��Biz0ܗ��(2
>p3���)ס��)/�aa�׿6(��m]����W[O�ߵy��x�[��m��hDd���ѩ���|ae����skuGy2��ڼ�Ӹ�ضn�UZ����z����V�����=Ϸ������U����!�|��L}��)yOcvB�V�봯��	���<�Z+�������ddQA��,�����h�+��m��ͼ�߯�KQ.x!�V��D��A���[�ջn;����s3����f9B�T?��E���	��~oMrk:}H"�>d����U�]�\�[�dM))0EFv�;0��nO"G((cB4b���c@��/�Oy/,M=� �TBG�@��E�e�d��H��bm(���u��V�(��0�Cߒ��Q�'�VR��5����+_��M{������J�t>�&Z��~ �nbm��0��4F�}`?��C��w�8�9�l�a�v�v�+(�s���9Ө���N�@�hI-��\����`�H@ǒ^d���D��X_�i��C_}����7^�8��x�{(����2��P��.��Z�S��u,���
Y�bY#�SX�jg-�=��e��*���3��(��q��Ou|',Y��K�&p�]�����8v9#�K��X�c�6q]^��|<�:
V���0�p"٥�����xWw)K��{�+��R����	'/>U�e0���}������31cH/�E�����/���k�\����ad�h�\o纮�0Na�|ޓ�w�^��R����!�����?O���,ԁ�Vy#���F��q283��c���d>�+�WW#�v�<�|�Kik%KH	�0�;�Ұ�]�^]�(�Jۓ�G���I)�2���&�ϛ$N���+�_p`��y�.�>^�_Н�w�������~|�IX��MJ�����dx	���#[�J�	��lfAT��b����ӛ�5�ź� _� +ϯ�k��@W��]�[d���;��n����U�j���S�7���AB��4������,kv�`Ye������0Ig�{���dAC	AD��2 �o��z�]�=����-	�Y	Ғ �O�n乺��i�Yq��:�l#c	�)c�-����tw�]c�V:t��J�����CQ� l>��׼�v^&:%�M��c-{/Ё
�Wd������� �?�y�n��y.�����4`fc0��i�؅qY����خ: =۳>�5�m�|�\wO�4�L�
�ϖ9�E9�Eԋ�gf�x\g	�T���KWnL��V�Ֆ]4x��Gyj�e���z��'S����0�-S}O��>�`���3:����Xy�[]��c���[.'��A3`� �ƺ{��>�V��i�w���"�,e��_�Ƀ�j��-�Q��9�	oS+��DJ/"?p�'��ڶAA���S���)�^(���}�!c!2Ǽ��k])�X��bƉHǦf\y�Ǟ>�Y��4p��ANO_;�-�#7g\�7�I�y��ʌ���Cv�9V������\�b|C�{4��/�Y����RZg���*=;A��ܤ�ױ���E܉}k�l�<�~��U��&��kr�M�w��Ӕc�Ti�M�~/����3�O���ϋ�w��߬|!�����tY��X��ڛu<Dc�h|�{��k�;ׇ'���._�vlUoR���>�5��^&��;�ݤ�2�7Y-7���Y�����y5//ݘn������l�Ϭ�X�N�[�e=m�j���b�\�����ɸV G��W��kU�7m��6�N�ɐ�p /�T�MD�K�8����ϴߞ�nhZ��{>^2Zº_s&`O�o����K��8�`��#F�BmL.`�h<�D�
C���ڸ�(}l\'�*U';?�u�p�(��Ka�3y�N�-Y�KY�R��f�9gP2���U�2v���z{�K�ر�v� W�&�(��ٲP�t��1�-�(���?#N���Z�)g�gqz�|kj�8�^�%[g�&��G���6��2�R�f�=�w`0&	�ؕ�F��mo��pT�N�f����Y�SJqW��k��P38!�0��7
���d��v|EE7Εσ+�X�w�^CZ��Ϭk�F:T��dĽ���k6VL�G4>
\)�+��8'6�)�7F�}�ܸ���j���G��U������"�@)�B�g�X_d��L8L}��6���!�jV�j\�G�Y�\�-�`��ޮ��P��D�:����O���\�-�*r���ȷ�Z��k��E��X,���h��,���B�?;U���qgB��]�:0x�B�F� >�EjZ�2�-a�'PO{�3Yĩ�јznܨ
:��o���%��g�p� �xDJ���W�q���)���3�c��}�qx�^q�j�.o=����\��D�����E���=&F2WE~+!�;�	Y�J�c����q挑���x>�'g*(���~Hy��]����?G��v�c�����o� J�A��9�Uq��<R�� �j_����{D�>d�D���h{����s�W�y<S�H�D˟!�T�&ռ��=<�:J�XӒ�J�X�
��G���LVo_(đ�&�K��j���׾����7*g|�4Oօ(_*w��r����	�:;���]���{����U~ry����C�Zx��D���#m,0��>r���MP���a� k_ ��n�kPo�1L�vɄ����t(*|�'�1�9@Kz{bV#펴\h�H���������%m
����f�)c�ĭ,WՔG���c�\��g�Ӣ�J&��[qe�{�_:��s�9(5��Sx����r_%{L�%Foō�A��D��W��Pͧ�x��1}�`��絮�TI	�2�5گz��V��z!m���/&2~��tU�ϳ��r3�U왍d��q9�43�-`w6 ��GIw���y%	�� C|v�h�Hm���v#�]?(�;}V��p�ק淼���j9'k }mn��=>�a����������R��{r��a�o� ��uz��])�d�Q�q�s�h9A���G��>U�u���G���Gg�������]�/�=F�_ϔ#�v�T��MnO��n�4��c��I"���`����}Kcz��ށk%�Yd<R�����:��T?�����G�?�xQ����}�u, �~�0u���c�^�U�A69���9��v7'��� �}���UrC�43N�!GT������ϵ��M�E|�LD��ҳ!�j*q-����.-M/�Go�Lԓ1Es��.�44kӷ�\k$�{��kն?z��}mu�5г���֣mo�߱h;2~��D�v��g�%��ʀ�?m�������Ϛ�����%����奩�3�a�p��K�5���zm��7Ў���vc=fs`{���q/���
f5iNtưZ��X�ɰ�q�،͇JO�\{�?���oU���_S5f0�+�^�nӟ���>]/�C��e�%l�?��J�@UxC�{r����!'A�sE���1Lv��D�bL�|�
A[mj����B���.�#ir���~*����X�2�J�]6#O3*Ga6<)������).ф��Yz�9��N#Y�I�*Ł�PP��k��N�#Q@��^^�������*AZgb6�A]����@!�k��}�c�i�F ĉ��kK'A������%C�
��Y�"��,�F���!ɍ�I5��������
��������^���s�Ԡ�kp5��c��P��Ɗ60�D�	��P�&���g�'��֗�^�	��A3��`�'�!�x�]����G�S�Vu��h0C��ݖ��
}ȼ��i����t;S4��[17;vĉpU�����۰E7����QY�5fS�s�,�J!�C��+	#hn��@�S�y�9��Ľ���M�p���t�)0�~�ޢ�B���\&7RF:���ݶ�5e�ӯ�k�Qٱ�W��#-Ʊ*h�C;?'�*��%;�$�t�`I�:1�L|�|=�K��M��p"���
��Ǆ������i��4e���G�>	dt�阿������>w�y��gb�Ei_����#�4�f��z��,�*�9�L��d�, 	]�=��w��w'����Iq��.���]�G忻��3\$��6ܖp}	�)G����J�����t��؁�I*m�%�vEK��q��Q���
|���җ}�hEb�/���$���%=r��}���wO�N�l88G����2���%��27''��n�9|���%��no�vX)k��ݮ��k���0/���؏��������aMY�}���E޴����]��Tm�@p����@�?��AnΊ�F;���Ery��g�J�S�A���7(�[�2I�C�׻]^���s>�p3��ՌU�A�Kr�1�*��f�f/���;w��g��DZ�[��"� �\��)2p���Ms�}'#`�Qϝ� �?��;�q�"gу������l�vr�;���1Ľ��nϪ�EȞ�vӎ������Ǵ�8X���Jf;���o�T	��'r%��]�'԰�M(U�-��N-��j�E� |��e]�s�1�OFbZ35�Js�4�C�AŒε��c�C�&?��E��꫓:L�O4��2�=%��@U�(:��y�)&��u6�Qƿ��r�?��z>��'wֆ>]�����@.32���G���X�|Z�y�̺��;r�aJ�K��01Yu��������+]�8�X�D/����� �UjƖ����G𼞽��tͳ��������R���}����X�J/�+���`ŊF�;F�ý�j��n%�֡m�$L �v�ko/Q.���Q;�<q��ME�-<Dm9y��Xd�M�1|�'����Gzmj���4
2��%�Ej�����!c���ً"L����1|��%�/�l�I@x`c�Ϥ��(������`
���&�c%h}Eo*h�����0t�O��L�L��}iE6\IoJ�c͆;8��[ud���Ɂ�6�����Ų��&��X!g���������[��p��kU\	X�/k<da{Q!��v��Y����>[}��5� �~��*��k���k�ᄓ�[���&�J· ����^����)�O˹�O}4����Z�w�9X�\��u�Hg��x�����O����}��r�2��]w;�U�x��\]��[z�� m�s��[��nd�n ;��|S�����.jz���z/��+m]c��M���(�rQ��\۰�B|ʎ܊~2�(�54�z�ד�\_��a�}�ݳ��_�1فZY�7�,��&�����Cq�n��x�Ǳ|n?l^7���H�	:@�6�@j�u+J���>��|�y! >�?�C��c�l�����W�۵�k����(�j6�;11���E�i����(;W��b$�]�2�b��Iz]�$q�
�y�>�o�	�_�q�N���r؉fC�(����8�{�~0����O�S'�8�6�[6��F��"r�5'�d���3�`\��F�#X}�Ð�" �:ʮ#������)|��������f���,	`��=Es��}V�,�K��2^�u�dڐ��3�U����<��0�8z�L��Aj���u��t��>qX�X7Y�{tk�H�����#_�,�ZMs�f�d��fpç��>X`���Dl���~`���
����H�~q<+�	B%9��d~�I��gZ��h����Ĝ�5L�p��d�|m
�3�9+	��*�P���zjaZڛ����P��8֮q7-�C�б0ܲ1&�g�#�n�W��>-%s#0`-95c_�1?�5���E��J9U�F��3Ϥ����x~qI��J������t]�|x4� �^���DV*�'�m0F/�L�+�=����u�^�z�I�f+A���i)܃_�N_����^ki�o�i�-�a��܋�m*���:�.����4�����mONhWd���^&���Gd|H�e���j���n�:���۾�~�W=������	�R2i$=~�� =V���#�QE�+�A�_q\߹� =�����$�(�U�_�E�������*F�2����<G8��x��i��z��܅A�.���/�������������q��A��Ep�|;��-	�+�7��.}����J2B�{�r�58#�x�V��Vo� �[��U^��?V�aʐ|B�U���~-,4kng�~m��lS���C�Cv�M��d���@��f���B%����)A��/����]κ�&q���ITy��;�fx�ĳ����7�璘���`��d�����l3I�!��!�� +�����0��K����B�rXs?��Wݎ��")�a�Ou��S4cO�~���ۆ.���?�>���=�+�幋.�;݆|��f��jw5���܏���r%��r�'��e��r�67��U���'��}\�����8൸#7�;I��/L��Y��ߪ���a�VK
����3|J�����ӆ���J�����xz"��DK'*�i�J$Y�ư�[2U��:��-���CЇT�����e�l�N�S]��a�����M4z��O�>q������&ʛ�Q��d6w!���2l��V�Cơ������cNV�m�Q�FqL9[��T�[H���E�',��4td��q(o54���K9r��V;%�\G&�<�>��-�u�]�!G�a�<ʣ��-*c���f�L�x�������=����9]�������c�/V�F�dٵҮ!�&f����j�"������ �R�Ҩ��F=��Ը�y �����3�.��@�m�������6�n`j��.����O�~��u�m/�G�ھ���U�w]7�O��i۰�3tE|:]Ap�F��ߌ�������	�K��2W�e���/�Yc;m߁��k����t��׮8������ǿ	�ں�N�����i��6+�'�*ʒ!��^�����:�OL#l�mq�[�M����Z����g������_�g�)V,./mHK���7nf��]3n� ��[q����&۸mG�oâ�ַ�}ʲ�5�✨}~
�-iD���r�ɸ&��_}Zo�u�����q�3���~G��\.��1��h>�Ԛ��8e��m��W�����UN�D�7KX���}��#�x�������
�I�$�gQ�k�z��I格�2��O�:6�o�R���a��c���Oާ55�[OO����>�G�`�m��u�E�V�� k��<|��M�����s�Q1��@j���N���3AF���̰�rs-�$�W��I-v٠e������~V  ��IDAT��mDA�Zg@Ѹg�'������[����۷鑳i;�b�g��F����Y����c@��Y��fA��)��e1"��c?e?_Z� R�y��XƑ��� 2}����8��&���,�LU�4aec����0xP�;$?f���^83��&��,�D�x�cg��t~鄏���<Q��Ȼ�ʎ����Y!����Ss����N����1�L�P �ݐ��u�1h�c��� / (���#p1(���CmCp@�y�|}�����h7���~�#S�
�'ʴv�����[�����/u�Q�J�-?�S�64d��Y>���2g�l�E�4�:6�ЦV�K ��� ��N�1xˤ;�.v���(����M�ԗ����x}�Zk���T��e�M���|�*���O�?��܉�8>4�g�W�^t��0�/v	���hȫJd*<�_�`+��:\Zt����)|?F��\"��I���DU��T߇!y9����TIG��ien�)C���
�Qqʾ��)���y.iq->'<.3)���'���_�����]\��|�n��b���<^r�h�Ti0�f�k���D:Ĥ-ʇ�%tp��$;��ѵ�`��Q�,�G�	Ɗ�N9:!t�Pv�y���Ly:ޞl7�U�F�qxTZ;rZd]�� #��@�#����y ���*��"O�69`b����13J���ORc�����N���;�#�>Jg��U�<� ��'�M�����:]�V��jtѣ����H��g����Ư"%�T�$R�k2���<�I�AGwɥ���vsJ'ۓ�^_��HU�-�s:��K�W���2��(/���4�~$Ϊ���
��w�"�w^��7п�;~}�w|'���dv�C`&v�al e���+��1W��.G��
{���}rm�SP�����?y	�>쥋�G�p�0��	t����ת5��/I�$(�ֻ����Q��H3M�&�֨��!uϐBV/"]̸u2��u����tgƷ�C?Dӥ�Uÿ�F�^�Ooz�黿���K��K=)CI;x=�qXD��-��asFC�I���� ��Sc��VL��]3xG�%��*0��o������Ϳ��雿y��g�q]+����d�<�;���z�0�*3~_^���/���L�Fu��a�pdc���vC�I��f�AZ�\��� 
G� n��&5�I�|p�!Z��u�9�q,[B�H�����,A��&sdMF�]�aؤlǅ��4�k:Q��,�Y��_��b����{r�Ltn���7#F�.�u~�P�uK�b���.[���g�ct�I�G��*T�:�mF�]2<��V�iHj(&�~�ER�m4yY`[�,��x�3]�_��t�eK��fSn�uv�x�>2�N{Ƴ\��LH�*T�}��_j^y�҂+$� Sk�dc�::���C���#��^%�Mˠ�m�&�h��~�H3�&���rP5�ՇԕW�/,�x���O��T}��`���\�մ���~��5��r,V�ܻu� ��^1�Ή�{�S�w���O��LvN���^q `��L_��
�R/v�_����S�΂���[�q�s���f��
?ƪ��� K䎍d�r�=���Ɵ��2h��e�g"���^C��ܻ�>��n�9��H���d��8�^���d�poGv�t���X���F��2��r��{[l��?/f�����l蓟�$}���f����sާ�=N{~)��fC=9R`h�����aJfS5#�^%���|,�˂�p��eJ�ם�c��5K�^�ծO���H���i�E��:�ِ���|�S��Y��|2����~I�=��DE��\�PM&�9�q|�Wާ�鲩����(���3Ng&ϒ�:�sx>w>#�*��AڣڭX(�#�uF=�
��7{�ggB��eŹ���e?f�́nƠ�z3�`��>7C�n�6�Sz&è7Z�/���4R���ںj� ��᝔AZ<� �w%&���3Ȫ\`�$�cVM��&�)̽�.#�-nJqnGj�ϐf(���
�c��6�5���� J�t>6��ډ��/�F���։���
�e�-�ɪ��ݪ/����|�uz	��9���Sr�����14a��=��Kc[��&�Yk+��ϔ��p.�Lo��w���Z�d��̮��V'�UP�-��t�+-A��ˍ�X/qR������0�o��ہ^���@�)�����y��$}�7~#}ɗ|=��C�Ѓ�3g(�����Rx�f�uW�4(E(���abԝ5��N*2�t�� �����n���I�;��؏��8� h�f("?CY��-PmU���R����m&��rzR	�`e�Ȓ�8�|����e��1���Uk�-�Q�u��=�}x>�����
J$����:s�S�Uy�@�`v�gk�bT��H��������L(1ȃ��3E!�gF�@S����N��1#tG+�j!���o?_���:��O�I���)C���U��͉|�LgI�[��C`Kj�d^���N�]�^����Od� ]pA����7�}xu5��w��{��3�w��m�+���l��*Ɍ�-S�!��DT.�e� -��'��C��h�m�k�tn�rp\۝�f�����گ����/��?��8�w_��<(�oR�d�����o�3�Nox��1>�.��3��nO�8vx�����g������1
s�nDG�4E�c��
����>3��h&�:���A6dH@���܈�ьÌ��2����}BD�%�� Rp�BU��<��D���g$�21��g$�b����'A+#�:g�1%=�d�e�S��2����o����S�VoB�.9�@���|���[�����_IEs�����ׇhv�)��i|ߐ�y�dk��pzz*�+���8�G�Q���ٖ�w"��]
�6�D�ˊ��K���:i�]�Py��{^�������@��m�>���HS{F9V0�V��\��s�p! x���%�/��㌢�c�O����%��޴䁹q�A�Z�� Ͻ�aq b���k4�hr`�-��=?�Oθv�~�������:>B�=?�n���gzz�<�Z���^d�?��z�~��l�D��g�#X�7�y@e�Y�of�'YTK��7��?���8��w�ٌ�g,?�=�i�+_�$}ٗ~����E�NB�� �s4���/�������G�Bȗ�f��x>��%��&I̜� 5������xb��O�n�C�9�zH�m�����#�{ׁ�ؕ���3�;*�E'^e��aFj�V���J����gv��L^�LC^����,�7�wq��j�s��cP9�n�#�RB���o��>��j\,z�Q��#�j�hP=D`��ֹ��d�ڰ�",b���a0�v�A���e.�͚t�F��>�ܧ�~���O~��O�����?�n�������e���W��F���J[T^n�=[���S�]6���|�,�f2v� A�#m��(i��c�پտҍ��VO���f�~�x�\��A�:�Y�`O��������3��C|T�8�M�LG�7(N�~J�TR�%��D&:7��M�1O�l
�3e?zwiK��Ͷ�:��:�N_�^�5CP�d9&���Y�s����5��o.qc�Ky��S�#���JP)vE���3g����p�� �GpG��<�)v��ϰ�p65c��	�ު�e�n�Y�4�Y�QNOn�u^����^����z�����N�bH��PcO��ʱ4'
�ǽ�����c��	2N|���16��@I�q���zYҼ�C�z���vlI�iG5�7���|s]0�k���c�w���m�q�;�Y���
{ɋ�/y�^����< �2�����wʳ������<C~����O~J�����f5	�B���	̻�k:i}N᾽A�V���6�����W��J���?��Rq�����a^��H�lГ�3�eة�:¦S�.����M@�a��̫�&��m&l�g��g ](h1�>����]3�a��0�i�u�8Q�;!d��92Ұj^�;� l�������(-0�ټXٱ��&��`� ٿD��wc<�n�@�)�E�YɂF�n�M�F��Ҷ��2�n��h��dpA��8<�:O���K)�Y�+>�ӳz�������^����+�>�,=���CO=E�<�qήV`��A[6kmD��ڐ:�����l�x���^��=�ٵ�kzIkO�Kn ���L��M������^���!u6J@҂M�ZL�A ��!풀������?�ʀfx�~y �+��Q0o�����Γ��C�,�
d衇����o����7�ؿ�������#v��)e�*:�Fz�)|n�IzV��ߙJd�D
��g�n]�5�
Q��I����cH���	F�8w��52#!��0#
�����`E�.Ug�r��:�9K�0�[��Zu�q�{�fOv{!RН�U�O�1�?k\!�8��	�)l�P?tpǢ,#�5�m!��R��2�{P�h�G���i0�Gv4�0�k��qWƴS�xd�a��r�1�1������3,N~sv��H�b 8����������aG��A_��iٝ\��&<�:m�Swp�*��!���(Ԛ��ӝ9%��A>��f8�p��V�f�t�|���x�o��y��O��?I���nw��ZШq��p�d�{�}�-�k7a��	�ȁ.���.>֎m�W�ᘢӱլq\��h�?�'����a^��eC�׉��m�y.������q��w	+V����h?�(�Ҏv|j:]���ϛi��dn(
�i��_/G��Po��+��o��9�vl����r���R�������SeZ��y�V�ܙ#�����8�Q� "�'�dЋjR�c��:	|�h�ʉ)2�=N���R��J�up�ݿ�=�xl��%��r��A�rf�0�U�?�uzf�`FW 5�����Gy���_E�\q�q�49� �t�ת�l���D�\�z1��`A	�!�3�Qd�/�s|�nor���'m2ȳ��;Rf��5��?���}�_��$�,u G���<n�T�f)���:tD�\�D_��>g�����w�N��[=�=��&Bv�o��j��a���.��gZd));�qȂ�����v�t����/��o�����~\e�Q��)"����L�<�0}���|S7Cv^@$�����p��b8��#��8�J�O[�U\� h�G�*�?�n�j�?0��OAv/��X�Ln�uv6�՗�?����y@�����B����/~�ӓO>�κ2R��D�YՄqS�e�2�u�>�����~��=�471AO����9"�����T��ыB�_�=��� ��_��`72F�4G���>�8ɹ6>O�7HdN�aL�o�nj�˓��Y��C��q��M�(>���E�.J�)��'�V���ŬdͤʽS���ku���ju8`!� ���I�-@D����3��C�W$X~�\..���7}���7�Ư�?�g��~�'�2��@[�c�����󕖖�ci��Lǩ�
58h����|��V��`jֽ�^�F�墖�UsȺ4q���	xΚЏ���Ro�9����f����Q�N��������k���Qs��V(LW6#=���$9�,��^�<��2��֮&:���b:'��W�h
\�:���z�����9�F����Yب`���a�XG"۳��d`�x��Q��}֤�G�l8N�'��YP7��->�уW�F�Sj]�u��H�E&BP9ڒc;�E:vJ�I�<��pFJղ)�?��[��A��
^�G�Q�A���8�ۑ�IZ2���������?�G���B=��tZ�J���X����k�����4�V��
�/�T�������C�c��Y�+T��#�(c�C=����(��*կ5�$�en����...��}��o���o�Zz��/��|���wHF�"GB7�?��;��|�iz��O��,҉��)YAن����u�Ͳ2wzVL��'��hH��ftn���$2�duAV3�B���	u�ߒ]�T�)�f�Ae;����]Gd��4���FÑ�n����'�3���� �.��3JKyT�_"�VE�J�u\k���-=)
���������f��XC�MXk�"��X�:	g���1��Rh9��{�=���q z�?�	:I��e�*�t�v���bf�_�����gdq̞�"�[C�!�4�>谀נvڵ���'i����Ӫ��	|�~��-	���{��s^�Rz���� K����]��������0��m�G���wѝ;�ض2lΔ��74���X���$�W�|�X\��QzW^d7O�k�K]/����<�}sd����zPà�g��0��iޜu�6z��7�����B <x�4.���c�IÐ�%�?��L�b���koPbJAd[q�\LW��z�W���/K*Ы��]�s�3����O#�`��W�9�!�S�z
��|��,�«Sm��L*��W��l�4m���@���90�Bäm�P�`,|�$gt���VGygL���	;�'=
#�� �!Ȝ�	��*���ZX�+�^"8�YU9��éDY��լ�gع�)�4��^w��c��hn���'��}�6�r	kk��ЮG�.�p3��1.�s�;�#U��#u�<0�3H}�1)4ePE7+�eM��L�bC���Fq�3��`Hi
#3��V��y���3�u�р������ѹ��#�ʵI�U�M��Ng�1Q#f�ɮ��E-o���qa39[�g��5�y}��9����K'�'� H߉g�Z�uuo!0�`�0H���C5���Scp���J�9Bh����������;�vu]��~����\SZJ�X{/)mN��a�Hp`8��\�U{�xׯ����r�,s�#���?�]����k��_�*z���H_���Z���Y�y���|�����y��ߧa<IǗM�Ʈ4���Fd;x�V��U�ʍx�K("���7q{V�sm{�ǒz�����ð�x����4~� @��\j���H���Cd^���ؕ9i�7�NL�fe3+�ݙ�؋^D���W����,ӌ4��vli<&	�4r��Gy�4�Uy��c�O��Q��1�crb�wɍ�crw�g9SZ�y-]���L��Ł ��⁌W&��F�����m)_��7��<�r�ЇI��b\i��je1B��Y����2o��B Ie�5�^gy�w���T��Z�u�=���(u)�@i[�</^���t��	�cy<R�(jx?Q��$`x��.�y���x�%�{��rFY�ˋ��p������6�"��Ԣ'=�G>7I�1�Y��'�K5�ȋz�����Wh:��r���(�%u����T�I�mA�&��oُ%)b��^��n���xǰ�����j��i���u���	46c��j��,ޤ� LF`9�8o����7RE�9@'P���ꊊ0xЦ�{�z�c��3X��xG�_�	���V6�����4�x9�i��^�H�Ʉ���d�9�v.�z	Y {F���k:�pĄMQV|�{�=�I#ۼ��T�w����*���Gy&�x���e.P�n�Y���Gږ�i����D�d�V�c3���_�����_�R���~�ď�8])?�1�~i��uC���)7Yz�r�X��F��~�O��p�ڔhg�D|�e��i	����2����eM���9�S���ծ�(c;I�O88�%�cu-���Q[�� Z�^����+m���I�������<��w�(������E��勞���Л��z��c;���?�Y}�9_d�rl�G?�4��>��:;;S�� �W��l2"7V4������k��g�^�Z�ll������iٞ���������R�
c��[	_:c7�
x@�o�����9����~$4%B6����|��^E/�˅w%��>�Ѓ,��ޟ�z�O�<��Ͼ������=��YV����ҥB�T����B��F�b�5Q�z�r�&��I�E/�l���s��h��S�OJ|�ȹ�����ި�џ͒�o��/�pc_:t%�zNM#`��Ά�19LL;K������~ۿ��������Y�~�����Oi��DNbǀ�W�N}���� �I�-=fs�3��Y��o��[]�/����dy��8���`��b)�m�~Ȃ�=`J��S2����H+��,q��7�5�l��)�����p+�mƜ���G�B�P��LU�F~\���#\��%��$�����1�S E����W|^wLN:�7�>2�~�! �ei�A���`�E
T�؞f���6�(Hvt��<B�a��|R�b�� őa��p�
q;��D�6��(l��`c
G�X�b6�`�V�3�y�`����tp�+]�O�=��_j_4�v�a��f8���1�w���Ao�-��~�~���o��w����,���zs]�'|����Xב4W^�>���,���õJ�� 1n�?�&�<r�l��ǸFU�8�\7�CP�%W��/��ׄڒ��A��t�+��8EJ�v�0��P��; qn0"��r�>�
�}�)��� <Wц	{��gP������..�X����b �A�&��yn�=���C��x�)�Y����+a h�9��
_Q����<�().�`}`��N������g�S�c��TZ�E��8I�[����;ꜳ�ˮ6C���}7��
f��z�s��	݉8�p~�)��\���A�S����A�`5�F���6�m%d��!�8��x�X�K6�uV8���('
B\��i9��n�F�.>�wW@!�y6� 5���u\�I���Oݕ7�P+gA��pz{�����dV�>�=�y�4���ǵtha��@�"s�q�:4���%%Onܰ��n��֛��H�m�2R�|��L��4
�q]�/S����Z>An�\���Gw��
گ�L��<?����f�i{rF��羋���Av�]����U �T�N/�6a�C�5Bߣ�w>�Hft6� O�F.|��T�53��囔���Z�P-B��RY��7������wfU��(7o��j�N�I���;Ƕ�δ�2oݾ�A%���[��l����)m�O��H�^���4��EF�a�sO�V[����U5%�b�dXE!f~�����@�l�0��UɅ6NL�^6��|���=��ȹe���N55�p��Ku�,�������#|i@he�@�&}ڱ ���fe��[sF����}�G7���r�:�r�������t���dl�
����+�|������v%Pv7�l!�{�m����[�Q�z��W�Um��!V�tñ��F���i�D(�b����e�(����)�v�1/�nl�L'J�lB��r�8}�qm�Q��v�]Ӣ�"���3��|צD�nia[ޏcg�N�p�2N�>�f�p��@A��Տp��mi�#�Z�*f��r�^땝a�7�mm�i����3��~��hGL~���zZ��h��9
��Е�-*���𜐱*�Zb�T��Ӗ:c�)������Z�+՜k��:���D�H���HǄ��|긥[g�x�K�-ݾs{���a�y�Qx߆#��l�}zJT�D�Qޏ��1�3z�����dk��Ƴ�%c���f��>�������r��U���(B���!��𰖸�6ϵ�yqu%ժ6p��d��>����W>��������s�x�[�u��J:=;��{��}��{�v��bƱ�gwx��xhƀ~�s�!"�2!��Ǟ�M��|~��>3���.�90�t�}��-�0ɲh��a���g�� ^��Yת�<��{��5e��f8���g��l'���G�����[�K���=��gi�����WX2V�|3��d]�6x#�,��A2H ݹ\���1�3�2�P��-ja-"�������Y��V��92y��5=�&N��U�G�����uY�]�a�?n�p�hv�oz���������=B�=�)�vQ����uY���O"���me�/Ș�%�V�bӛ.l��8�����kc�7�4�M��Z�=A�x�F�%��8���{<�X����`����_~c�k�]V��\]��
��﫷\��>�ߟ�O��PY)d��ޏ�)ss-�_��|nb�F�ll��2d��X��XA��B�5�F�1�����;
bv����5,��6d�m��܆I5?��N��%�Jp����ތ��D7�Lz?S}66�����FȲ��a8a{c��b�,�4<�����3���I3���q��|lP���g���}v���-�����	��0������(�})�Z���S����\�+���Q@fbk��}^ ���h46��G(%���[M�J�_k�۾bGX�y����w� �N���.Յ���~l���w�nݺCSI�TA9W�dC�J|ʹ���F��O��oC��5Wu��w���L�ҙ�v<�k��&<���KR%��$���S!z�Nwd�AH���|0q^���O0k���2Y�=���z����\���_��P��K|�^{�wX<�[�M��f��-�D��}���w����);����D������D!.W5kZ:��V���7X3mqH��hhܦ�$`��t�6I��3B��b����M��ʀt�UB��ې��g9ze��N
0�a+�78u�(g�=��SͼcAmd�5�}���Tϛ;��
S��ϱ���1e��#8.z���>�	%��}�^-�����4U�x$�F9P[�Ꮍ�u|�#��������f_�`�f���v^:;6ҭ�J�p|vzJ��Ϳ������y'[1p�RIeϙt�*}����C��9I, ��TS�r�M������p���>�'���ۻq��L�e�!�u@�x�!j�CQ��t�T�.��م��V�����>��]vK��c���^���ٰ���J�8�r��P˹ϟ��'�o�!��o�f2�������S�p���N�L�$�6\�M���P4So����v��wg9���lĨq��VH�a�b,V��g����7�&}���͙e,#��P[���J�˖�mk)4%j�]�q�C@Yn���ӎ��Aa�[��e7/}�����tkj�1lox֚.��}fO�o>��4��=ѐT�{w�I�������җ����ȇ}�T�u,��'>�1z���~�������}���04���ĝ�f�i��na�KZs�械�!%s�^���|�\�Q�z��B���������V:2敿I�m�^��K��)�)-�MÄ����T�&=o������%���M��=�?i�#�FkeIOq�V�qxv�$�]��L�xt1�MC���^Y��df�A��2�j���Y�@��a]�hA3�&C�e��8>h]����a'q0\Yݐ�������O���a�� 3��R2��˪d��#��F6�kP9�v��֨לC��Lv�2/��G娮R�6j�MR�g��M����ql���G�8Ƞ.�.�JK��{X��z��bm�_<J�D���`ҥ�(�q1���( �׾�K��g����Tk�S��M �1�����c�����z�s�����/���k���J�@h	x���C>�G?��zKdM��<f2=]�>B�<kS�k���a���d�$�d�B/�JHO�vO�L+A�/�]���/��
_)��ɭ:=�E��M�J���Ͽ����&�����mˎ�<L�,g
��֦cf;\�x��;w���O����D��|�i�o��p�L������g����uZ��Z��e��P�nU�=>�����s-hT��J��v�?]F�}ɪ&�Qrt������$��{�wY_g�6���N��*E;�چ�"/�>F�b�P?��_�}VQV����`�l&T�,ȟ>݉�#��d&��΍�w�5��{���w��v�ī+��ض�l#8��#X�e�c]&v�{�׍n,Jr:i϶,��_¤_S"E_��yik�\K�g�l��̿%��(��Qjj�,�L\��OL��m�P�4�p)WD=��g�
6���&LZ;ݙo�C��n���5�������k�CVs����y:�r���.��h6������A�����.����3:9�l��lNg��j�ے	�6=�9O҇��Q�t&G��LE؊s����ܭg?[{n�׫�3�{���%G�x Ң�Ĥ�,��)�;j�H��r� ��C�!���u-��ZA�oal����@[_�޽X��;�T��8m��#���i����R8���g��^�������z�}r���*�I
rZ捰;MB�� S)[�і��hg�(���Ԓ�n��ܙ �/�q<�K�1�y�)�#J[�q\�M�E��OA��������8S��p4��)!��p.���h�1C�Pp�މ�ע2zS�w��WJ�Qz]��K�G Ř	w���3�hV�a��p*N�!Blq�X�N=����we�����,z9"\��ƞ �H� X`v0~2��� ,'m�}L�D�0VX�n����K9W�V��|��+e~N����G�:�� J��crL�������Q1�N2���u��@�����r]�>H�����q�@K����[��eL��'�t�ӂ�k��L7iq�Wy]C����|�г�k�M9�5�|[_m�'���\w:$z�W����������}�Y~J-��Q�k�-�F)� ˔��ǃ���G��>��1�cj���s����*���ƃ��Z�C��N2��.c�E�Ҏ=Er�*���n<��\�	�;���K�'[:����~H#��U���gI�]�{ �����@w����;g��q��:���_>����]9~���)��yP�*����:�������;Rc���9oxg���;��������t:˧؁��q�X�D�fq<H ���TIq9�.������gߙ�|f9�������%=���:RP�`.�����K��vO��^�P��k��yy���{~������*�K>��s��T�*���#I&���W�
=��������O�x#BZ�H[�Q����������T�c�T@tp��>�K�L���w�Ŷ2���yM�kD���.��M9�f�@�,;�7�D��ςj�*���5��b8�� �B�*��[��F������;)��U#%蝮����KT诤7Ç$Mm��H�g�dz�t�f���	�nh���I�8�-��йs�n��$�����Yw&�Us@��tjm�?:�<����3����]���d1�r[
dS�Nz��಴�&I��L1�͟�'�^�a�����=�ԇ�%���0���9D[��
�7�7��z�9?��q�v�(G=ۃ����::�MJ������kh�>WZ�շj�hh�g�����!\o�����ᪧ+���ϐc�T������F��&=�DR�߾}��櫿����������t�Yw1�����c�6�>o�ӣ�F��+r�h}sY l|�8H�sί:�̾2e��Vɭ�S>��9)�Sz%���%���
-wǀG�29 +%�}�Q��L�� !����%�z���o������nz�O�$'�#�w
m�E'A���_:5���{���O�6��;�:��f�x��$�9TTE�@Q���[&�_�+��zr+'�HG��b�R�,(ՁIKNm��k+�O��p$�݃�jP�����պ��D�
X����cbڹ���w��x��@w�ẝؘ�K��_۔��R���m���
}�����7��r*kZ4��w�ȧk��ϒ���g������ʹ��*"t:S�eE�K b�R>:�+�y���"t�}=K�n���1dYy�>�2�B!oJ}�۲#;&lp�4�#(�o��k����QN�r@��Jc��&����U}"�]V�A.{�;�<S�'+��4����O�/ǥ8vj솸���F��U��v��uE1_,hf���j,�˃g�ذ���A����e%񉊽�ȒM���O��<���H����]\ҳ�ݥg���v�S������Kd�^�}�����k���r�m�@�K�m�>��b
���gN��V �릲G��Q��r(B%5�[n�h)t�yG�#�������/��1 K��pC�$��O�����w��������#/�[g[�u*i�K*�b�`c=GJ�l��`Ɛ�82F5�T��k8�
B�����H�q�i���01���)f��;��QY)�ϛ���N���Y�g\+�yf�M)נ)U��C�mG�����-��[v�j=���D�?�9V�>����F~qL�5�aN\�5'����s��\��1�i"3T�x��	�~A����|��S�9��@<Ŗ0��rTC%��%2����Q���<�Q�v�	X������%.v����\��R��D������9�5ۥHr�x������#�2�ǖ�\���4�|�%�%��#�$�x3�p����������$Jp�Q��e��N
 g'�xE?���������;���`�)��f*����ct�ƏP��[�R,ڋ�#pSքG���7)*��0�s��Zp׻Sx�����$��O�<��*�,�+�ђ����?J������,�B
]*FRd	���J�/G-�g�WR�F��VF$�;,wr�H�IZOo���^8߸��vc�����:�ISY4*�oW��,"��SUQ65��U����xG��G�8���=�ż�#�w���/�[�F��L��fҸѵI�^x{�w3~�������������^��W�O<A<� ��>)ΥA�Za�-E��T���! _��d�w~�b�kKox��5�;�L&J��~��O����������������N4�%�IA�-��qqqN��я�؏�����T��-�����VQ�^��l�F��O�(	4I��YAᰇ`l[�-=��[�)��~_���ݫw���^OGY3n�3ޯ�M)�s4��z��ӌ��}2�� 7uZ��>E���uz�/��#O��O?M�|�i&t"Ǎ�/��v��������
������M��׼��n��@�+���I*�ÐS�����_d����	�`�[�c��I���2'>��2~�a��ȷ���3�_�y�����c��<�S�YIeE�(-ZQ��������ݻ璺vw����il�4h��h��뛍�'�Qy����	sY
v�T�a�@�@�E~�9h��QV/Ի_8�l	����KIicmܬ��'���u����j��\��.��.r��o�qD��q��>ʧ����w+�]<25�Uv\�T��� �X>1]re@a�E���i��5R�b���L��0���Ca��m�g�is"w"k����{J�+���~1^^�9�5�g��<�yz׻�E?��wӭ[g�Z�0�;�|mV\����g�N�B�m���3��?W��hM��Vye��C\����n�ꕞ�[ޒ��'����r.���~�����Œ8�͙�з�������z�ч���;�Q�l�%�u�^�m��,e��<��!y״>�����B���
&�W�k]�\�ϖ��0��@
^��s���^�&Ǐx�Bb��cԡ��s��U�e�[�Aj[�vV�4��d�x�;�g��[����������5��:�o�f�,Gn߸)����^ƙ*���e�E�lӑEH�!}��'��*4S�8
9cQg��նS��^�O���O��z/��t}��21���&$t��g�������o��_O��|�A9�*�Q�g�n��Xb>
]����L{l�f��Ҏn|E�=nۏ��.H�*[�E�\2�Ӑ��b��̚�{e�pO��ex�
�#�����/�S��)Ș�>�l����8T���$��A�C	�͆���;)��p/��I�eA?\�v�wRY2�O~*���?�AW�v��|b�'��"�C|�����������,�m�ID_u�T鯬� T�0߻��2 ִ�A���M$�ӋQ)����ɭ�ր�����
<r%�Ps��.�.����E�<�8�'M��QP6=:qM/�f�үb��d9
���>����;W�Q�n3ӎ+�����ߧ��/�����M��6e	��1��.��N�-=���g[>U���h���v0��љ��3��\;b\Jo���;�����8�r� �'��-y��E9I"wN��M���4���1U�{"��Ȋ��lF��#�K�%:M[f��83�	g�ʎ��	t7	����w��r��EM��1���Սf4�c�#ȁ�e��6�;Q`�bC[f�� 	�<2R"˴=ԓ�ͯ3h��:��+;q7z�]9K��Z>{[���l�y6�Bt��!�uF��"����iOɢ�� ����T�v+��l���R�z�֌�Fj������GEk�j��<��0�A��v&j1�%a��f�`�B�ʤ=�.��q�h�Ƴ�uL(��SJ�j�B�pD'a���Fx��0�}�|_).�=���h��� %�d>��tI{�*�e8�eq�m$��f�^���	!~NZ������>:�t���.���zP9��(�J���rh,�����Q�%\4���%���N�-�E����5��~��g��_���;�^�͓�+U��+zd���ia��^���z��M�V��gn�'Zwk�N[���^�=��}-�x#�<x'|;!V�B�=�;�ϋ���м�jިD'�A5�!�G��#������#{����؍�ƢlA��E`"v��ͤ�p���^��7����}���KpQ9�k���?}��黾�;y��s�sn���s���d��"t8���.�h@�Yx2yqyqN/~ѣt��tzz�JQ"���)6�qWB��kN��h�8�Ȇd�����v���B��}��f�����l���$=�ӯz�L���Af�r8�Ϳ�o���ۣ�W���&���%��O�8���1�,��'���<�~K�[ߊ!*��Cj�*����|�)�G����������
~�׋1q�ݹwRe�1�H�h9Fq»A&:�c�to��zzp��><`�
��J*ڹ��~x�OXF�:����3�*g�[����-$+Ϗpxuu��WWW�3�%>�^�J_'�K ����(2y7'5��l�9�`���ydN�F�#U�eӍ܀�_j�`�뢿m��ou����!���J�1a�7WB��� �� ;>�� J��9B��Au�B��B{t|��1��.`�)��j��c)��ؔ,�h*c14D
�$3F#�!g���hp.<a3��]�ؗ�#oe�����V�^�ԲՂ�]��#�6�at+�2ޤBY�۪�2�5k�w��Un�3ke�_7-M����t�e���~�|�&E�=w�6}R�2�a��ڻ�|h�hW��Ě�q����Ï�o~�[�E�,{uyO�^d�q��I�K|k���}j`>�~$؍<@k �\�����}����{J۷�M��R�CP���̝��o�Y�*�lM��pdjt���ln�q���y2�+��<���m��O���蓟��d����춶�}x���~$�,�O{j�o���Y��{-�m듊Tits[��I���U�כ\��d�5�폩՛b��t��ݪ� H�w	\� Æy�6a�A��:�Qt��y�����D��I�u���f���,�ly#b�dQ�O�vv���v��g>5�/��l�o����z5/!�G/�� ���vL���v�3��}�
"��F��R�M6�u� qC�c�W��͈��G�(�$	nٍLq2��\<��lӮl��?'y�l�� ���3٘rrr�>�Ѳ�s�$&g����#6������ȶ�I7�l�3R�>�=��|�6v�`xm��g��cfˎ��:�v�[f��H9�E�E��"Q��$��8���F� 1�8� AG6L� �#HĒ�XB$H�d;�m�6q�)j	II��eHΐ���{����{N_U�۷���͛!!�%�|ݷ�=�,u�~U�N�;Wg{>���]#�>Ug�)0Hw���`�aV�g���x��K�!N�Ao�~,8��1�ة`�k)ܮ�����9G���Ck�X\Ğ��+�ӭI�*�>��r���*����lEk?�e����:ߣ�m������SS�J���F�G:�>������F��"��Jv����u���{��q:b�;�;�r}u��l�{?���_�*=��3������_�~�7����|�.��>ld]|v�=�}���&u�+���i=�u�����>�E�h`���6mn#Ɔ��o�_�b�$6�u]4�Jm�8�9Ma���UV�B�l]�x�6�i��U���6#d��9C빀s��{�q�~����w����U�xrvBy$�j,x��_I���Wӷ=|�0�ƢA��g+f�����ɸ���ucj|�ƍ�t��9���%��A�B�4p���`�0�$J.8��76Ǳ�,�(����N�T��u�FPl.� `�L98~���PLj�%�Z��p�yWA/�"��u��K��u���8�؄=ݴ�)�P�N�I�Ojw"\�;L��0�z*bP!	#!�� ^�Ly�G������y�]��;�@� �����Q¼��p���z��� F��䍭NBB!�9N����)����H(�"���E�����,�nS��������Xy�5�8�G�G,D1k�W�a�<�D������7���C���nW5�w�� ��L��ww �������O������_���|j��?	�Q�����}�j����EooU*S�Zo��m��26 ��׵m���`9�f6��dy� ����=�JY�=� �Wy��<f� gc(���4�����P��wldm��M�oqB٫}3��_t�����YVaC
;�k���LY���\�d9we�׮]�o|��.�K;l�^Cz"�mU*�k�K�$x�ٰ����Ŧ��רI]Z������q|t��n�1-�_k���ﻗq���:,Ǽ��/�X9�DL#�d�wE�:�R1���W�T��O׬�����8t,pIV���7�i5$���`�)>�U�8��:6���e����t�i��^�vٳ�V6뱍��ƣ���	/��@Ƿk���:�ѣ�<B��?@������폊���Um��,~:�n`/4R���/���]I������zr�	'�N�Z�U7:�o��]� ���"<��%��s\(����NYu��'�CD���M�������1c��ｇNON���+t���˜��TC��.*�j��^#:�>U��%��k�&�:�ئ�q��:Q����6�"��0$����2����r��
Ӏ8��������O�}��dB�x��f�P��vࡨ6A5S��m$���9R��uc`�SN;p
>�V
;!񘇓i�I=�B�����T��;3��]��8"=t9`�):vf�O��Xt�|�z�FĎ�#���B�:t>���:M�/�Xώ\W*�2��s�i���V�ؙ��C�����'����K����ǵ����߰hcj!�����vkj��Û�߼u;�9��v�4�ȵ �{� �(n�C��_(�m�]�}z�6ǧi�� 
~ԇ�?S�wũO�O��������ҥKt�=��͛'#�X[�5;n8�r�����I��c
�C�9���\�jz�y4����>�wW�]��q�wMi�����Lߝ���;�`R�W�1k���|ͫ����?J��O��t���0Jo�v����mc��,3����aϰ1=B2=���R���̌{2z�^>�A�N�lyf��3gڶ��m�qŅ�_�dy��*�Z����>�����J�|�;�G�O�ۿ���#D�zv2�OW��G��}�7���^:>�@�Bk��e�w�d��hk��W��T<.Q���X놹�\߀r�x��A~C� ��ٻ �1�o`�6�K��p�0 ��$a��l����H��X-��B#`#]J��-�veu�],%��ѡDq#�z�M��Bm1�:yȿ�;�TЈ�}���n�J��b�~��`_�S\�>l�2F��:�G^����n����k�ÇJc���:#�9aH$Ťee������
G��j�1�y[p6!ӕ�D�@Duv������"�����~U��V�tн�J��@�zP:VZE�֕� �P;�V؟2s���!z /���C�Inë�{B8�0��Dr���v9��~M��.�w	���;�����ܖ��#���ۥ����|/��m�M�Gt8�y����SOsZ�_��_������N�2�^f/z���f����/�����6;��S������k��ƺu�Kz�c�s7� %rpt����8��rV�0l��6��t�����_����Gbn6�C��P��F訢���P��:��ic��AtPO_�09����7����?�������=w�I˺ᮂ�^�a�Q<�-6�ONN���;r�4ϔaV�h�:��!'�څ��2!�m��bKؼRA.9b�2]����=8�l�� K���`J(�hp0�r�ӧ��Q4�4�8��K��a|�E��#=�ɦz?�Ѐ���F�5,��q��w\b�l�}5�fkh��D'1ڲ�#7���ܑ�%���9;�<7}?��ڽ�=�"<�i69d}u��B��2^�����8W�"݊�.B]�$N	�e��oW֐d�N�,D�b ͅ�Dyލ{��t,� ]s/�im5`v �p������?L����󳋑^��IR�ztX8�`[�i�0�OQ�v�/���_~���?���E��HW��f5�r�J�[�����V`�k"�O��V�LKn�`{{}�~���a.�}����������n��u~�J(�W(v�x����* �w���k�=�>�ȓz:����ҥc����j��(:�T��۟�7Fy5���[�h���|��]�Bt.��-�\�QB[Rj0�GW)濞��iT>��/T����M��U�LaSWڕ,ݗ�R)��l�Juh��Ku2�F�VF�ҳ2^��8�����1�}||�7�NO��47f�'L*O䐣�⎠�����B96��*E񯏽ˬ�8~�'�7D���(����6^�M��6�����=�2SzZ�O@��"X�19lce<��׿qZ���/��#O�X�:�s�]���^�ȣ���F����������Gd��離F���\��i��H�7�zn�1�*�L�zH��0�Q�b�{���~GT6��8=�NX��U2C�b�F(B�����N��+�����3�F����s��P�ɤ�y���+^A?�c���u���I�P5�q����σt��b��@�]Rh8b�9�o���h��ˠSD�Zk���F"��yp��<]�|�o���j���ͼ�6D@�/�U�.(�̓��ZS�A"G��m�#�T�tMI��^��A��b6��Sim�йЇ\����LDqЕ���F�"���eO��ӝ��a:�������;ݨ�B�)y��t�;U'G�9yO���a��9Y�m��v�s� |�;��%�vR��s�ޠ�����_{���>�I�z�F��8Z2fY��Ri�����mF�5l�S�D�66��R�of�'���V9�R��D�+󣲳+���J�Z�����z�g��"ϔB?��*����!�	��d�f���7�<<�Q�R�Ӡ�W�&¶F�$�������P����z�����R����Ǿt�9sz���]�JL-�4`�w[$*���I���:�p��<�a��8x��CkK�'?�o��ݟ�Y�X(���Fn�l|����7g㙾[��s���"�������'!8E�LH:o�f:>����l �ۢ��:�"��ܛ؈i��5-�>L��G����8st�kp���M���:_�~�b��2��,��ǾD�~�>��[��F94ⶓ�����p��7oޤ/����3$��Ep�Gn�~ہ�E�c�?�a�1p�׾���'+�:Oի8Bs���z��Ht�������l��Ƭ��u+����%�}��`���1y^m
���˘�:�A��+Ҭ��@�g�	���"�Lŝ��^#L�.ώ���n������<��EQ[�4�8�v0�����V�Xu���f>p��#�H�q�rpd��G�H�dt^�!ݢ�V�Ɓ\��u�&'�jb4��'�v��Iy�vDk�ۼ���>YIuw�k�?����K��v����@	�U��ޖ�bN��7�$��9^����U	nP?����_���{ﻗ����	�O?�4;��i8]�W�|�uQ�^>��Ke�݊܍�6��o>��Oy�y��xΚ������}�5{�R&ֵK����2�~]ԁ�xI��%.������q���5��o��=��u��׮<3'�>k���4/��&0Km��ђ~�O�0��?�������k�'�q=�;�'�va#�Qf�ЕKW�C1o�Ő�y �5%D��4�Q<��pZ��=|`}��~�fV&���@ 25a��t��l*�����(�1o(����(d�"0Vu������8z,����FM��^O��lѱ�d���&,((J�����,�[c&@�$Lhj�	���䞬��vi�����s`���PTd�z-,]�}�J�Ү�+��\�����bG�D�[ZO'�qt`c~�`��j8e��$.�)��� F���q�C�!T���iOe|��rP�@�a>�����-���� �5�$�;�B�V�}�ޝu�5�]Z(0�}��O������׿N��ߣ��)u7�1��j����[yI�C�Y_ϳ�k�5��tҦ(q��y�<ל5"�߇���kcSw���0d�"�u������E���] f��m��9L�M�3��X�Sq�������T���'���r4ʂ���*�q�� *ͧ�y5}\Ӑu���~��A����﮲߄�]o�F���_o����ל���b&����"q�X.�U�z���}����l�x��H�X+��@�0�6h�6��bÛg0.����5z�>2*����>�:jX��������fy��8���6$�Ɩ��T�T51Z��7�u���|3��N�B�BP�kZ9��X�3�����Tًs4Ǜ�¹�n��F{�>��͸���ߤ�����g���n�����B͚�@1�l�,�7����;��;��.��G���~;-�u�}�{�����ƛ���x���qd6#��\Qꑮ�C�tc�0�������)��l�z�����Qv�C��[0LRLfS%'����&�b���^�!֣8�;/Y�����=���!�q㆜&ʃ��R��nP�N�Y_��:�-�KzݬWÕtvb�E�Ѵ�M��d���A�EC4�&��F��A\��D���?��ߎZ���}��0�M1
e��b�U��CM5�N�t����f$T��z
��_�8���t8��"�6�>����ЏvKt�э	��UOS*�&r�e9�ɇ�FL��tS�wL�
 N#�!:KcԮg�{i7;�W������Q�A����Jb�DW��Io{�;�}������?M������+�SI�RX/�>��ߠ�2i��h#�<���<�Y������iJ~?�7/�n�co3�z����fʁw4��Y��bh���[��b�Vg��6�0o�������H�K����1�E�s�VI��GZ���6�mr^�u��-�s질�V�1;��<3C3��Mݝo�����b^ez�ek����:8��d�J��Fw�^�0�z���-Vv�'�8kd���|Wyu��Ѓ>H_~싚��ib�.���6�ىӡ����<���[z�b�G�FG�(ob� �%����� 0}��	?oeU�qn�3v7m�
��]��3��Y���r�Rr=���mH��*������L���>@��w�}��|P4U6�C��K�~^T��v-ӷ=�m�o���+���Г��7��()�!���N�}-���q��N�MH�pQ�	����7�+�3_ˠl�q�0'�M��mؿa]k���zw^`G0��TL���^�}�����WEuf|X%j�h��Aĺ�b���V�K����Ѩ8$�;��E���J��M�Q=}fr�F>�7�v��8�;ew���30!�l��to���W�4~WХ������k���49!� �	C�Y�BW�T>4�Ӡ����7��-���b���?����mA5�l�F���[=�oX��.����-lu_��ھ���T~�n�(+���r{v�U��>R�#ƺF��tzr���J��H3�{��^N=�2��+�?��7ON�_�l�k�x#N}[�#o�6d���aZ)��ó��?W����olz "��!3$E�6o�l��&�{>6�z]؁#�����F�i�c�-�����X�I�I���5��rH�]�=�+ef�mz
��1.�K��
��0:F������'=@����ЙY�W�eͣ��7����_�oiypL��3*�����7�!��l�Kt��JN|��丬}?><�TՑ^(�W=@;�s�����[җ����F��(a�e�����������$��7�8p� ��[��5�o��Q�2z����h�?[lF^nX'��ڦ��f�3�|����Ÿ'��h��AŲy��3�����#eM�:�|��K���4OI,���a�4h���Gf��!HH#�h�vʀ�����[����c���R�Ų�5W�d�6�UI
����bpp�[>UB�8xبT�+�a��}Ii�F��1��(����6�G�ڎϻ�tp��Pi7;U��1����t-��;a�_�c+�t�X�N�����������~��A��ƻ(�,��Ͻ�A� �DذI����tŅ�*3 "�a����0Z/I�K�\Id�����:^��T�����A�gaIw]&k�?Hdrv���h�sT|,������Z���}θ�� 3o�����Dy3���cY1�W�[C�-8�|�C5�%�*�CZ��fv��W�t�S
���S��Xy�	{ϫuޙ�?\�4�B\����$*�P�$��(�W]����:���D�t�F}���<�4����-wF`��L_dW۱F=��� A��i>Z�=��)6Fb�\7��Y����9P�����F���H*��oIY8�!Bʒ弞KM�2a�X�tT8���#^�͍��\M�q���y����(�u}_�j��DW��(�<�[�'�	�'��!�!t?����3c�"��*:�E�_������ ��dӨF8z�{~������-G;▼��ￗ��z��'h��+zqZ���R	.�z�'�Xt�G����u:���ۙ���+b:�mt�9}����9�&;�Hl�{���3�nU��U㪽�u�����嚣mTcO��:qq��p��:2��j��=�.$�K��m['[���W��2��K�Ϥ�L�@7)dy��iDW��)���e��r�g�dV�?�߂�_�u���tR��@�?�t!G�U�=�#��I������R�=x�8�����7����CD�)M�y*4O���Kjhڞit�����8��}
s�kb����WI��/�� Qy��O�����Xn�߅6���GrǛ�L�z��@�o������ag����}��t_�9��H��,�>c4T��F�<-�se]���k<�n�K�E�f��s8I�����V�{/f���z��pZ����<r�;JkJc��)�9� ��+G
��³�C5{��^m���`�9=G?o���J	�;5�nr^y���ŶĐ�ma�#�$��T%��$=Q�n��FR�,ͽm:�T�m������7cxA���|=/ޥXʹ�.iw�۱���1�{I�`K1�4f�*_K�Ԍ� ��Ƈh=b�;�J/{���Ǿh������vF�;��ϵ�3�W�_��*e���}�k5�Z��SMcK�Zj~�M:�c�Tq^������m�0�_	?"�1�������#$���aC��+������u����0M3J�nCl�����vIɣ�!H%�.�w�ևC��ӳ�kl���W�/�w?A�x��9�A��F�Y}�xN����:-i�:�,à�(�f�irLƧ�Sx(�-ڑ�W�2p�1�_�f��.N/��&9jL]!͈�^�Dz�!�o�0s�D��=�H-.G���z'���s�N���+�3�j���x;���5֜�9��!����T����"��D�5���&nh��ԣ�,�	dr�� ܴy�Z��#6�v$�a�#�GH�әd���7D6x��3�>(Q+�"v����JH����5�[]���vZ��=��-2QF��\��B�a���l�!5 5���D��ݹ�	�{�"�NU��5]�o֫�}���8�T:[�c���?I?�����/����3�H���0#��c�9*�d����Ý��(ȘQy,E-m�8��:����ЗG!��ͽ�dJ�$��H����4S�C���o�.��1{A�l����9���vK7A ����"I �)���
?��i�t�<\��Wl��L�;ϩ,�:���r��;�y�ۿ�x�^z�Z���RR �4��|zìN�`��/�AL�I��|MH'Dh��s
'5���HR�=R�up�&",��f�1�7��<O���V�ԓ~�����Sf�˗��p��������`�v�v"��vq��
L� f0h'�
�� ^�Z��;�1L���J=����e����S�ad��"�gL��%�"/�:��~�v�g�1��|���M/o`��Z�5���%h!�T-5d�2�2�.���6�U\SE�R��ͥx�6�*(����?�0�����Oc0+. l���_cN�9f��<p����w��K�i-���l�T6�'~���ᯎ���Jw�j�%D'�U�N]�SUʕ�-���w��l�eY�.�n�"*o
�KjC�_��ͭ����X>n@�3ȳ};u�|-N�z�X��W�3���?g�V7���l�����2h1?=88r��D���	�mnޗD�=�(��5j�@�b^��w��WJ�0�i�ޢ�C���l\y�[�B��\演�U�S؂7��,U�8���$ϧ)�mn	�ʬ����!�+�*���i]�tz���
������1tH�[/������������T��d�rvR�H��5��#`�s�s�2[7Pv|�zHlǜ�Ʈw��E[W\U0&$��D�m��#VM"c��������k�9��
��H�>S�e?��Sz��_Nw�u'ݼy6�;�Z�t�=w�;��v��'>&��]��{q�J�4/�6t���
�5�#[+�x!�����u��ļDC~��&��cto0T<@�&)Δ�����H�^��#��7��<G����%3����c�Xl�M��8�U?b�ב�ӑ@ԏS�H��'�0�#����/ʁ���*l5q1u��a��ڵ�f�|�B��������!R
��Í�<���I���w#//�e������DoOt#5
�iߔ �8����?8M��C'�ρ׋���)�+��f>N&Y�j+(]tXKdɺ�j�u<5Ő
XY�Ig��:��R|�2���p���]�ٟ���U����J��v�#msT��?�R�4����1�fC��0�_� ŋJW�ΒB(|g��"<�k���������L�s�2�)><;J�{��^Ӎ�me��Qg(����6*-oˁ~�c����1�r����)�a�P�˺MHk������ޡ�9]ˡ��o�3;�h�F��=ozMi�J��W�ߍ��V����S6�DJX�;�*$on�no�s��������9�4��/z5v���֮-����^L��~��S�]n����'�^���5s�\�K�i�Zs�ͨl����ϱ�2��qI�R&Kx3�{��ٌ��8�����v���5��ܳĨ[�S��9M�%# #��ra�����z���M�:舺��b��Z����d��b�)<G]�}O�zJ�|��@�am�"4��>�W�;L ]�ސ�\���ZY���a+�V���5$K��Q.�>k�.�N
���_�����^O��m��&X�UH�5M�8��~�@g�bs�����|��������)Q-k@�D�yf�������P;NK��甡�nR��I��Hs٠G{��'a�B9�l;�E����9/��H�"�aWz�s�5b�Ȑ5U�ӣ�
"�)���͋�w�u�5�\H��^3(��W������G����W78�'gEH���n�r[����ч��� k��n�n�C�0��x_|jf*�-g*�a�m_+��Mј&���8}7>Ӥl�V�q]؁��9��޼�e�nl�+ze]�~-`�� 9I�����B�rA�dS�a�{Εj�4�Q�Tܼ6�1D��G�!�7�q���'k_��ؗ���OO��t�m`c)�n��qߝ!�0/�m&�l�T��� �7���_F�-!��S(�&�g���BÆ��oã�@�YI B�3	e�E�m�R�K�<�5��A���t 9�y��"�p�0�V��I�BlD0��1(�x�C��;�k��Q�z3����ԈL���fr����|��đ��{�-k)�E���<�]��i*6./�r�	\t"��pcNIx�	��љPBن�+�����os�?%wf�W�� �n�I]���J3"���bҿ�{���ӫ���g~�aY;�9^7,Wt��3��k:=�I���;>�7$ݕ�8X�.|򏎇J�ƭ�CD���'�/)(c�(�wq�P��Ͼ�N�7R36�R�M^�����������5b�ڴ�@�_����]dw�������$Y_Ƨ\���L�o�b�?����7;��{�Ы����/��MM����{z�>��OqD�*��Hri�Fa��tbb@ǫZ�t�Dce�4l�npe�`j�[D�K�$b�:!���M�M�"졿��ꊐ,6��I]j�:X��,��w/����tvv��uO���9��[��W��%^s��Q�B�Л��E&�q�y�H���p%�"��G���\��wƢ��!0�Vߡ�j�K�G��O�t��stp��Y�>��5��;��m�3?�S�]	�4��b�MYИ�T_�n���~�Ji�@��B|F�}YX\��[�Osߵ�s�KX��d��c��Y�Q���o���ҽ��!���v-Bf�3갓��D���NYS��uU��^�L�Ģg)5���HhB�A�X}�#(�\)lEł�wu�Q,��ƺ��<����&s��.�Q�m����x���'���8t5�?���̈=�׀мn�*ig ͥ��(�����,B�i$e�����=L3�]�>DK�;C���}���u�~���S���u�m�D���=����!�F�I������G�Qnj����duv2�Q�d񣓃3�}\�2������i�:�s�ӿy#���_���bs���3�8F�_�;,���6�m�s'��U�`�����ofo7��y���[���o�Ӵ3��q���M&aTp��b���|��[M'x!�}����6��MYC�x'���@._<>*��G�����;���w�Z+�3�ǶL�T\tOb����Lmc���y�;������Z��s^\�Xv�.�k��Ժ�Q��ܮ[��ͳM�<�ok�������(��o%�38�&�Έ��d݋�λFPK=G�;�Iq6��©����4}x���.�M	z
���q�4��vWI>֢��k���ljzVr�o�6`aj]�d;�+��{u�RA��`r�ݾ��a�?��O� ����c7'���:FE𜥩L����:���0P�vQ��͢�T�k��k����s<��,�ѝ;|��)�v(���k;�GB����b�)g;�)�|�E@`i��T�ooˁ�sPD�5�ug��)�z���6H,�-�-Q'Sy���E׺J=ۇ
ѓ;O'��h�l+�Wdmeރ!����Hk���㬃(v?�U�}ʴ��?�PM������q����G�s}�Kߐ�Ŧ(����z��D�Д:�o��Ā��5�%��
��*]��$��[\�S^��x��3��r�����4��qŅ8R3eE�ؙr3@���_�n�xۘ$4+�z��&�٢�F���`��1�08*~��	!F-���u��,�>��ͻK6�%�T����(��G~�^��WW��2��.0�_h���; n�����5C0I�E�����L�ZZ�I�"	 �L� ���Cp�@�0��>�2���t���`䪒��3���š���쥪9�\�&¦�4#�����#h!<7K�*x2�26�kO�@;�o*�I>�MX6�IQĻ����^�XOT����~����<qG��AxAg\k�av��E�r#@9dT��H�qa�Fy�/�p+����#z>,����p.�<��$�H}
��sO膂�>�8��O?�)&&'
�l��d�[�6��S�D��H��jd��xt�G��$?�+J�3��ʟ2<��p��_��u�Sjx�|�Ă� [l`���2�Y�� ���H�����"̩�z^N��H�5gę{v��g�b�m��:��5���`��RO��{K(�M��J�8�a߫|kN���N$��ز�7���H����ԧ�?�Y�,T�tBUSfoK��p�5�؈�|�!A�4�79@�8W�z�&�g��\V�P0ڦG���H?��t��D1�S<v��u?�A��¶���P~��tW��i[�P�	㞜^��K�<g��`�SC{W�q���,�-���*s�K�w
a�7�ƭ��mb}EN�2�]t��?�}蟿���C�a���Z��H��{]�|��q����J��mcW1���rQ�D���k����f҅Εk�֊��S=P��i{Ú�"�W��AOo~�kx�:�Mj6*K.m��J@�4y��'���l�Y�A�@s���N{9$���sLQ���3��ŝqR��S"�m�������g[ߠ�����������:q>���ן�^��I�L>1%�8�A���k'�I��
¦WzX��7ոi���۝�k-.��i�TԎ�=+���`>��*�rp �>�u�	���*����U=R���E�lݳ����>��t-�]�v����>G��SZ�v��S�B�Q�I%�����4�fr/F���v�'Vh9�-e���;!5&=I[��E_�`�ܢ�:m��;�O���6�ݿ赯�Fl[����������������1��:�=9O����Q_�����QsX��2K��.���cV~-�E�]#�t�ہ��%����:����q}f�z�A[�e��4<`K{��m��8o�v�mc9�}H��Hh����dS�a/`C�'�g֮��n��>�6�m��Z���>�M:kj����݋F��-,Ə7ّ�lѥHj��6�GI�Ρ`SW���	M�lP��5�0у�o��ɰ�Yԇ�~}����P�u���>P2�D����>7ZM��G��Q,��(r2��ҡ�y�Y�`A�đJ9�`������������K���z�WR�ܞ���Ug�G[`/�;u��S�5��Ҟ�������k��������;�l��)�F��,���[�l~�7�␅���@�P|�C_����}A�(Q;I�����1��$����ߒ��X*����i�`?5k!�b�uD'_Is&�z�u�ݬ��J�z�D5�d�X���e�[,�o<Ki}J���uL��q�LGDE��^Y#� ͱ�� �ű���}�����o��Aٗ��+7���x��[����K-�q]<��{+���4�w]X>qX�!,t��bt���w�^�#M0��&�ǫ������t�qk�O��s=wy�����t�XNsLocc
��'��>��Ұ.��'������5�S���л��=t����88������!��a6X�U�CG�m$�NKҦL�������Y o�K!���Md��!�D�GY�Yff!������ȑ�x��go!�+pY,������իw���1WRC5sZ��'�$��˅,-f�¨7��v!D�PF�-o0� D ;��m��'��^Re��{�t�)�kGq��0����\��w444ݸ!3,*�����akAJl���ע읭Vv��7s�@I��Vtzz�)T���o��@�~`��>�Wg��y�l詒�����y�f�#8�=�K�J-��;̥�Erud!��Y4R7��&-�1��{�<<��f*xwQ>(|�\gu��m�z����G��oӯ���O�Ǉ�D���=P���/]�5�n�z�p�Tt��2Un�XG�=��F�T4�Zb'�1��tj�I��G��b����6\��XfꜸ�y��´�[�v�cWݻ�7u؈N,�RhR' �b�}n���$rO��N�<�+�G�J����A��_H��ז%{!�.�8l�?���9ojMW���hz��^K����cM�S�b� R���������%���f6�����=���Z)a����&�ޞ�=��T�:dO�Ŧg���k��)k?�tx�б��W�߼q�Q���1h޻絋��:�)n�g�nk�E��Tiu���'��!4�҉��5�^ �{t��d��Ƃ!�(�^�-�R2jA����IQ�A�oY���t����پ����}��OЕ��������]'''t����]�MO��ۮ��}�o�4Ә�Y �;�	�'�8.b�0�ӱ��܅p�v�ԁO��隡x?�z_��p���ۣnaEp^ǥ��z���~z��O_����5����;��ˣ�K�e/y��;�$[���D+�[�9?)��:M�N���f:T�{
�B�]lO-bT&�ѯ̈H�^��'�������rG���dUC��Qzn��F9����f=�y�e=��1�A�q�8/�j�o��Z~�mj$�,Nu��σ��u�:�W#D!���`z��tv�����`}F��$yj-�9\D��3)l(%99��n��8&�Ş�5<U;���ɩt)>ܒ�������/��g>�9���Y:u�Z_��q��=��o�`��=�_	|x��S�4���w&��Xu/�0�zU�G��@�:a��$�1����|=��h1:��'o��-gw]�m_�����0��(�t
�2��}�.b2��ȡl�ŉK���������?�_Ҿ}�i�m��t�h�ȷv#�~�);�9~w��^�����TXu���T&t6KL[��y������]�k��z׌�t�ҭ\ns%�7�smk��	?����d��⁈������NO�����_v�yk�uh'�a\�c�v3Z*�wx-2_�s��{�SF4y���T���3���?�Iz����Fl��w���G����G}oOHخ&Y�K������^�Q���F�	�d�WAG�8%�+3l��8�X�q��"�Y�L;�SJ���}��{�bD� �Z��`'�ɗA���N�Q=ى�:�g�),R�Ч��$�Ɂ p�?�@cχ������T�Q{�����o$�k]w�� с�ue$�O &6�{F:טd�q��#ۤ�pBqw%�CR����A�,BCؿ����!kM����
���"�!f)ؖ6��t�R�N=)�{1W-��Ȟ2D����YP��4L x#���PDaM�ZL���nJ�b�H�Ety�����Y�#���(=�OJdݺ'Vy���7���ߣ'��.%q����:����ڶ�̣ɵ��L:���+p"��v���)9�^�����B�!s�ˢ��X��Bn�i@�h��1f���M�	5�G�Pi�A���x��:� I�8r�NO�N����N+��Q�?/��2ӎ�J	��[`�p��7Nx���
�f10�:^j��\���j��{����O~�~���._9&q�,tZ���$v8At�Ă��|ұ7�b�I	����Ĭ������aV�_Ø0�q:_,���- �"�l*��%=��v��q�hO�Ss�s�� l��{��s?�2Mf���b�\��>P�.��������˾���`T���H՝I���ҜYɸX�� �x��P��ǌA�c�'�h)6� ` �8�T*Xew4Xu����k���J��P�py��ب0X�E�1t��r���C��s�D����Nצ�cz>8n@���=��,9�;��Y-0.j݌  �#��ϓ������Ơ��2R@rE�g73v|���8��?�ē����8�<�B_�~H}�ٵb�F�H�7����Bku&���b9��Cʷ3!���+�h�X�u�:��E�Q�HH�$�HD(� ���o�{�/v�f����s
6.l�)Ȼ�^s�_�j5���ֹ��7���w&��G̰��b�JC����ʅ�O�`cj̬����Ṿ��&�i�����Åh�De!�<���٨Se,� e�c�}�kY�WN���~�|�'l4Q�;H�%�e�`K3�v�8A��r[ ��=��k�ڤbI������D���*���-q3K0��`!�0�̑͹�7#o�81��5m���6c�gL�m�2����۞�נ�����6p��Yw̬�n1 ��Dyg�gs��S�U�Hrފy�:"�s8�~���W��' (]����`ㇳ�!�s�7���c�}����/�?��������G},�;�����O���.Ɇf����u�͕̓�V_�q�m�u��箩�[��i;[٤��o�mnmM>є>��F%1����Q �q,�v7}�����0}��'h��\nY�9��Rt���=P]%IJ�Z���ꕫt���8�e	�Z�lu����T�,�/�s<��â�.��.�c�/!t�ј=�s5�1ӵ�%� ���Z�s��S�D)�hheK3�t}��*9.$��O<1��� �H5��k:9=���!cȊӉu��\�8<��{uZg�C�����Y�s�K�+M�&I�@S��Y��+�L(ݬ�*SQk_�uJ�*�,"?uY����Ӳ:����kFVvD��C�ցWT��Zv���|�)��=FO>���j+U�Ш�T��(�ش%���6T�Z���S0�rNj��-Nv���l�;OY7J�nޜ��Or���N�0%���ƌ~Ӯ)n��V��l�ގ�����ȏ���V���FmQ��ixw#�?�6�)�)�{��v�r4�K�ӱ�,��7=��f�ր�v<��!�iv�%u�ſtwm�7��|F��]<�`�ؓ�g�F[fӖ��ߊ��+��.�B��}��w��>�ڇ�wm�S�s�����\|�v�cR��D���p۴�.�ϛxQ(c
U�S�C��]Im��8�@��pz��o���J�~M�1�}:}�~``�U(�F��4��P�ڮ�}�i��_����?��Tv��c$N�����n�ڡ��vU*��T:���0gk=`���-���ս!�>�:Sn��Ct��bM��|2�j����ay���q��8~n-;����-iz!������QQ�bُ��v��K���D��}]�1z���eL{�uwq��;�v���^��ԍq�2$[;IJ ��Z_a�:�k�LMz�\7�!ǵ`�!`~2~�t���D��r1�^�Xg�ݕ�)�g:(P'¡Hj���]x�8�cv��3��ܦV�$2�J����s{rM�bz��y�la-va���OE�\������s��*lZa՝�^}ۢ���+Jѽl�����TR3i& .���l��bϑ��N�@�ݐ�:�1Я��F?���o����C2U�gǏ^�4��ɞd�rt��+a�<�+��:��=��7�Ob��Z����:�̄D@�G�w}z��;*I��dx�8g+���d|�}�#��W.zm`�:dO�]���K{��J������AM*��j~�}���L��(Q믛�����%ڑG���X.¬N�V�%��%�ԍ��5gV���5Z��H`ݴLל�$]H�A�G"_�@�@[@��pl��>������>y�
F����c����R��b
����Y����!K�0�h� ����͍[i�_s
���F���_���@�D�v��W��/�y��ʪ: ����P��$�r"��W�ٌ�?Ō�Esc�`�� 9�j�kb,�"_��a�Q�q�XD#eJv��q��ܡ�f̰a�>Gы�"{?o��!Vj��t�bT+�nq�bCj���O�qEв���	]�֔�"�lS^�_��-)9�s�� >�����L+�9�R��E:��!u�)��8�8���~$Qo����e�6Z����]���7nҒ7/�V�>��<��U�+V�_'W��na��v4��U�4Xu�Iyu�u�@a�
�k���YX�:xP%����4,����Z،�vIvk׭}ȑ)}��v�o׆�E.�#����5��m�}��fZ�)�F���v����&͙n�Y�Kk���A`��%��0֦��o�X�ҵ���v��q�R��JY�ڮVg�����=B����ة�z�W�����B�H�.�ҋ��1�m��9����0����Vy�՝?$�("ΏڥԈ��:�m���z
�pįx�mx��g��������c57.sk�5s��t~{��07d�DNJ.��$�����I�Z�XhQ�q�:n&q&���7+�W�5���W�&uuK�~�Cd��ƣ�L��Өh�Vϫ���:�� ����;?��oq�Ι�\�J���'��c�_~��|��>��s�h������E���]/���ќ�'�"�NuQǃ�����N+�Bs4~�t����p�e��a@�9��S�O�gw�C~��{���G���Ɉ٪1���)]���O��!N� \�7=TǎopN]�����+�����M�p�������-f�!qЙ�>iV|z�������9*�;����93������"���:5m���q]��� ��Z�r:���bz[J�S1�sj��ɝ���0AWi�șW�H�5�n��A�r��4n��	N>aC�]2E��
"`yy�s�CG'��Nv(H���D�n\�ݸ�e�_�I�&�ڂ����Z��4�g6�׍֫ss(�#|��!�s�Ť:��t�HW�FnVMQuc%�
c����G��u�+��$�t��~rS�@�?ٷ火�ڶY�ۚ���(��s:�y��\��%nj6�mG\s��2��ض;�}��F'1��]�:�nm�g��������\�\���&$-v�N"����}��Ԓ3��`���}l[�4Y/ӟw���7�Z��l�g"�؇�wElȟg�i�:�4��޵g6���թn����w�b�G+1&.����'~�tf�Wٞ�l,�~6��g���&��Zgx�h5bU`R���wjP�5c�!���~�G�kI?��w�w\����(�f>�V���M�-"C�>��d)�~O�=��� �� dN�@ݺ� �a-α�M�XW}�a��1d=��~��#qeagRM'.N2�������Na�a��^���d���r�ͺ"���傀%k�$�֫�q�\�e/�vY��Ճ}5jz��F_�����mǑP$��&�U��Q߂��;t�k�C*�e�uѹM�(. ��\e
�J��fa��E�)N�	kg��\��j�M���ht?�%dR�S^�������qhuR_1���"HF�M0��{��')��B���EWg}�S���8#a��WO)�v�}����t��Kz�zU��^�p��e��d�z��#�-���r�{�w8~^���C���<+t���pz!����#��h�0y�-���C�q�nޤ����O��_��>�,]>:��);���:�98}���Uqg��6��>��(͑��Q��݄��w��yZh%옢����!��EZs}� 4$î���u�}|��=��y{.��X�O�b�-p�����5j���d w7������TP��Jz2c�t�{60�U�p�2\�B��{����hq�CT������WK�$:���Զ���sbl�*`)�6<��
|yC����۬G������V�L6�W�p 6a����dF5ǧ#R��� �Q��Z�o���D-X�H�݃H7c7+��iC�Ղ�P��%a\r�D�5ǯˬ{ڃ"�b�`�_e;���8N�X�X�	w�iƞA2BM��bԋ�1���>fa��j�[�ey��|�g�������đ��˔L�����\>�r��L"L=q�k!	��h$�ߖ�F�� _���8>2�d ��:�a��T������E���\�!3��+v��Z>��0�oA� �j3�&xE/贡X�l��v(�L
v���|�\y��5E�K�̂?�c��セ�Y�0����y! "���H�6�� QJZl��"gc]�S�׿A�s�Ry�Z}��T�}v��~��^�"{�SL�` �X��6Q4?���ɯ}��tCr?Y�_[|s��=O�ϐ�o���"�J1'H��}�(�H@���O�1|N�1g����۴����&_�nÕ&4�\��a�:�w�}7���������]�Ɗ\��*q��w��*v�}���wo������(�;�; d��I#�q�^e���̹��ޞ	�K�Ʒ�����1^GGG�<X�B�4"\�����۵ٔU~��挫/�f������Se]�b��O�_��6��鴢��!X7���g�#���.����tǃP?�6ݥ+#�u�q.�_Vk�F�R�8n�W��ħ�a4�Ɉ#R�M����C,���e��˞���A��/���}��:�p���W�����'?�i�x���<EE��I�(�n�MvT�<�FW�X�mZ_{ͱj[:i��v��F���t/��BI�=��M:x����:����%�9��Wk:]gz��h�N�9��?���`�i��W�N�pD�qе_����o���$����0�KX徝��kfFؗE��s@;Α�F�T!ӏѼ��^����{'�.:�sy
)�'|�@�������iQ��@/����s�}���e�x��_h�m�����o�����PI�g�N$?�Nd-�SSglS�~�$����:͓��Z���1�Z�:NOY6{��Ϥj��I¬��4I����+�'/#�%��AE�M������JN�:�Auf|⋴~�+t��u*��j~�-c�L�ǀk��D�js;Th�yמ:�N炀'�����(+Di���l�Ķ1{m�y�����v�n�p�=���|���c4k29��\��9.D-O�>m�nX����N�x���\ �Ssk~I42v���mы�_䭑�8?ٵ�6����lZ`�}ۻ�c³3x��\���xE]�x�w���wM���;��k��)R������:dj*�����ܣ޽>�Jt|����g_�e��\��-G5gI������	r�t<1_8��`Y�.5�bi�0]u���9v��(���O|�~�_�kW������h�5����bp��:���hrŜ�#[�cp�$��2��:!6Cm�Z��9~
�P��a8�P�(�ǫ}~P&�6��>��Z;����.�O��,�
�`m��[��F��tn��\D�1%Yi�D����?�p�����f�|����O:�/�W�%���Mm���Go�}�eb��;��$��=���h������Q)"�m�^ě�u�3R�ˮ;�#Kp6�sC̘PB�� 'K���Pvx".�}5�rӱL!�Ap���'�#N����aR�3��ҕ��)Vz�B�A}=�ZkA�}8�}D8l�P�*r��2'1���2��ܞz�����l:���t��o�a5�qw@p���c�S4s@g�!��zYZ��w}#}�OY��x�Fyϧ������4<������-��ђ��N�RM�[�G�#��Ɏ���K�X/&8�[麸G�ˁ�`���>�k@jDn��-^�ˠ�y�5L$}yR�g&�L�9��:E+��^�����ѣ��K�x�W��p0.���6<
a��	�4q��hx����跖c�I-�:1��5Ae�#_�b�c���5�D�����Zۅ�������E/Q" aD*V~��9�F"Yfb�#�Ft��e��q��WV��HlH�N��^t�f�QL� ,��Y?'#,�ԛT�P�)�2쓁RA��eR@����aA�C�p;�x=���)����Yn���Y��h����G������$h�6�i=��:5��S%{��G��Z���

��6A�;(z��H��x�{�^QT���F��ڂ�L�Di#��%�	m�]Xq�$�		������Q-~O�3�n�T~��T3r�����B��Yӗ��5w��
T��X���Hk���oh1)�B�Ľ�h�я��mt8H
�+o{3�/}�n|�St�������W�pv��FR�K4��ƺ3�m3��\�(6Mv��[�:�_�����^8��5� ��k�eʦ�}�g�<��hm���`H�z��=-mGЮm퍗;��`���ߺ��õ��o�l1�J��)�4�X�y�|������_��_�ǟ��<�iI��І:JD�"�F3><���	>'�eB��"�u��_9A�����m�ARb\(�g<<a3��/d�}�����^��5���lE�<��kj�s�#�qMיӆ��|�N�>Vv��10#VU�I�n�^.���-x�.�����C��s�\.E��J��CX��N/0 %�N'o9o��F��nB�' s�[V��T��w��tu����������V#Х;������Hi5�ú�]+��_�$wY���9�xMe��qpn�[�<�a��m���9 r?���N.�a���gqI��Řr�s*�!����t�������x����8�[6���N�Y���R�Si��qx��z�[��rq&5yɍwa�F������lȻ���X�h:����M씖;��s���7�o�^��������E��>� =(X1�pH׵�8#�gV%�.�+�	l�'�P����`p>��R�۞&�Ѻ�,��lS��#X����=��ڊ����i�u��ި�C���E_�v��{V�!1��fԱup����ӡ�:� UC'#{ہ7�������=�F\q��_��/?F��'i�O�vHìC���p��Vt�mr�\9��i�ϧE���X��G���L��Tw���������#��܅�	��,��ئ12�l]E��8���1a��sp�Ł.� ��7����%�c:�?/]��KxHg�$��	X�-̓/g�5#����D�x�6��SJ���r���\�7l����MMTn����.�ȥн�ʻ9��F�^i0A�ƺg����W��hײo5�=�� "Mk���o�٣Ny��L�z���wQw�
u�:���D젩A@Nƍe�)�Gqmc���>ͥ����`��a]�``�xP#�m��Zѳ��^veG�(74rQr~�S*�N>��E��|�@*jS Iy�$�G�Mq������q���S$�	�00E�E�0d��"��W�7ߒtr�lsD�w�m�{=�ǑD�L���K�������4QSᔍ|��j/�vJI���G*������jd
��N��
Hݢ�\!)ѓޭ<�ژj$���Im6�:NpTsv��uW��q����HY��/�+���(1��3
�u�����NRu��S��ʢ�����ƾ$� D ź�ԑ�ozyq��v�vOXֺ��"��D��{8�l����ٓ�^j�!�7 W'QK���0�ay��Ҿ�Dm#��U�I:β�$�bR'�N�W��T�	�~,�CĂ��q��|�P�~-D��e7#�0���,;��zѽ�:ϕ�+��Z�����gi�������ǿB�����J*��#�r�A����Y>��U�O�lԵk4��z���o�͹n^r�H��6���5H
�_�T�(-��F��Z�~P�T���CBZ��!���묧�;�+o�.:z�kiy�ts|�3�T`5j��T0)��`/��Tݣ��ֳ,
��{	�6Dz>\�t��*�	�Rs��Y�cf/V��ǽB�yGtn�p�I�	��c,L�7U����+�� �� �_t��j#K ��1#ٕ�4�O2!��t�p��g��Z�J������`���mJ�~����n~�ܓ�4|5`�����"h�HA�.�I8�����������$f/fVf��O��$�!M�M�n�P��[%Ģq%++#��,�2q�6����7~��8��
�c���陻ڹS����sam���Q$�� �DQ�/.� �
�����Ȣf�=��!�"���ug�P�evJ։�c��^�tRI܃w�G��ӕ׽���'���'��*(8[�R��/k�Ϝ�����ۻe���@��mלC�y��iǆ�����.���l�g�J��i6��ixR���g�#Gٻ�g��ȱ��6��щ��]OS΅Qu��Ů�A��uM�.�*�$��]P���>_���o}��������~�'�
��gԏ��0�Х�c��r+l\��,�h��fDs�ZO�tR��U���9J�n�1w���m'=krB��dLT�d)��C��"�
�.K$��˯Ƒ˗�9G)}�.�j�+O|�n�8i�Ӭxv�Oy�đv�ʋ^��x"6���ל�6A]�c�s�����Pe���C�~�:|�w�ݯ5�{�nqL7k8�a�kVg"s�	��KQg���LL���k�O�H�$�z0�`�Z���qj����dT���h5�l�I����t�o������|`Tk40�	� ܛ<��Lg��rAO�(zo�{g5L�#t+�v ��e����eF|��I��P�J%v�_d���t3N�[���������x��Uf�f5������	�X��a��K�{����8<
d��.����h��	����4�������l�Z�ZZl�u�sm=�&1��֞<�	�9=C=f.�IQѓ��wD�C��H��5]`�-�P�{d>mN�a��t�̲D�;5��FU�i��bc���S���s)�J�B�K���1Zd�4�݀��p-[�>f���y#�Ӱ����Z��j�������E�o�a���Gv9^�$��:.�Se�8w5r�i��w�Gt�t�5o�����x����ߠ���5���X/�� �a���<��胶^�,r�e&�oo9hk����i�M <�V�{�S�⼚�:m-x��M�Q�T�/i9�[����p��ӥk������u������Ϧs�������Ο�}�K׋y1=)�vݴ8���6��a�d?o��̼n����"=20;*A��v;���h�
mY��5=����?}�0��m@��׹q0�`�)`�PGF:�M��&�㻜7v��m:�c?�ڰy�&�lN�r�����W�[���x���=�Lw���������?D�Q����k���?�4)j��B�co<�a����p+��鎁8���`��,��FܷZ5ke�H�H���c&_mo�I��6��ʵ7p@��$���1w�����|�C%h�~�r��.4vǚ�(��Z���'/�C����WY0��B՗�Wv�U<�kK4}��®3�
��g8T��\�e�N�Wh:xs����v������7*�lx�P�FX(}�Y�����e'��+�3�_}\��5��Ni�q��[���8�އ�0{��(�Xj�� �c[g7�O5���.��������В�{����S�\��[y/��&�n��{����Q��k*��0�:�f��`�����84��,`ۏ��[�tn>ȶ�I�4�Ī#QDP����VW.Sw�]t�ʗӕ7����u:���髿��t��`��G?��+�X�౑�'8�wX����<]aj_��s�a~דS�>ז�Ξ��rΘ֝��BE)xw��V�3�F�U�-�AC��o�� 0,[���𿳁�u�;��V���7���%=�:ㅐj�"��I4Sf	OhC-E���d�`��K�;���A�mX/
��؈�V�w�Z���[�8<��Z�P�:�zY��w[�ݲ�zj��Pȥ��>���CJ *B��!���=5�=�!nu&�<�� /<�#0�����W�y <�L�Q�#���toe�<�����ii�S�I���[�d���G��������V�d��c��1���.k��T�0d��C���h��)�A�n_����#65t��?���/)ֻ�J��4z@�ܢ��>9���ᙫʃ�b�f�P ��zH�s/z����� �ۙ�5BK��v��̋�c9�#1� &�׉\��x���9]��z�����t�ַ��?H'��{����]F%nX���W\d�6��>�k}����D�pG���o���s�/)|Y�Ôo�j��7x00o�i6�mڳ}�x�v6X"��;_�2��r=r��%��uF��H�\�Y��}��u���sQ��`Js���l�2��$RS%Z�W\�����瞥?���k��+�~��t8b���n�2��`n���ą�ha�\�>$�϶�]v�V��*���&J1'��N�>�6���'mߤ|���,���K�n�.�ݒ�ֳ�<k��}��9Y�sm4t?��O ���oײܓ[�&���e��j+���W�D��s'����壯��;�h5����^Q�ٜ�V�ٽ�uN__��u^���5����~�N'j�;����:yu=�VR��ߏ��񼤻��V��|����XU�����p{iOvPBB�3��o��)���R��ҝ�ڷO�L��F�F۳�*�lY�KV*Ǩ淾��_E/{�;��|�e�XMN�e6|��#��ܬ2[�"R���)њ�9�����%�s�~]�:R��n�j�o~�^�6���J�9�|`o9��l^�1���L���F��n�5�w��g�Ӕ�QW)�)��r��&tΒь�V�Fo�q~�ٞ�+��"��嶇~�&�8E�����Oq��n�r��%�+��"��i��q����}�N�`sk~ol���Xo����
xj�k��\�F1��<���%:����=�w�W~�����/Pz�G��값���t��}j��1�2��s���X����SZ���lG�<]hW���E�vN�l��)Z�VZ9��Mlc�1�bB�4��edE.k���?�Ͱ�L�)�T�U�	emc�*����-~Y
�z���{8��)�4|'ANǒJR\����� `7���	o��������k��&��C��F��}�+ɰx
��h�j0b�m����ĝ7
�Y]�`�d���'�s�l�k��#/���u_�k�C�}�����?L���NׂuKH[P4�A����I�sm�	_`�C���B��a�1l��#�Gz�ւ�����t�0���X�w���^]ns��A~ڦ��ǌ���0 nw�s��s>мg���aӹ��4S�i{�c�%
��g��i�5��S�}�W!�%��-����r��^:e</2��v��3��	*>�6v�Oj�M�28l��ǡm��.�v�;�@�)龧�l:�9ݓ8�{���2�T�q�KzK0y�(d���҆�u�/شK�1kh���1�}lM��,f׺\n�)qޒ\�t�>��L)�&��+��~�&5<�Ӳ��*m�o�"Ї�%�}�=ʤ�X�3���#�]�|��ҵ{獵?�a���cT}=�ي��D��<��2�0�vx���ky�s�����~�Bʧ����[I�rۮ�����aNӉQi "��(XHEO$�OUOo�Ъ7G�}��0�{=��T5�z����G�9s>"�Ukn��O� � ��R� � PBX���IX9��?��~R�e����k�ɠN��%Hܠ���9��L�sskf��o���$�`�tn��/;�`�pX)�
�o&�Y]l��k�"�܀�m��P��.t^��{��wt�&X�r���^�g/����a�* /IѠ���.2�.m0>|���g��^�G�iq^���S��������VM	�Ba.B93T��6����o+�Dٸ��tFc|�+����p�ҕ�yƟ&7"��ͳ���ic�g�q���z�S�N��8�xLhT��"G�ۦ�,
sʴW����偆�zn�{��Ct��w�IZ��o}�����B��<��A�]��p��(��@�s�w�����e �w���\�QA��%������r���z_4 m���a^⳥8�C��Z�(H�"��qc
���m�~]ޘ�ɬ�K�F��R\�)CL{V��e�9QƂ(8!P��0�$���RO�ɟ�s����?��~Agt:*&K��B�0�`�f�-�1�Q��mY��$���$ ��0S��r՚�V'�fC5a����fT�d���7._���5l=�S�Nͅy��3�v�	�^4Ul7�Q�q^�ڵǩl|��n�
Ow�k7��F����̽�?H���0�]���Z"R�X^����參����޻ݖ\�a��>�|�w_sGw�4�f$F!4h`$H�g0�� ��ġB'&�P���+�8?R���)a��J�#��A�$l�K�`�KI�y�����޻�{�zu������{gF�-���٧w?V�^�^�\���V?F��<���Z~Ó2a(���pZ3N,�*0̸L�v��x!�h�S��!W3��b8rt���M�-`��p����C��w>��πK:��F�}��S��e�N� ����ݱ1���v㬖��E|���m������-A[�nL�t)!ufH�"���n�}�qX���<w�[P�n<l�k���p+I��0�_2l��k�-:��[p�ל��j �����΄��}$����fD������;c!�=	c�#õ�[���U��+�/E����	n�����C@��W񍴨��*��e�� ^ nubm[pSWx��.���9�QRT�!/��Nu7���_�;ڔ����F�Nx�tK�.ėԕ�K�/��Ax��JķR^�.�=E)NU���:
#��k����тȚ�骯���6ܶ�֬��}/�{��7�>�!�}����3>(5�lœT���Rr.�ߧ��Ti���Ԗ`�%��ݝ���<-)��r�m)������&��b�ϩ�����щ-�t/�\��Ts�X����^��^��6A�_��R|�W��8�A���db���6�n�].<k�_Fތ�z.�2� c�<7v�T<�=brqy�Q���1;���vp��N4`�D�SU-����ԉ'~v|`�(<ʮ��õ���}��Ư�Յs��z	u�����mh�;��/:���t��ᛍ��9�qKm�DʗE�����K鯤�q.b�8%k[U�_x/{�.Q:�������'H�l�g�h�Gn�C���խ��IT쪰/��i����`h	�Y�8aeq�!��f�M���a�imꠜ��g6��� -����x��n7�#�{�8 ֍�����E��vN��\��־��j�W��{��\\IK��%"��D�ɼ�OA���涶<$�hd	b4tO�X�Y��}�<~Q�C#��u�@��[L�b�����X�Np��l�魾��g�/�%{�A��xt^ik��l�a�������� ���O���O
��i��TwR��yw@چ�,f�Y[�u�|Í�;�b�eoO�w��5
�Ӗ�e`����}:���s]��|.}��@{���
`��-6f�HL����mm���O�;I
`=+�ѓ��
1ԵلA)@T��;����+ڑ���h��6�lT���(��r�&�B�а�V��Ҁ�����On[�����0H3���3S����3���+1��L�
zx���!g� ����"(��D!T��@�C�5v]�v�s�+��6W'�T]�3�#.���n�g��T��yT�o��Fs�3�W� P����M�����EoP��7[{U*�ԑ�W2͆��Ĳ���Ey�<�*k��!�+s�)0]�;����A�c��3�
0iӮ�i��옲\�/]jx��~b\�,���G�0$\������������p�����as�9��#�T�'d�ށp�(��9�Xe,
���-��)�I�3N^���U*��c�{�şoZ�t�}��*$'x�0��p�`�Q67�3��*fǤc��z�Vh����/�<��LrS���\��Bb���(������j�Bܜ�(���W+"G��%�aBɢ�F5ȫ(4B$�}��E�l��������������gz|����!r��Yu�vt~6��O��;|�g.�ń���7�A�*EU��?g����^H�#�ۇs8wx �iz�m�_�z�t�������f�V�L�����&���h:�JR�oQ.�����ެH�[z�
^���Ŧ�����"=�-��L�>�|���3X��{���
g��pB�n<\#�pb6T�2��g����j`���˚:�V�Bһ��ѳ6�8C�n|H	Hl��y�MHcP��#x������|}������ �$'��$*�8�-?��f�l�%�tb�@�S'������q�'z������aƄ`�[�p�﫻}�x������@�bz��m�rD
��'�
;���"�D&��i0�H�t/Ќ�r��4F/b��1QC��و�k�`�"Ƅ�$_�3z9i��"Sz},$(�3���Uk�O�� ���f\�2+�Qc�3�J�@�#�Hr������Bp�Yz^3���EJ\!�yC���򳈿q��֜�=�M��l���%飮(eR�*�Wj���6E� 8*�b����~�?Sx��������\��k�솎G���!=۬�e����/������GV0{�30�B�9Ge�"�6y�s�Ƅ�)-����&��A\��u˻��@uu'�O�I�����4���Ld��on�T��U~�RR����Y�9&�� ]# L��y?��1O����=즵�N*!��u�9�nS޹%e[&a��26gY�t�y��s\���U����/��W{�Վd��b@�卐�#��{���9�%b��vO�\_��%ŗ�����0��}gl�f�E����j���țI��(�2���V�"��̖qv�,��X��h�s�S׻�������;�ꢆ�d	�Mm�B�t�sA�T7;A��f0�%by>�r��l���t�n$�H�Yի)^F)�E�_�o ��3Ĥ���p%���E�1;*2�a���&���,h�����g���e!8
Ws"Oeg\qn�������`�\�-9�&@F�ZI��Av&p���h�V�b�KX��7�g�\�I�|E֦�u=%E��{b{��M9�\�K�Q7�2���e�$nؐ���]���W~�<昆�Kˡt:_�w�]���~#���$N0��
�:��NCː�"��YTj_bxߌ,V�0�Õ���7""	:��@}Ͻp�{���+���O��pVٶY��B{��n�$"���E~߅Wc�1�3I���ʾ�A2�!}�s~!S���c����.,!~�۱��Y���S�u���~sp�y��p|��Í$�F�3əօ*ΙKi^	Z4�V�/;�D��x���%��]��0�Cj�E /�}S�*C$���y�q��⳿�� ����B ��x�ICM�E��ӛ�\��� X���w�9#�X���o�H�ً��a��]C���O?���A*hD�?��.���܄Y�j��K6;�k(���e��� (	��֭�e����G��<�0�~�q0�]�	c���uV�ư��q�o����	W��vA��6R�0>�[U�O6�P-C�qvljiu7��L��UX��{q�q���WaO�W�N�3��:���8��n=w�8����ի0�Xw����� 	�³� ��m,PN�S-*D��k�@�ΐPe�gc���"�� ^��?��իc+mƊ�>�f����H���Z���;�Q[&�:wj�o�X���]����|���dө[����6mm ���`��-�o�ȸ�yVH�X�4+X����w~ ����\~��!�&��1%�;��o��/�9D�=w	6�"*��PRR��� �W�O�
Q�Y���E�<�Mb|��2��������z�!����M�>�,��!2�,揍�1v�Q�.s�w����7�eP2�H�x���a䧔�����P���J�'j�3x"t�@C��w��/{\�gдk�i�����8�Դ�6%��Y�RL:�EI�����]��f�}l��Jy�� A�+X�HzpX�����[A�-�7��z×��������8�:�
QH60�U(䷀�I�D�w�����]�[�����eŨ�ͭA��@��R/͇��	2��������Z�s�`8چ־�e�oכ��69b��IÏԖ!;7����[�>��w�w���e�K�1�I�"��8z���̀���f���~�) OA�����q�!��:�a����h?�8�&^�x?��Q���b���6��2>�<��}�̳��x*7�-|F�+,�M���4�ث�&(��7H�Y���� `�ͷ�t)�E�y8]�O5��m-��eϺBZҎ-��|p�p盿>�Ͼ چnG/�=��5���qǼ��[yk���&�Ω_���H��I�so�3��a	�P����	�-)�f�)ꌽ0��[Y�A�7!���ȧ�·���� ���T)��g���n
;t;h?mA
�|�t���_/�rkg�P&��Gp�u��Ň���,s������Q
�����;0V�}�E	K�3E�$0|6��8�)��wVڇ�޷JH�޹��㮼#�
��R�It��{+De�P��>�nf�L���z�v�up�W�^�����Yp�^���"�xī&D�Ϸ�c���D�ڱ<���2�s�vi���Q�8�gs~EOh��zC��]��1�G$�u`�x��#���8h��]�����"O�Ο�x�e��d�)Ć���F�N�L�(�N�q��x�gx!}�d�ŋ9b1��c������%���ٓ��=��+�b168�Q���0�/IY��9"#�������3PLi�lF �h�ضLMe=v��"��o�� �x�Kl��s+�wT��t�=�;�o{�. f<e:5�Xm:�΢%{�l�
� �R��IJ�������*���XQ�@ŕlx�2��T�}��z�dnf��������bٯY��?Ȗ��]�����N�� X����|�ο�mp����?�r�s�^�k�洄fR�]�.���_Ƀ�fn�I[�ҳ��mw�?��I���ޭ���9�af�0�	b�D�H9x}����A�Ĝ�!OO�6�\|�xݫa=�v݀[�q4F�$��A<���ͯ7tlq<Ť3�8k!��I ��� A]90��z�e("ș��1�y�ڙ��r�%��/H���X����v�P7Z.9>�͗?���8�s3���`/+���9Zœ�_?e�e�43e����rdn�`�a��=œ�7<�BB\�ר�?qܻ�'0�>U��DE�N�f���\��*�4����;�Mƙ��ޔ��q>b60_[������q�^�;����@�ʄ�Y��c/�&тx\r�:�(K�_3k����cX��fׯbF�Dx5��H�k0��Mop��{Ec��DpN�]�%����U.{w����~���SN߲�0���D,����ocB��x�ӣ�h`»�n�+6ao�}˓\���_d�;�:��n<���"w�i5�Ӗ���+�a�Rm��x��̑��v�4D[{�ج�p�}w����{���Ο��\]�z����j�U�x�Q �%�B��5�9�Y���9��Ӵ>��QYJ����v{��rF ��C�O�%ϡ��������H5���p��������
��6���f��2_�����aV�ݩ��7����y��;U���q���939�?���Q�UՖ�V��ʙ���2�+�X�%)�AY�t�~����t���z`����6b�"7#���ӡ2Ff�9�d��N`Ŀ;6yO�� �~%�#�=�hp�d�P�t;��ͺ����ft`�\���g�U_�.x�3O���3l�`<��j��j�ќY�H,ƴmd����^�s�d�H�:^&��O�Òot���(M֮0��H���}p�����z'\|�����	��S�G��$ur���P�{η-ZN��9�%���ow���{��l�qeW��v�i�?�p��]r0�fĦ!�(nG=:��Y=B��`�q]�Υ�+ ��a���\�ӷ�o���Ӌ/�\$C��(lA��Q7��H�$t�9��J�V�a�XQ�Pfv���G�!��<*�Q1r��P���qσ�kA  +g��į�%���V�,~�O�l>�$̂!�5�[;�5�O�u�]%t%�(��<�w�H	c��Y�7�$}P�g����9��C��q�B��;~��]���L(�mY�1����=��ۍ�>��yd��:�^�3��)4G�ʣ��Ь�u�/��閖[����/9sO~5).yj,ON��1��VS��@�~��ZWtOu�1B����@iH:�P��u��"�z�ښ>х	rK"�)Qw�U--��ޅ��CU�έ��rB��9�<ߧN~ ��<�ˋ�_ڤ.���\��m�_�ߎ������3鱇�{^����r�aT�3@�����!}�������2�Dv�&c��fd��rl�L�?���i'���սWݟ1 Gd{�ӦxW�x�Z���;�	����!և�9]uj;%]5���:W�r˕���}�߲j\'���{����}�(+����M`@���E��������2:!�����"RZW����l�U��ӊ��r�����y�G��_l��2t���S���ɋ#v"�'0
�L�F�N�E/��֩�b;�2���q��wf��3'�*�����xL���]c��o�����뫨k��飒�ʢ�������>ߋ^�M\��d5���88⅞�80X�oD���ԉ�ߵ�G���'��`e	�"Nݢ��,D|�c��G~��Kp�9y|�(��h�)_�Fh�M��&}Υ��"�ɢʅ~cKa�^�� lK�%eo��%cr;:�Ӗ��sr}6�CF/n����K������G5,�+D�D%��X�$F� 6����$��A�g�S�(#+f�e��@������
��N�I:t����W��h[۽��ύ`#`+�TP�3n�ȅܱ�e�YS�[�hn����ɝ=J�m��:�����iu�MY�Hah�����-7ĵ\(�E�2���fe��N���b���֧�C�饈Bö98i9�����q:DP�2��F�~����2Ģ�nCN)��~�8x�k���~!��b�N�&���*1T8������q�@�i1�Ѹ��|v��d2��a�E�tY�
9�L�Z��p�.�%��-ð���(����`@�J1�X�g���@n�G�B�q������Ag�a�y�PH���\9b��صw�%����q;���K�ܾ9�<Q��=���E-³RU��f=j�?P�J���7�]�?�=>��_��������l�����zxc((�AY��ܘ�쁪�{��� �B��m��L���H���n��.!\qU��p���S�g�!7v���/6�jՐ�(|>�/`����|��1�n����4�*n$�֔���!y(�C/��+JB/�ՙ�>O߻��?w��]l�G�\��A�ϳ�KLǥ��<�	�[N��c���a!�ƙ3��Gނ+|�ói9�O�����{��& b��yP: 󮉍6j ���;������=�U�e���\-�����-����/�����u8��^��	(8�G\Ŏ�o>��3��K�Ke����\i����/�1�y/��<ޚFCG�h�:�:8Y{�=�:����ó�V=|(�t�xr�\��r�{"҆t<�,3�p~��_j'�ҿ�v���MW���l�3�)���,��r{.S溹�U�meF���d �7���l�0��|k�+[���Ї�|&������qoi���ߪ��IQ�����F�о���*�
=c���s��*-��n�8w��m��'?�Ӄ%̑�4^y�'񶒾�����0�oDCp��0^4���|���4�����w��֖$
ZA�����M�����El�0|E����K:	h!.J�Q�	�M'2��q����th����d�l~uJKZq0�n޺��A�*wʙ��=�TM�����ͳ@�4@�F~�6P Nb�tGY���sx�G3��=l:Dtd�H`��CŒ�DS��G�r��� �OS��������{��lcZlq~�h�c�}����`�"����}?�IN���K��L/�b:�3���;�W�.��jMi����s+�����B�42�-�Odm����Qs0`��n���2̳��^�a�M��׉v��j�q�4Cq0҅�"jm��2?}l���@�Tqڳ%q�0Q ��R�[
��!���3I�!�J?���(�f�i'��ȭ�|MW��LhO�;ٯ��a���#6���Շ���{%|��pρ�Kp�!V����Np���,�T��㺵eD�x��dwSu�kx�H�dkƳ[;���w6��[����h{�ק�o��*dpu �۱���"����8�s��!�{����'���o���pv-�r1Gd��Go�3�4���v[�t�䶥Py�J��Pr'�A{�pďU^�X�q��%����5��2ƵZ6�K��u)`t�|�1L�%6t#�Ȕ����1(3�Pڼ&$A*���7ƍqd?�;��ƶs�%R���#���q_�s|�>�1h�%�[&�r�?YX>���P���e����⑎1ǖ*]��)-���ހL��m�C}f�"A[�9�P�O4rNzhm�_C�k٩"!���%}g!�d�j\N��WS��Ǽ��7���0N�!��e��=��P_{�B-
/��3�,��>K�3"Q���ޱь���,�^�U������4�t��e0�f1�%��̙%z�w6V�0��Ng7�����c�(C�a�p�L�b���`P{����ۮu�T�~X�s�zJ|u/(��"��gKQ����*����_�b������6Y[���8<ExQa���������~���Y0J��,�*.��"��] 49I��r���N�!�#	���y�Q.��p�³�E]yH:�qS��n`�G/���4W1ѵ�jU���¹sG��t2	]R�k����E���et�
�a�h'Ca۫bk�x�G3�3[����Jmf�F��~G�xm�X�lR��!���d��g��Nri;d�z]����;_� <�^#�
�PQ���#�:�/�%iWִp���\<tj�{�H�R�Ln(��"ͦ�5:�pt���l`9_�=��^��/�'���4�jV���a/���P䯘�3T��8n0b'G�[`�>"��8�a�i�8��(�<G���bC���
��{7��;��;_���^BGQyBH����� �v"������e���4�`l$q�Fg>�Gnׅn}I�E^cT��
�R���=�î-�M�F��FR�B�������t1��{[Wc������q#�}P��]R��6�̶1�~�̭Β�	�	�W��T{�M�Z�M���~����^�?��p0#YC�"8�e$�	e�>��ź�/*'0ܬ
��N
����`h�����c>�!�]e��!�Gg�$8���ڬR<���w|��Rԍ�(�R�XF�̂,�#�k��D�:/G�*�����]��u��_*�hd _�
�͔\��"8tO2����DQ�1�X8�;��ƽ�2��Drd���0�����;�L�?�����:�7�E/�ɘ2�RD������1�w{1�%��x�k��D������	o`'�@(�D{�h(�20��4�Ν�N�%%BV�aBV�M���Kw��+��r�xLXk�5�!B�����J�:&��M��*a�!��,��.��F7����
I�G��I���ЛX]��e�YE�M�/͘��v_��c��ouI�`(7�
RZ"�����Sm�ҧ̵��JK+q+�r3p�&2m�����Z�:��E+�QN�J���9���!�Y�<Hx�M"ީ_-ዥ#��M}��S����=m�qVXg�׈ē#�d"��O���9n��R��f�f�Q�D|�_d���N@�Rp��"uU-��;w>�(|�ӟ�����QO[�s�M���n��$�M6>�l�h�~/]o*�޿�Ɠ�yg�6�D���u���3h��~�Y�`h�,�`z5�I�U
�mH��t�'����;�ac7,R¹͠(��S��%����1�Uf�y�t\Ӆ�q���DdJ�F�Wf��7u]�7���H�Z��w��9�>���R���p��Í�P���-�l�w��m;
f�XiyҸ_ؒ��m�zͦ��i�ul�����*Eq������sI@.	�S�ݼ������ۺ0�"=���z���{�����o=s4Vl5 ��a��Q#6��$zS��Nh��?,��;>���ѡ���Qh�0��p�ۆ�^	�4�W]�dR�j�7��]{j�s�P�JfZ'��'m�r��7q�؁C 36NCB�i�B;5D��8W&�jd�r,��a$�J�(Y�f�/4^�Eh�/�����r.�c*Ё�	��n�\zH�ҍ2�GZ����U�랻�G���������Ǚqb��r>b�jLgR�ӆ�T��c����Љ�Q��m12�1vT:y�����{PN��u�ڑ^X)���˽`�{���ȗ�!:D�9t��^@��f�Ͻ�G<�j��=���Y��*�!��k޷��H�th�B:�yD��e���]����F�#�׾*�E#J4f��@n��M�J���䖬g#�1
��xcHj�o8�������0���X��"yw�<'�#�+�c�Se���\�(�Io~�I(f����U~�F|f��ܼ�M+��y��=p�^�����ְh
��x0�ȍb1X˾ץN{���'��U>��#<�L!�+tJ��lz�u��F��Kw����=0{ͫ����~�5M��l�zׯê�0B6_�7��RT��a�#��a�d���� 7���V���3���t�T��u�7�w�Mڲ�ʹe�LdM1.�z��=Z׸c��6N�˳����=!�mrnj�g��DЩ����������i�T�|~�F�O�b�Ox�xO����oH�R����b�z\{����n�Y�v������d�JƗ��B�E��+��=�L�qH�(c��PiA�jF��1��`h{9���U�ٔ6��x�f�DK�q�=[a+�BRR��s��1��8�J` ���8"���5�E�)yڞgΜ��({)���ۂ�>2�8�-�B}o��/� ݌9�����VI/U6�KL�=��:�G��6<Wl6���otT��$��:7�L���|���*]��=�rw9�Oh;��������(!��]���S�r>΅~s�AS�%�@>�X8��HJ
�mJN�h�;8ЃB�c|P��-�l�����^wV����8�Y��u�l��� �+��O(û
	�X�W}���Yg@z-H��z�8�*���OZ�\��n$ą����,���� ���˖̇���v�TJ�'�{�O�Q�9B�{�]X����!�ϝg�:�r�>;���oPN��P��x ��mgaVN�j���K��������ɽ�{Gơk��(�[]v9��2�筬i�G��BK�������y�'��rOL`��X �3��Qz4TG���uƱ�a�"� >����\���4��}�f�{�Ń�擟��H�r%3�0Dn?B��ϥ2f�U�w�����A-���mSaޠ0��T[_���r
 L/�$�o#&��M0n��~�ˡ���^xY�B��M������rM���]@�Dq��F@;��s�� )�_����>u]Tz��:!|��R�b�l�q����'o^o�3��8�nT�R�)�c��7�d~��d�ڏ1�"��P^#�{6�l]�F>�H0�7�����(����2X���S�>�$��I�n�W
��LO������R��B�[�һ�w$�*��6#�zM�$��e��Dn��]�@�0�g�,^Cb �C�d��C\�\޵����p��WE��I�?�ɒ�s��L8s��6Z�
�N?VJ�҇�!Mp��p��t���|G���|��{���u���������B'�M��|�X��<��A���x�$�xn�R��`@���N�p0�9���F�$�K�ձ�0ł�����v�~Vޜ,�4(���2���~b�R��%+��'c���*T�eTr�
6(�� �q�4r㉷�;V�`�`ZY� CCә��/C]���U�S=<r�����v�Q|�@��wd(�["qx|�?Q���x�V�sll��st����-���M��J˜�'.-iO����K��t�*w�����*�ٚ�gBW�jd�� ��bX�J����fX+��ú7�^�ڧ�f�jx�#��_�������7��\���!���o6}C��K�@Bڇ�/�Q�f.��R�5*���~���W��A�Ͱ�$;bR����Ӿf���3G@�
����?P���o��`�#��*vNO�5zՇ:� ���9���,����BF�y���q_�W��t�`��}���x��.GQ6��~C��!=�(�g��3�d"��J�H���[Y�dZ����������>�9����Y��!���ȑ��1tղQ뼑D(��+s��<���E�bH���x"/���=�굙��N4���#?i�S MI����_��BK���=��7ב���Uq+���	���xz���ZE�y�֦��!���<��:��+�������\���ߎM�Fߟ�9���؛�C�=x���K2� >�U��t�����bG��K���(?���L����Mo�2x������+'+h�{���� �זprҒ���["��!=��,N&1�{
#�y�*�>�e��{�T
��D�<�5-��#���Zmk��Nj�������L=�i�=f�`��K��i�7k�k&�>�X����!�5	���߹.$�O璷�;yi_�vI>�~�ۈ���3�;�)�i�n&�t�18��2���谵��0��4�<]/gԸ���9�K;�(�AB�m�'�F�j��dbL����Z���Q�Dg=(�/W��*�;^Ǽɧ��|l�8�$S��!��X}� �M{8j$5r��X�2�h�����0��79P�B� "�<N��ӯ8U[�e�Oj=�&�i(/a�x���d��qW>�WӒ#߬��n�<j��c�`<j��O|���N>�O���F����/	b�U�����rL��_vr"��]�3Qn��D_�{*�n~q?aXk�/`�*l�G<����VN4P�؂��|�0I�I����C>�@'�`�`�$�/	����ɸ�Kad2ć(@ӥ^�S�����`g���3]fKS����� �\J�'�wٹ��Z2#oNS"ݏtN�c�Ձ�J~��JM�}�~≟7aA��Oz~�纺E�p�
�+�C��̾�R���ˌFrc(���ɯ�/ |j�mU�o��
X6�HD=��<���K������	�+�XN�T���|��-=���Dn�XY@����f|�d��9�9?K[����l��R)�U�cq��d���̞�����X�����~/�R������R.���k�PNjx�tX�\5<�q�����s�ʔ}����E��D�G�������8_�m9	ܡ���n�/ �Q^���"t<�#˹��О��I��ո��R��8��G����}r�����tz� ���4�l�%�����p�,�!��z'"�ʁ�ICF�s�2Ջ�JN����q7�
�V� ���'�34!��J>�*yͻ��{D��~;�H%�H���F��D1}W#̓����ߋmng�&�|�n���:�1�J<8Kuh|~g��7;�n/�/�c��v�i]�	�ç�ɧdT+�r��#�%|�{��8c[��[Ӳ�t����hD,��/+D�fqd`�GT&��6�?9 vqr����%���)�>'���4�Jd��u��g�T�⟝����C����R}T��;�Qu0$9�b�S�- v��d�@�^�k�6��t0����.����l�V�Li(_,���o���+1�~³�U��W[3�4'���*'ܜ���igևs����yp��M�5$�i�����lY���8:Y~d�-O�� (5������2�28��W�	N6M���XCt��óL d[���MQfͳ7�Ʋ�-'�M�./���^�$ʗ�N���B�0�}��#�uNM�� {�s{/@�B>1-�Mgh
6?AaJI�Bl���
�aO
A�g��wl�{zO��P�
��
iH�n����p�߸9�zx���������������pp����l��#R�!�cc~H��:���<gR�ևgׯ]���������|N6~/�ɕkW�W~�cppx�/�1�UԼ7+�m{�Z��{��9��1�xL���<o6h�_�����aSV+�P�a=����3W����>Kw ���?0�#d��hu������U�pW�1�GZU��9%>l4DZlj@7;<Ȩ��]��`�:��C���܎��L�LĎ��H�U\'*Q<�\Z�~è�w\�i����"�/�I��n�Ύl�6cHe�Ny30�o�7m*����ع�`�����p�͜n|�N�}�������W����ȇ`ѯK�9L|�Ƞ_����r*�rc�(��3J<q�q�{�s�*v�Ӧ���/pX���)�n��~l�6��������о��v�ڞ���5���M�'kXn�{@���_��T_�3����#_����6&�:������}�뽭�>��-�C����I8���T}����8YG�^��)��W�&���c��ﶶ��e	�h��9�9����.'��C��MK��^7Ý=�Rs"ʄϳ9̎QL��4�LX�H�D�@����y��H|Fn�-�\xXB��7]E��ʆ'��wt,�];`��
$ʖ���l��G��+���:r�������2^>�w9:`N��|�-܄v��j7�;O�:�����b2/�#��BQ>c�|����o���+�O�?�j�)���s�Gp}}�3�z���g�:�b��*�2�f��弯�hM����tn��%���� 3O9�4lB��G�5l���=K/��J祚�䱌z��=<seG}�F�z½U��rT� m�+|T�؞A�{� �*���VE:����Vm�>�ӧ3p�����CN�p"P�;F� 8�yB+��`YH���9�V;�tO�/��8N��@�8��]9�`cq�t�۩���UY*�
��q�ӗ�0�cVm��o���!�p/��?���a��z��u�Y/9Ϊ��`Q+�D�ً]#s|ơ�s?��t��~Ž�){�Q�=���;{Y�d�p�b��y���QGڧU`�iH2WZ�a��K���͛��FkG���,2�M�K��&峗ZI�c��ģa<���`�F�4�uF֣t��ρ�����T��.��X�7�c��{��5��|q�]�8d�f�9Q��p敞n?��8���ľ�BlH���)�����l���]g3c{�eu�1�Ҧ��/�1������<h}������|��tYb�ѷ�ޖ�];�"�[:+2�i�9F�ہ������+r���7��R&9�X9��W����Ş�;�7������^7 ��dTv)u>�ȡB�+�9G��T�~�s�~����vY��c���S�3��}�C%Xl#��K��2d��hFZ��1�����A���L}��V�y���ٲ���o8��5��S�R��m0rn|��a��Gpq�4:ֱ~���$0�����=aq1TB����]��`F��]���/�^����	ky7�\�3O����?	¬�N׉G�m�&�s��9RK"���������^8��N8�?�{�������4>�JHD��AV�(�������ϺhH���}*s��Ѥ��S�4Y��|�v�����G�gM+|��7�������If$d��A�������9����?��5,�ЮZh:�)���_0�x:�y�a�I��4��묆s|�r�V��!{��1��n�[����aԥ�k/�[��Cw��`��=Y*R=�����ս�
�!�����HJd �g���O֔�a1�`6���ݞ��p9�'�����_����/���
u��r���4t�4|�+s��N�&D�F���X�C� ��|�������߃����Q3��
�o��o�?�A��_�%<�j��Cń���v<��{��K!����0��'h� W��j���p����3�?���34��0��Z�x�:T�Wh�x��y�[�4.�w=���@F�:R/t�ƫtN3>�9�i���������vW�k�v�\BN��Ip�/��x��-ҟ�O��7*<���@V�N�)�f%*$�q؝�@�������5�9�Ts��f<�a����Ĵj�C1��"Zѡ��a�(1VB��̯V+�,`�=n��	\�/��o��~O����ρ;�]Ҫ�x�q�<1�Qc����9�3[yϖqZ�R��c*� �)r�^.P���˅�/���<�5׾�]]��h��@�]7k��q��֛�z�1��.S4��/�_&�(#�_7�=��ʉ�4����0��>]���s��m3�~�\D��:�=Ɩ��%�C|n��Pv6�g�F����a��܈��ԉ����=2�7m30��Oɸ��Hj�S�! ˾�FE2f"Ǚ�xЅ��s�dX&�2]C{�[.Ea�e���7����Fu��������sP�u���,��/���Y�z��Y'\��k����A�A
��w�r�1rx���QG���K�]�-::$��{�+��U^35}��^ƱG##I�v��Kd�^F||��'��N��h���d5#�qq�]�ޘ�Q�M�'k�_�&�i��98����ec����H!�4O�4�}6���C?�p^�����*Q��Q��'�ӝA�����'���0�rR���L���ʒ'��`B���0h?O��u�RG�y�U�[��.�E-�A~��!L�੷���W.��E�AW��Ԏ�cG�{XP	��s��xw��CG���C��D61�=�?�D�ɲ�iD[�iGȐ-A\�������Gd(�T�4ľ�BlR����q�����σ�r�䤗�[�CX?�n��y�3]����i���<��{�-S��͓�iTΟ��6r�X�'�wG�lx�K���e����d�R��y;�u�e�\Z�1v �R/SƘ��)��\.� #���4�St�1�1�;�/{����>zI	�����O��v�"�X��C`N��q3�����1=�4ޱ=�p0��mMű�o��8?e�y?��h=��+N�e6�ћҳ�N�FQm�s�_8����}��}NQ�}���7��/�Q���ol�7Uv���8��/����I5,i�"'[��`	�B{����z�/�.C�
}\~	����a3h�]g�4���6D`kJ�{�#Xٶm�1�q�� mV��m�F�kJ��+��έ�!e~%xh�e�0�cmo+%��O;�ƽ��������.acW���P����(ϭ��m��F>����^B�6��i��$lHoüO����C@�q27l����A�)4��F��c����a/��Z8g�E�áڃ�y߸�[}�׫<=��mG���P�f��ɺ�����y��o����p����������B�:�i(�S�¿�� �/t�M�6³����9��7�@X棷��Q�$h�x��--F�a��L�L�nO�mJ����G��N���+<�<ޝ�.��"w�Ѱ��B���	��V��[h����E��� :\82rX�f�7��hW&�Q��s������y�_b�Θ@�a�"�Y�[�=衣��������y9ܵF��&5WRRy��Cl�p����y<�#"+z2r�sPHGt�	8*�3s{����k �^}�"|���o�g�����?~�66�l�� 'r���'�8NrQ���I��Q���Ưѱ������SO=�O���n��O��؏�5����pt��zVs�nм�ֳ�"N(�@YQMI�  ��IDAT7�iZ�!���Z������x�O~��?�A���5���Z3��v7�+X���o�0tзw�7�zZ�����Վ���D8�ι�8�Is���郤�`:�SQZI7Y�~p��dU���`w�B�
���O���qx���?��߂��..\Oz�b1CDw|g���-c���Lzu$�+�{I�L���9�S�plp�Tא���T*T>�	�>dwI6J�y�� M��F�J�7���'Q��3���@�Fo�N����J���&8��+�p����1��G�)�T+��.�(�H��ÿJR�ɐjHg_�(��*�2�D~4Դ.8ЭB��1��?���m��!2�.�U|׻����-pܿ��X�iuE�񻦃k=^���c�m-؃����R�(R��[�IAPz!���K��O�s��(%���ѿnFw�m���B��$\\��p�Jt�zt:�[ӓ�G�#^�oe��;��v���c��O���{�z/�Ö|���a&��a$�.�������wC���_�3�#��(�!UJ��\���|�7�z�L�+/����_���-o���;a5Ng{����]�:Mdl�e�S�Q�x�Q �1�i��t�����������ɤ�H�W|3[���<�D��[#ME��d���7=�,C��x *i^d���(�@�8���$ℏzE� C8�鞇�������_����{~����(4�&�]Ǒ+3;#+��ؤ|����d�+��p��f��;*��Pե�z�:L�z���vgW�O�~���\���K���������|���CI�ϴB��YyQ���=v0
{Jdr֙BE��$���b6�UO�������W��a�RG�S<�gj��A�@�j��҉���Y���(�:�}��B���5N2��u�
1A��>08f��@#
Y�=Ȗ�X�f[<�uQ��� &�4QC$�7;rՒ:�ӭ�Pe3���f�z���|fW�B��߅����?�����~GG��z����k�e�
+�(B��t���4����Ǚ�ٳ��k�';q�Ni�\�Q�X�#��]�w���`�4}N9���)�=�f��$
�G��*���)7#�Oų��y;��B��YT_�t�\U��Sp�K	?�zG�NRw�N涐PJ:Cn)��l��3��;��]�<�E�Q��cEz�)6� ��.\�ŧ!Rw��$,�سF`�o��=4���
{;p p,T�!܆��L���\�� ���0:7�	�ٌn8�p�M0B[	д�����`3����!��7��U�l��Yy�!�iϴ00F��-�t~i���C�ǋ��ߩ�7�; {3q�hE�,?��;-C�m�����]e� ~�2뛅ǰ]Y��W��B�+0�K���/[����wC�t���:�3�AcKk䔺I�d��G7a9��A����x6�0���r�O�\�g)��\?�İ"Nh��f�aB[���殻யx������}V�^�+�3x:8l��в���Z4>b^����Q����"YG�xn�
7K1r(�k"k}q��'��e�ފ��p�Q历Z��-sc\C"���� ��2	�I�wr�YiG:b4�J�LϷ���{F��n�U�]�>-1�XS����E=��f0tI��j�����w	����|aX�Si6���z���s�靈���>r���Pg��"j��>�ԨA1#Z�E�(~�g���4{��8�d�(�uS����,8$����Uh��C�����|�#?��L���d��j�`U�ъ�䛴:�ct�0��ﯥ�)!�����O��~�Cp��9���U89���V%�*N�"�.:����s�6�:�Ox�m�4� R�4lV�/���o����}���.����a��u�b�u��f���Hψ6����΍�'_�64u]�nHz�ny�CqF�h�����Dp�9��� Bݙ���98|�1x�C�����xӯ}~���c���}\s�z�]մG�p�Z�4/P��JqIo2:6�Z�h���.�=�eŕ�T��>Y�-d�$�mD�Bƅ�E�vu��.O���K"�p��P'���A͋2v?Ǔ��?랟�����145\��p�;�	7>�yx��O�AR��8U�)����psTR��X}��v7PJ�,���\�0�Fk����ס���z^��Ae]��D�~��7���z����cX�M�K��M�G��vc	�zx4>:4I��4���T:��e�Ω�X/��^�K�э��m�Yj?C�>�[Uvuk��ۃ%}��âkD=�c���@�kҎ��i�Q6Ǜ��)�\o�/�P��(���]���S3J��w�7����}��^ls>ʓ(�О�t�lz*t��{���Ư}7��m���E�L�{��j�����%�@�P:�;N ���zh�t��Ur/Iq�zH�60�>:.D�n����0�4o�\��*�F�!z��2>�G{�K^�H�P9 o��/�ꄂ�n��bG�t�Rʵ k��6EjN�D�`����@2���ގ��K���!\�3��L-"78��,��yk�
1���kG�&OC���}���G�>Q@�3�P#2lR��`x/�7&��t9�t*���ؒv��JU" ��$"�Acq~��h�>���tv�1�T;t8�xAe���c��u��Q�nP�16c�G���B��#�����cK���)�`Xe ��ƴ���u�
�bv��@��D�����b?�O��=@Va	̫�`}�8s���ǿ
^�[�_����|y�׭C�����}�@��V �@m���j�l#�R}���lq��l����;"S'�Q��c3&���S���ȥ��/�v���f�]�$v�_J�SK.�Eۡ7�uXn���ir����k�zS���^*)������x�⥌��3�)�A%=�t^;F_�����L�4������3���H;��7�{]c�X@=?��|�Ӏ��� �n"�d�ӗ�~�p�w����8H�q� �Q9���kU�s.C^Gb�g2.i�$��v��ς�y��5�a:�@��)z�
(*��J�n��Ύ�1��{���	Qҍ��3~�y�J6�|��O�Ǔ#�.2�c�W^���<o��]��f�C�ȷݜ��������ݶ��{�[����b̭,��0��:��+�7wBa���7<S���FJɹĪ]Zo�V�>ǆ���v�c��1�����[�Ny����gKgs�&���J�ۧ�
4�#����A;J繾�cj��Ϸ��_�?PJ��1P�yN���v��
6�z-w�\�sP�[౿����G���hf5�L�NV �J�C���ۯ:��E�[[d��@Ó�^�8�"��wIF�|a~�\��=��Eg*��F����j�7�J!]�aqc�ؘ~��*�k!��9��ԜB�1��bD����_G��������Ͼ��܊ҙ��p�m'�2f4��`@.�{[8�X��'��3~�M���'E*���u$	J�
g���!�,����-��S�T�)�߬¨��
�{��o�7��0�������3O�a/���������^Q	^�!�J��
��t.���:2��>�=������$z�=�q7B8�y���k<�����UxkUn���O�;�HGy�%Z�pH\�jC�fM���.������'��_��uk�q���Fh6����iIBDQ��G�1H(������BgyW�J$������_�qE�[���#$x��d�����&�+��/���z���}-,�ſ�_���g���'�	qD0�C����3tD������8\	{ӹK��}�{pBxUTo�����-[:s��z녷�{�T�pDcb�&Gt�<q.�r���0G�<vCy �蓤b1f"Ḽ�Pږe�^ê���� ����	�ZW�=8�Ż����?�����������kt{���(0!�L��	'�9���oe�i!�u�%�*�8UP�����&/���!���s!
צ����3����y6�4�chVKLgn�����rW�a�It�'�D��1w�P��d�8�d�A���NU��F�U���i8%��>�V��bd������z�]F�k�pSe�n�zVi������wK�W��� /��w�Ȍ��AX!�#˖����ó�~�ӹ^�j��[�o�I:���>�b�Sdh����;���/�O�"+�2_���c13c�<�=o���ǰ�p'�x�k���~����M���|��其��d t�L�F�l�X&�^2M+�
�=������e9���6
*�	�6��ֱ�Ju��V�_��2�gtw��^��wy�b���Sᑴ�V8� ���[���F9��8s��Y:�m�G�Z�R0xg�� �^��Q��,`�Ru`��F4I�u�WY�s�D�Y������y�H6�'OJn/��4��bٙeՓE��i%�9�F�h­q�N��ϨF{^@W�s�d�pmA|����Φ${$�g�
%�O]�m�6M�,�2!�3�f^�tG�^�� ���$�eV���|���ƪ���;~}t�_����S��'>	���_�����p���¹Ep�ZC�Z@���J�� �5%��_:��z���,�&�3sh�p���}��H,F�E�dO�ӑ��+o��o;4�l���sTnSPǋ��n.��H��G����{Vο��/F)����<"��Sz�,��.���Yr��r�(�R�;c0��7���8oW)��t�m�/�^~��k۰e�Y�b៏�����U���=Wҕ��j���ңށ�)�&?����{���]�I�H '�Y�s�^���p={��Q�)�M�RN�BEF���()��$�����г\F��soT��-�p��I����x���%�ɖr�o��{Q��yK/g$�P��q����ĩ�k�b`���r�RD0����R����Yg��?���2�ދQ��Y��U�G�!���9fȖЧ�`������Q��'�����O���^ޞS���\aSH�[Q4:5�D���bc����WEH����&�4�:oH��X�P�|���{���[�/����պ�E'�L��v�Q:ȁ#Dڈ��<9�H�H9��H�V�U`!P9h�R,���.�7k[B`�CF�����s �o=��Ԓd5@9�CjD!���IÓ��؄����>��+:uػ��(�c�6��`�.���������-c�ʸv�^*S7�K��/t�ձFx�aT�	u���jH�5.G�/��m36J�{�	S
�^��Us�����jSç��W|�7����.���������/ f�amC
�@���FCc����+���x�)'�t���Q~j�R��"��+�k��P��
fͩk��&К�f��[�����o��W�W�w���;������ޱ^�1@p����&[�_����v^����60���� �B8�r�.a�50{�i��tj�i@�8�	Q5`�\�I{��p���	�x��p��?�����ys����E7a>�s(A�l��C7j��ޚ�)����Ý�M�
�>|8����JBW��7�d� ���qX�cI_	'�
a_��7�W���a�������o�8s�x����]G獮>���;r�D=1����U�g2�8��\�QH�ө�:o����@玦���?�MK�+�ǿ��G� 7�y����	76���������2D��iu���c�-lK��6�Qh�|�.�O�ioU�����SJ:�M���Q�����v�ld>�RVKf�����J�gm�ŶClS�+��;�=gl6�v{���.��5�o�{ɸ�tQ�J�7�o���7�-�K�,ȝ6��87gT�sn)BF�j��{�G�|�M���#p�Mo��!��@�n������U�,@�wt{�F�L	��K䅩"c�(|��;�=�0CM��S9R�nXvb���M�s�$�>�ͧ�^���e�a�ZKi�����wVe ��^�PA)�%QJW<ґ������u�o�^u�߫B�]+$�/|#�ʹ�|
0��w�"��`a�ُSf0���8ڐ�d% �%�Q��Mڒn2�_�:���_r��K-�zG��]�@�h;r>�|aƗ���M�����q��T�:�O�w�'��K+���NB�)o{����
�4ϒ�3�~��0��RegȘHq�	��xM�9�^���o���䡇��-�c��]���_�������4�봞�{]r������@O+s�H��x�	�v��8��u�M�	�����*8aH9�s�N۳�1�unS-��m���N�¡b[�c�ʶ�l;���!�K�0��K�LՋr�zR��^�3�~��̶:S�y�~�۵��̭�y� [�0v=�b���/�I���Aɻ����%Q?��Ob��D!�Ԋ4�K�c����/ܭ*1^�d�N�-�T4e�Č��00����X%I}�`�(�T|�Z�Ո���>er�J�2��s`�)zVhI��<߁�Q�n�]�/.���eN��f�Џ��B+�����Q\��=m֠ ���K��\|c[V�W,Ev�~���Jo�7���]q�7�O�qg����Y�����h�#������7�m��X}��Y��1ǎQ�c�L�}�o�im�za)�v������Q�(-w��B�c�8&���]��:�n�n���[��?�!$�jm��R
�[���p0n��.%�cZ��8r��ޤ������툡$���ɰL_�44��Y-�CG��3�~�-�r��\�]r�dd��`�S��ȹ$}D��8���$':��[6� �5�A�A��_��7��,v�/��Ff2�)�4���v�>���z��;{o�V�u�,�<��G��(���g��L�4wm����|��g=	�(yH2���_���>�Vx��;�?����?��C��Sp�0�6	u�ЄC�p���hV���(��bG.
5
:p��7���n���o~�`���Ixq:��N�o!��_m�m<ޤ������-������^� \�^���6e�iR���)�3GKtQ2��������T\f�+�S�I�zM�	��y�:T��M?E�6Ƒ ۶"�A�V���7\;8��>�����o�����8wtZ	���y����'���y´�sK�<�>7]��������T�Y���;Jπ�dT�C�����C>ו'��1Mp��%�f��)����ѷr�,����/�����<�[���eh�j�����H�E)��"��|�X�L������l�'��ͅ�]'{�?�dEK`����F��G�y�}�Woz�y��=��v�{�m�����׎O�ڍe��:
 �JD�S�f�J�e!�b�3n�%OpV�A�xd5.w�>�}�ƌ5;�It���[�sX�F�*�/H����Pi[I�������H���f�i�kE��؛n�.�JTAYq�^��;|RCd��㴺vi����\�O���s�2��;���-ȆZ�y�f!�j$�y �L��t��������~�@s�\i��o�:�!��v�~�����!AO�V���CA�D0%���9�窲W,�4:��Q�7y��Ƽ�tO)�t�\L���'aw��J�7/�M�6�O���e]2M��1�j0�D�3O'1t��-ś	�[B�=�DIHi��$�	#�m!���Jb��X�ʒ�+�;ȫD&����M��\6�&��	E(M�c���A���U���qvQDH�=(69�T~#��7�V��Ws긽��tF������b�b��n;.�"{+�<��[�/�_wR�9I�j�-d��zt5ٞ�qYp��p��uh�\��������?��w�.����^��c������7Oᘀ�*\�)�],��<�th|3��c6�)m���r;������>���K�L��u6���Xݱ�/F)�a�\O;�)�J�6��F(��1�}��F��9�Q���|�e���$��βn�l�}J����}� �ʁ#��,�
��nE��]a����=���xD]�{��mZ��0�YK��}�o�wfhZ�M!�y<P�1�5�1��~���n�t�^G��3$+ic������ʒ�W�LU^��G�c�o/�@��[1*F_�z��>��E*�5�mX8���P?�Kt���v&,�<�PTT��=7�a����c�]�@�X_n��;����)e��IHɵ��^u�x���m?��9׋7�aZ����Yo0�A���;�=l(�P��"���Eo��΃�YF>G4r�B��RG��\�ƨ�x�?A��N���~��XKQ�_����%
$>ּ8px�D]�<�I䃁����Ɲh��-�����l��?��I'S�:�ɊRTI��e��Rȱ|�t�w����Nm��SL�@�!��P�-yK��z%��<V�u�o��h��������������~ӷ�/��߇'?�3��|����#����}��cY��vd�N����sE��n_�-AА�FzDoײY��6�ph+Mñ� <�Ӭ��%8��������G�k�%\�l`�n`u�Bc�q���[t�������'$Fe]v����j�7�e��Xq�k�Dmz��V�J�ׯ�G�ԔN�_C7���n`�~���yx��<�x�>w�0��1E]�h��X]P@�^����&�bUf����!�d�̠�~���MP��x��T�R�ɢ����E�T��㔵�34q����8{px �������N�׳3p�W��� ��߇O��G��o�6��r������k�:4{ZP������	�#s8q����*�s��9�cgOZ���'U�K�ټ���zx��4�ϟ��~�]_��qzX�V08�?;9>��7������i�Z�CҚ�T���_{H�u�M��9\ +�GX��e����إ(��3��Sł,Q��%P$oB���	!�w�l$�DBU2�Վھ�����Ȗ���|���9���p�h>�O�q�����q.���b��\����NrB����<<���	_�.w�]��cO�7�n"m�Q(�8N���<�\.@)�Ð{���5�f�o9�B\\I����G�%8L�џc�C�:��s�Q��:��o�V��񛔎��n�^�i�z�Z9��$����Md4�(D���Biћ������"|ۧ��Ʊ>H_]z�)������m��v�Լ�a��a�N�pj����9_*M+Va=�W�Ӿ�H��}��eB�9ϰ2W��� �@J�@r �D����"N)iO�K�n]A�����ťt��fN���G�fg觥U��."4l�W��9��7A�l�5�38��	i/�\z�1x�_�?��~�S�����P-*��(��s�x���aN?�DL�p��"��<Ɇ�����)�`>%�@�2tF��}�VJv�)�ߪ��/uGR'��O��.Yb�{�l�S����◗�ڌ�-9��:�j�����mc�c��X^�DF`9B۔J;�=����`w�{;p8�������f*!��e��8�� 7~@�莕S�AR�n8��NL��O�θo�	a�:���QA����
\CPw|%�)+4��{"���3
)������1���J��sT���FXIw�J�#TjA�L�*ăx�v4��i)W&�q^���6G�xm��/�J8�P��;�'�����B���Rn �Z%�e���TKY73�\6��%��p��86�VJp{�0.�;k��{j7'���`���e�RH2��h��� �Ms��&ًUa4�jL������E�"-�/��2H�	���p�r�:���Vp+xk�E:��lr7H�F�iF	��tV����zHAp�n��/�o����޻5[�\�A��Z{�#��H�-[�oR,�1�-�+	�N9<�!�y�
ި�*~���*��
SNQ@�P����I��8�eˑ�|��.{�5�ٗ�c���s��k�����9���Zkξ���{w���������;� ��]Op�m���}4h�s���dp[�h\��v�'s�z7���.ߝ��&\)Y�����s"�0��c�k�u-���Ѱ'�4�y� 92��cq�`�!6%
��A��<�Vew��c�b+3���-#+���k�?��2,�1���Ar�и1k(u �L?��ш�Z�À-���C%���RQx*T~�Y�>���Z�r y�j!'Nt��'�}v����S��p�������������������g����݇x�[�4��]��P�3p�����m��YpFD���BN%��aP��91�-�T�c�Oz}7�𴇧7O��7^�w~����ֿ��ٟ�����w�w�4 w���v����H�����U�t�x�RZ�Qi�7^R?�Z��-��^��-	 ш^��=�C��I�7.��=�w�w~�Z��wp0O���-��������Ë����@]��P�q��vW}8���骵�HE<�dó�LO$H&�tWo9w�3*w�.�0�=��n����8���I\��)��%6�ީ�'�-y�Ql�	JGv?�~7��\�C��kO��C���8}� /�2���|>�}�������8>�n���;]�Ɲ~a={���'�v�yЇ���&�8�`��7�����m��3���	��]��� ��0<ہc�/�rOބ�?���C?���� /���8�5�$
a�����|��� S�$t�A&���%�4�]�i�W�m��y�|g�}xd�i@!����3�j,�kH#��K��ԙ� :�iQ�N�l|BƔ��Cת�b�T?7�OW���pX�;>���"w�<s,��&����y�~�Z.����G�9\�5��t�A�qNؐb�[q��[�],`2*;֢l�H����]Nu�%~x�Û�'�����>>��@�b�#��ۜ=F�]،o�6E�,R���u�{w�+%!��Z��<4����`�+'�_��������ҫ�,���z�0O�Pm��NF���p!��-r��+�LE�?ȅt����m���a'҄@�(�;��{�h����p�[8�$�!_�{z��ŋ�=�iNU�V0u�[�c�|_Kgؗ�w��x�/dA��������;���$�N�6Xԏm6�� �`�t2L��Va��D+�>ڳ�
Y��N��m]6�g"m�(���J2~,�F9��y��ہ�k�����	"�a���,���W?q�{^�t����w'�˿?��m߹=���_��w�-�{�� o��7|;=�dOwb��uO��$>V�d�n-�?R�H7S+,Ql�0��_��`
�;v�s�f�lfY���1��?��o�J���"He	\,8��\��� �M��_'��hk�1Ѵ���J9s@��ok�����F`�	I���p{'7,�7�>oʋrg�c��0�G�
u����|���l��AB����6���VA�����N�m7T �n9��u S��/*��:	W�\�cR�����jx_�C��Y��76_��9�Fǃ�4F�A��iF�V���>A�
%��10�->1dè0�\p��p<B��Q�)i��`JoG2���5�Rf̃0K]}�����޳{�������'��;we�1:LO���qD�0����?�Q���$2P�,��葱�<) *+Z4�{$*�&�2�����%���|��7DCq$A��D�ٜ�Jc4"��.����Q��,�D�,���{Q��y]|N#2P�L����6�"�M�4�\R��6�'�;�������+p
ut.(ș&����'s��w;x���w��5��/~����W����+�����a��?����nC���`���dNެ��v�[�v����.\������s:���3�9���퉻S������.���� ��ހo�n������˿�����v�n�g'���m{��c�m��t�2x�z��3n[&Oq���|M�=`kǊݰ,MxGA�Y"�����-N��vH\��Ӣbi�倹�<��'߅���_����߂����U;ww On�i'a�#9�)pd؄����rZgh��\B�)�^eL;D�|����[u���+�BϣQw��C��ҭ���ln���»_�x����o��o��~�C������bH{�>�Ø��{Ì�����#S`䞸0���ލڻ{����C詃�AF���?}o�����W��/�8��'Gw��.}��~䆻�����g����] �����0D���,P�򙄲<ud ��K�=�C������ )�\k5݉��K=��˫-zИ����,�-�g�����#F��%cEo��E���
�sr?n`�9���ih������p:�X��N�2{��/�U�?����)�hᯃ���a>��x
�7�,e�8k�)fG�1�zH�T��R�RЁe<8� �u��E��ъ�Gʐt�d��@���C,2��^kQo��}L6I8'4���Kx�c���򙼬t5H�T��7����.���Υ�qB}EJ����#�ךp��,���`Ź��@�ibx��<�s1щ�
�Z�`P����t8/��>��D����Nd�O`��P�B\�̈́c��M�+?���>�6�/���b�d��|#P
��qm�u>��Gw�c��@����6��{~�+�����O������|��q���;޾��i�2�kd�	ǭ�ɬ�w�Q�;C'L�1wAqlslV-m��mMZ 2�E�8�rzh�wZ��,�"�T���>��K�<-vc�g'���Za��-p�r�d�t��:s������\�
]�ˮP��F��8�M��j����>���<|�$�#�s������T�c!�X�Q=�֊��7��#Ӯ�3������d\�NpY ���M�zbK
��p܁�rY��	���f�+�k�Z��А�6����+�&7W���>�K�AM���������VL��ۢ�&�V/�<���Z[Q@�h�#����Z�+�H3cَ�fƷ�#��g:*�=�8���p�ӳ�w������n/����!��n�c��T��)���0#ۆ���eBKSR��mx�Xa8E+�1 �/-��f�q��h�}�l�d;��s�j���d�&�I(�~.�͂��B�Z	� �Ch��#~Ӽg���1�W�O�  �%&� w[��a��-;Y������n���߭���p:xa����[������_����g��;�����
~�����=?�����qw��A��;��s$�Op;�Gk,����Wv�)i#k��{wb��*��;h7��|��G��/|���~~�~�w}7|�鋡����=�C��Κ�?}��O�8�S7�4����t���<\�]��8�s�5�w�M�1 �qt��r��QaL���a�[��p��`���f�!է��/�?�;�
�_�{`����8�S8}%�.�Z�QO!�۳�N�
'��s��ƵzS<JA7��t�FK���/��BpԐ����ނ��>hҀ�����������g>����o���߁?����������g����ϳ�+n�w���?����q9�^@=��~
A'�I4F�vC�<~�������0|��?������?tǽ��)]w�@/���_U���ܽxw�C�<P�#��F}�:m�#\�á�c�p����C�0��.)����M,hF��-��L[-C�!I�RN;�hJU�˞QOg�O�`HW������Yy�h:Mb�,�Q}��Z���>�)b��h���>�|��~�ux��)ĩ�B:mJ�8�)�����m��yl6�ț���eƓD,ϻ@���B�!cOh��2��O�&C�)�h�;�$+�"��+i����<���#2�;u����"���z��9|��S��D���?;�4�����IO�g
\�l�2��b��<�m�s�BvE�<E.��S�����:��Ni�'N^J�]���5)rIn��6e6
���v������)%F���t&�<��i2�p]�O^;·�s�o���~�7�v�IO��'���RIFnj�w��R����ʑ�'ͩ�ۼ�4�W��t��^�d��PV�O�yM9���88�������^�ĵ�s��m��K�{��Z�+olM͇�V��A����nm�>9��d�\����m����K;[��0��A�ރ�1=�����vM�;�$�-BPz��e��ה$�@&��3dI��EI�t��A��Z��D��.���s��%q�f�z�MXn��3����A�1G1*T6}�ؘe�x%�94��)$��������E	���q�z�b���P��@h�ҹk;�Db�����t��ES��W�E tD�7���Tz8����S_�QxϽvqw�ߵnO̠��
�FVϔ����e��4���\���ł ��@j��$i��`��~|f��T^*Ʀy���H�h�U������"q^�iY:P5��c�ٸխ9k��o0K���!�R�@�^�M';Ǵ)���&�-(������_Շ+��o���������7}��韃����|�������w᛿������s���$8�O��k��JZ}�N��ñ���n'�����x{w}��̧���#���G�����G�O�x�����;x��Ο��N����"[[��p�Ǿ���f}����/%�2�xt�hƺH�p��OwH�L��=p��]_<?��7o��#�w��u�����O�o�N�n��0�Yܿ� 
�!��BېS�QK�ݬ�\�|h4���F�S�XQR��2��������`���'���;�}�	V���}x<�ü�}���O}>�
����'��������?����1\��O��9ޅk	l���7�:2�Os�ע��_�k���"|�'�
�O}؛����������>.� 8k�p8�ӧχ��*���O��bߙ��9c<���ӎ��O}n��]������#� \�ibz���lϞ{]`6-�H���!����H�SfC�aD��D�ܯ��u:��ĎC���~�������޾8z9ĺ �x��?Q���Y�P���ٵx�$�8VL����-�w�L�6wخ>OP
x��D�Y�(�q�&����vGF@'-�GӘ�ҩ�d�׉r�����g�M�'ke!���)����1�v5ZgR�E�B�bY�	ԕ��/�,�{�oɄ��d�U%�WT%��C^Ii�3$3}��Z�E<N��:oMI[�<&^��ö�8h�s<����>�vv�A{|6�}�����}�������?�ݱ�����}G�(��K~��!��o�e��[�J�yj�2��19Y����F�_[{���5�5�ƛ�����X�\����v�놱�.���������b���:i:�|���6���e�,����Lӽ��P����a�%�*?}�`Ҝ��2I�"��g���^��&7�{�fr.q1��y��>���wS�ØDj�C��k�)������X�W�n����� q�|���T�Ns�"Rƍ���<H�h�7��2 '�*�^�P�Ā��y��8�'�X2^�w�[w�{{��_�y�p��;ww��}�p�ʔ��Mw�Gd����N�F��L���D;��R�l���������ˮ�!����Ւe�hwj]1�9}�8� ��ǹK�NV�b�����kFSڥqzr��z��E�mI�&�Χ�tD4�v�":+�;q�ޙ�P����R)�?���1�O90�w�c��38B���[s���9�><�w�=�g7���_�E���:t��x�w��������?�Cx��߄���P���w����	�N��}��{�����o~�cp���O~������~��������ٱ��߁��������,�g��c�2�9�]�������Х��N��C4�}\����䜮�A��I�~2���ﲡSܽ����}?���pgn�S_�
��>Ͽ�-�����-��F�F5�ӛ٫ݖ?����-��Xڒ��3��4$�/+�
Z� ,K����9�����&���=�~XU.��vo�v;��-ܝ���Ʈ?���;߿����^��>�%��>��{����C���|�o��?�����;1]�Ep�����1�ݩ�ϓ[��н�6���'���� �|�Sp�O�����U)���{���}�ֱ;Y'��uw8��g�B:w�M�Q '!��r�h���oƌ(%3�6��%�_6-��P{Y�f���f�����e-rI�T+�	��V��ۨI��a
3���;�����nL�wb�`���?w�����R.�N?4����E!�wb�*�0�r�I��-��t��`�|�j�v�g�DY0�����?�x��A�'%�Q�Im��!-�ڀu�z��4�x��hש��c4~�P�#�<��r�L/q[[W��ny���Vs�5@�K�eLk
q��"����Q����L���W�}�:}Z(�îvA����Ee ���6���'���ٚhC�7��ךl>�N�W�m��D;������?K���>=�}�����>��_�?���s���o��}8}�sA�x�$�'�J��!��#�����t�F�+�7���11��C\~�8���E����[�saNY��^x�f�ƥ]	un0S,�]���k�A�Ër-��(8tQ/1 �=����芙e:`RMS�e'pp!�0
�gI0`�a����!q�0f�Z�^�K�Ƿ��c�Ï:]<F�p퓤���-�{{dD�`b(��Wm�3'w+-S�
�N���#�F�HqI{ߋ�c�"3�������
�b�4ai��Ԍ+�?փ�v�+ݵ��176w|�Z�sb�<��: ۡH��m]c-h��i����<��4�}��7�G�]&��R��`P9m�ŵ�u��Ʊ�t;kbt�r#	G��i�e���r���[?��8Ϻh�s<�hN�Az�|�{�������ݝ�n��Ǡ�3��j�*L����Ɵ%�qg����T��0J�Ĥ���O �a��H~���c�`��8�٘;~y8_���H@��ߧ�����3L�O��<Z�)$�ꩿ^�#�kyW�c�)5��[�^8�tGn����S���U-h#�W�Fb�e���i=j�=pA;�a����~t��n���i�S����~�t�]p��»_�*��;���3�������~���7��|���� ǃ?��t�ܾ�7ނ�>�1x�㟀���Û?�#���>7��4߼���#<;�p�{
��8L<�=������ѷ�4<�t�;���Q6N�4�-����Is96#N*��nXc�[�����h�P�7\9˃3 i=�2~�3\�쯣�\?�na���k��.|�+_�?�/�kx��	���p{�3g�;)�����#�:�~��uz��r����+�b;�<>s��A�A�K} I� �	)��8�1��?�Ih}*��yk�0��w����T���	��sAϟ��0�yx��q���y޻@	�gC�o�C�>�dn?��"���/�w=��Ú����ٟ}^�������?���3w�����o���'o�o}n���|�]���������-���P�|�;u�M���ޝb㜟N��؋������������������O^C�Ųc�+dul��=�8���r9p==`=h�o�y8>����ti��v���.�5�+4��fB6NΪN�/ݷx�U:j���PY]V/}6��w���0�8��A�p��r���<򨯁�PЩ�=Oaޘp��nx5P�AV9������?/����ׯ�q����=a}�nl]���qEG�}E)e�.�j�F(-�7a���B�(PI�NM0�C�~><f�`zjk[�����N)���.'�K�̋\߷�d9��F�Z`/c*���Wӻ�E�st�5��w��Vkd#B����2�;}!_ol��Ж]\'V��r��]��v��>9I�*����� [@>?��YAI?,������La8ι�����3�_>��:jc�o</_��_�t$\�}� �s6:Ό6w���xpW��y}�f�3��ҏ��~�������_h��q��+q�db̙�B^7�Q֏t�*�8��ybyE���Q��[3�j�
QW��i�f��[�=6��1�&�9�>c�^�XHY@�|��i�����2N�xE��:<A8�NJ�� yj;�`vN>,{gLɸ,<����s���J�<BF�+ϋ_��N7X�D*�������c���s.�����뵆L�����F�k�X.���2���r�z�}�c�i�N�Q[���WJ�$��ʬE`�~��Q~M	�b̨Nm\J�X�8='Q�ݜIB0&�S�X ˌ)�"��$c�?.�d��P�'��0��.x�w��C8q#�	m������WЏ(��yP3�i���8e҇�ݓ���jȦ�lЏ�V����4d`:z����ܑ�ec� 5)W�-�ܰ�>mhQ^/��>�1��7��v�`�B���]X�6Zެ�wOɵ��NCy��{��)\a�&��78�ܕ�M�"��vxw�ć�|g����-����w��c�?�a��;���x���P��o���пv������P��ߝ�ِ��އ�;���$6ޑ|���p���'�T��:gp>��f���E16f}�t�a�v���g5gX���$�!2xƹ}�xl�����On�n�O�G�_�U:p��=`T9��t]K|0��u��	����E>j�wuE�����S�5��ǵ��t&>1 ;f�v�v���>��0��������s��-�]��hLd��`�������ͻ�?�Yx�N�����aX~�uq;����� ��	�5zt}1�����������ܕG?�Nn���G����p��a��h��(\ů��<���0�;�|��}�J�����X�Έ4<OX�/���N��;E�����������ֻ�VӇ��?��v�����ʓO���O�3'k�.A�Y���ʒsT��ԃb0� �ڔ�"�4�y;Mo�4z��O��'�����J�9�V���Iw	��e�I=��O�o]:��`�	V�q>o��N�щ�t�i��X��-�Jڽ�O�8!��r���m�	k"��q+q�J5�ӏ�K�R��n�~ʸ�֏�n\�.�c���X�:�yԅ�jcz�R�zL�����~��|��۰{a�9��?l:�8I�e$�g��d�L�]^WAD��-g��C���i>�ll�*�n�����,��r���E��r�@&(L#�#e��|�y;���\c��j����A�ѝY�,}�!�sAs�7���Zbl���u8�^�BN�j�A��w�..^�uU�`��jΙ5q��V޵�N��m�%4��p�m�6�/�_�'��}>����=��x�����ܽc��E�{֙�5E>��#�io�C�^(����ۆ&�GAk�ˢm�����<��Z����SC>������i�;d�P��L�Z�r���>�p�����/��X��6��C�v��Ooq���Q�'8���̽���J��ޝ��J�A��B�3�3��A���va�ہ����{cHc�c�;�K��;`p�GO����Cp@?sAf�p*����&����q
�q����Q-��M��3�(q^���v�a^W�T���*�&�8p��������a�4���n�7����# ���p��SX�����i�og��vR�s��0o��P�����i��e\����<��������ݰN�p�d7��ݠ����*nG��v���nXk�]8��9���5����ׇ����.�ats����O�q'tx~禇�S��?!��k�H�+��ux8|���p�[�HG���%�3�OK@��2����	FO�x�ۖC+j��.���Aև6f��A���){x�K_���?�DO�����J5���F�i�Vs���4�A�|^�
|��E]͈�teu�W�)J�%��%�婾�F�����P���y��T�R� ��!��Si��z�f|�J�aJ�z6W�A��-i��j�&\���Z�ky��?OF�d��:�u�(��M����4�9K����P�~�W���Iѧ�)Z��N3'`K�6�+J��*%��p�A&�q����o�������?{?���t���Cj>6�̞,�l����T��q�.��-�Ly�
�L��WQ��as��y�:?�����>glyT�������B�jh�Ы���Uq��	�� N�圅�q4��_��NshP�����GHsC���|0���rU\���m�KZ_V���ߺ�Ng��=9ߐ�V���w��� �	kq�	fbhRi�?=�f�}�8�#t��9a;�#F�*8�h�BQ��J��p͕y��cԺC~:�ҕ�qC~���ɔ_�R%s��I�o�a���_ԯܰU��|�廾����v.��橻@/�`�}��X���O�A��]���e�퍍}i证��)G�=�!|�Ӽ�u�љ��7*�q�9Nnד�����C|��{ ,]�ⵆCs7|����}���4��}w~��s���0�|_�~:���A��S ���s<}��*�y|:��dY?���௑��.��~+�{��@�qLՈ���|�H��&4�)���wؽ�6<y�cp�η�����$�alWr�A����'��8��*I2ꯇ���X8��ڱ�����zޜv��>>{w������:��n��6���{�.����r� ~���:?�T���}���.7G\ �_~��7n线�h���i�cp�F�;��Z��3³(s����`d�.�!�!�Iɧh4�� `eZ��6�u
�as���O�l�F�&�F�^�QS�T}�#-��*��_
9}��m��(�`N׋_�	���(�[�n�h�Q�ۡ���2��>�52��9]݀�M�=����g������06���-K/�{�����
��Q�d:J(��č\�Cx����l=_w4�~��L3O��^�9��h͍k�&����z�0^ˮw&����/V�u�m��l��#~"��W"����4��|����q�,4L&���W��̓�"���x}��JX��$���aw�n�!�nN�e�7ނ�wށ��~v����H�����FqH���C�6�6E/=�������l�8�XZ���µq�~�|���j����o���o^W[y�N� �8��y&:��%1D$IǼ����m��3�qҤ�^���ow�s���yݮ��˄��ek�T���h"�0n
GޟJu���(�nBC�R_��<����W�I�]	�����,*���zlQڗ)��冹m�Ì;o������w�`S3�f���F�brNA0 ������G�����$4�S���V2pY2(Z�]ޙ7�3��7O����ovp���ٴ�.�S܍�ʠ���aA�k�6R ���NI��N�\���{Zi<Tr�8��c�O�^�{1*J̍����@�]>7�Y�N�5�"��e˝x���ܑ��T���+�n��
�'�l=Y4.�X���p̶��&�F��6���E�Y<���3}�vN�?|�����awrF�W�:׹S:v�3���N:����s�;����O����� ��+1��_Q�F$���?cqQ��w]1]�Ѿ>^��SE5�!@>����3H���.�t.�<�7�8W}���;�ORp_1_�&Ւ�Ҋ9/�<a�;qP�b$�υ�P-xROin��Hw�� ���,�}:���Js��Srr�y9���ٝ�����O�;��r���9����n�K���q����8����n���f@��;���X��i88��(ç;զ�S��R�-�8?���A(�P��>	��]*�;��z ��RM�
s�'N�} \עs�#O��.���K�<��گ�3�]:�s&Ε����yМ&��qu�=��oGO���w����A9�p[^EFD���h?�+�d�vPh�l�{����E����l�>��ƫ�2�_�;� ^P����%>W�[u���ϬF|*)�^��s��#�.�#�<�ʱٜ�2iG'*H=2�=.�Y��=<#�-�����������+�
8�A��֘/S�(_�Z��HW����k]2����u,}�'7���R6E�]3U"�1ó����ڨ0|fÌl�f���Ay�P���o�ϩ4��� ��HE ?Ldn�~�mOwM��A����pr2��O�{_��N���IݟڤV�>�s3���l�������h�;˺7�`�Ԃډ��E�x9=L��F��Է����Z���K�ee>���	��~.��MUZ�p�BSLB�r,���G��� a�~/$
2g������H_m`��d�ԚQL�	�22(, |��,o���ȇǯ��)n��o�g�7����d�\N�
�����һD��0��1,G�E��0�"(���z����ץ��hj��Jˁ"d(�=���<�1Bm�h�����1�(��.և��js�U�T�p�Oi<�N@c�n��],I\)���֋�~L��p�(_z�y*"=�$lZ���(kGR���-��`6qFҾ��]�d>��> �2<縿�!���Gy?]9���0�X6�:C֗�]T*��������X�<�D���E��t�A�3\ ;���!r��W�q�(bSO*�x�������MFT��B�O��͖�+���o�'cA\kStWN}�������_�&p���n��:o�޹�o�b����N��ױ�B�[cS��+
0��!	!�j����;#�Ե�t?�����l���|���}7�a]D�=5��	�y`J�m����GiF,�o+$y���REb��~��S��� [��4q��ֽ?U�R���uO�����*d����Hؗ��^%X�����L�}�������2 h.e9E9��S���:;h�k�j�^�B� J ���d��'�]�-�]�v�u$.���k~�xM��V���N��U�M=�\�qhw> ݉�'�ڿ�F��`����o�
�m�mht�+��������.J�!�1��>��W;Ԇ��mq�-����<v��1�:Y5�Ad=mC�|d�=�7)@2�a���M+c��e,mD�A._�h�u�O��^���`H�jiG)��h��_'C�r���I1�o�z.1��z4䩺��WK�0+=_^&�^�(�j�%��4>�O�����T���4+9��5�� ��΄}j��G�p�La_����0Ǻ�*�ѮhP�9�N�h�����<mi����y�Y����C
|E��t)SiJ瞩��>g�sV��������b�3��.�����C��s�Pl 
�&q� ��=/w�:�0�u���8�ܑ�a�V'*����(��,�Td��w9%����v�Jj��<� �9㕧�S�F"]\c&��4#�d��#p9OZ��<��n�x�pu�u�5�����E;���<��Df+�S���6'�>� w��7u����S(�O�b�z��b$�;j? ƛx��縓9��3�t$�<�@���I7l���C�+*��h���h�xP��cّ|[ ]�:m��V��l�-���N-:�t�v���Z�����̥)�SxZ��˚�;�M<SA�ө��3�k%�x;��y���
F_��h\�W�l"8mJ~l`SA�4��9��Zm��-˛�߷�q�%�!�UF*��d��+g��4U^;�"�m����|Lks��	��KW�i�N��7�뢜2(5o��^�%k�z�FKC���8?"A7$}h����'��]GQH,Jߕ6M�0��\y��d�6��Z@��Xym< ��៻xw����Ȍ�$T�Gѳ��i��>�jt0�f��#��q��H`:����D[�/+��xR=�'�үw�l�rCu�[����H�EN4��Ђ�ܩEF��,���X,^+�u�aWj:�{��)�)9@�[UaW )\��ܠf��3j*��u<j<�Y�\�h�dp�\��׊�?���/����ϞN��r�	;��#���k?PBƐ���*��X���r�kp:%B�`c�^����M�w�`[ȧb�Ji=1Jh�o}����A_�����؏�4Klޟ�\�%���2�{�	:��r�x$�mđ@iZx�z΍�r4`�ά�h�:�}��p�w�*�ʇ�1l�M�C����]����� �'��J���9IN=�0j�\���%��X_� ��XO��$l0��~BO�,��h����n6�+��(�Z@&1���V,K��p���2P�(r�� �%��Ӡ;���x9��%��9j��FiA@���5-���Q�>\�B�Џy�0^�li���-�n�?����'���TR�8�.�����G6�`��ʃ�Z﷙M�'-���4}���+T�����]E�	�Mt��̝đ�6J��e6Q�0lW#�2)I�X��ׄWx�*|�<��'��E�����d*ޢK�^�Q1�����u���8�9tm=ȯ��ޘ��ICS��YtF��~~����<3w�DC&�A��&��
��s�b��mD#�uI��DG/�!���/��eP[y<���~��C��Td8�u����^Y
 N�m`�ɝ�|��7
(	D�.<�����yO�0�úk!J'�<)�� ���Nmg��S�Ah=E$$߶��o>&��@}G�.���`�t��@�'�\B����u�?}_�R[Ҍ��z�K�k	x����0�=�8�~l�1B6�9p����� ���s%�ИY�@=�*7�4�u���V�4�#o��S*���N��Y�9V�(b�b���	�kQ��;��w��@�3��Z��}ʊ���]d&��|��[Y#���(�;H/$�Y�$=l�;1_�l$5fp��䂁��Lii~��d
z|�&�9�_E�������sAڎ����1wν�sT�R�}~hcV��X_��-���qxs��k��x����?5��ˀ�������m����h�l���1��e����)�Χ�u�����f��a�7�����;[�14,Y(�I�����B8de���un�3�OM
w;�v� $?T́,rh��#2n�x�*"���7<ʲ�S07�m�����k�'�Hߖ*l��@����P�C1�;� ~�������:ݱ�@E�!K�r�����R�9!C��N���{F�v]�6E�
syL����/n71�+r�l|c�Wp����r���c�E�U���r;�t�8�cɭ�S�����N`G�3��;�NZ�]� <�������J����1P�Գԧ�x�@��Q"1�}�h��9��{S�`L! �`g�Ȏv���z�W����E� �X��6�q�
w_��i��f�f��߬�^h��oͻ�N���ǆ�wT��c	;H�$6�2QG�G�r�Ӓ����ǂaFo��pt5_-��IƁ�z��Z?]CȊE�|�1�նl����9����m���>��y�.�u��0"R�.�m(Q$�,�	ev`� �2�7������x��՝�p
Z��1�c/�!��༾����K7�a�޺ol��6��ͥ�t����|��Σ�5���At��ޙjg:=r7h.�y�6,�N�'C��)M.Ư;��3�:PqʛW������3%m:��b���h��2�`�^:Xn��o�s��/p�����>���	�&:�O2)�߬u��1��匵�9�L�<w:�w��10ʌ�p �C;�T�A`X�X*|��������*�9ߩ�=����3�Ĳ��zI���M��`�jTj~)�3�Ӻ�U�,�
�d���ef'4�Z��Y��9�l�N>t�0�ȑW��gW�����в&��L��m���\��RvC��g&?�����?��XA�(]�K��qb�]�����h*rp��;B�S��9!\��ݒ�>,�Č�Q4n��:�)�OB:�'{�,�6F��\;�6�|*S*]�3���N@b�_��P�2�!߶��N�O��+\��B1oCp�M�z(�!	�>�ל���\-�F
,��dq��M&p���aP�-�U@?Ǵd~2�_
��SU�/[6`l��� ?e �7к)�:>2�#+��h��LxaWV�(gp�!�aӻ.�2W�ߒ�!�Gz�P^���5�0%�m���p���՜�������&��~M�1��석ѓ^1�΢6����t���qi�.�F��+�k�y,
�@c���Ԏ?����v�v�y�q��c�A�|�9.�ߛ��,��6'(,���u��`������Nn��!HF�1&or'b�v��cϲ���\�ۼ[F�z%'�.@��|a,��:�9f8OJ-�{�3�`�w^��P1�e�V��k�e��M�sש��Z? QW����@� �el+�!q�x��T�� �:����`>�)���5pW4G������Z8=n�xݹ.�������Z�<FJ8���IW��X<3'���	e�I`10�I�ᩉk��'i*�ϥ�<&ל�1B;嵾q���+��e_A�?2 f��<�y4�;�����ZhvSk"��b��W*�f6.�gQK�m�Naqu�����,-����^�9�˵J���H�ʜ<˝��v=��q{ä��*�[����n���
�c*7�������t��&��74��ڦ���\0���EiWq�O�²���:bT�@�&S��ۣ�C�\j@ρ��a6�B�����*�>�_?����lp���R}h�E>Jg�v|�-v��A�<,��5��:��XH�E덞�O�6Z4j�#���o�k�r��q����6�`Skb9C,������q����dd���N+��xsw����m�(e�[HQv������r
g�e��؞�X�]�ֲ�	R��=��gD@໷e�JvrJ��.<�\�.��[v�"\���?�af�r��G�wɧ��7$��ڼ�����)?Y"�#�8�-�\���Wm�j��Ц��q��0A�q�l�Cԫq�`��v����S���+$8��$)'i�#E?��d��I<K��z	;|����7�w@���A?q��}�1=��� �!���Cy ߌDt=���[�H#ow��@\��yP��\��N�e8�g��Gl���-'�^���NYcrZ��@�Y�9����$	��.įXM=�K��ۘm���	������KÎ
s8l�M���{NY���;�$��A+[La!]Ej[E2Pj�v��o;��/gU��쮧{�����=���.h���&x���j,(��9Q���J'�"oqN�>�7��n��@R=#�w�Ffi(�DN��z���}�0>vl�@;�|��?�Xɡ.��)=����,	�:L)|畖�fNf�����IG�V��F�s��u���B�`��0�y��F��11�/8컄��L;�c���[W�PP7�qJ0 !�0�N�	�>�� ��FV�1EZ≊�ua�;���4|eA�9�k^��ɲ���4iN���
@NM<�%�-�I �b�#Բ5S���,ǈ֚�55��Þ՝0�\���;	c��K��z	?h�6��a���8g���F��+=�)���]�%=�"�cTɯS~_���b$��T�β�/�,x2,�$�1�������t��e8h�������?֥��uu��6͆c�cPSH��}��� _����]���`���*F�}ɗT���k]�&op/��?���`���i�4f<��v�KY�Φ
��6�&�>���kR���;R�K^���
g9���.앩�΋��3huV��w?]��\*Zh���}��qߧ}L������M2�I��5���;F����Xr�����*��On��F&�h��	}���DϚ8���j���#�`�5�pa	6y\���l76{<*�i�K�
}�}^~�v�F*}:5�0L"��ml�I��Zi�8Ⱦ��L���j�kl���hJ��x��R)�6(��p�8�8��>�1�F��L;�B��:��epC�����C��!�Z��?P6A��9��>���-�� ����0vfd�w*N�P_n,���'ܧ���#/#��^d�j�Y2�_۵ J5`���bP��@@:%hn�����s���"Ig
��n�аT�tp�㇥�"l������_���N/��T�|�{���6���MKp<��;m�k��������b�y�j}ǃ����-eҊ��t��L��~��;�7��e\3]7oc��,�ᛜ��� �]��tqM�l����-�I�(5�%4 ���C��[y����h��8zV��#� \�B��658��])wGc����j�&ĸc@۩1^�/%\rhG��\c��T(w��W�F�;�0-��//K|b��SШ���_<�p�8t��q�%�vT<O�@�8�kրZ=������J�Y���8(���V��42O�Gp���P��ڋ�i��G���D<����yeM�m�5<=/p}�M���p�s�'�L�;��5���M:��v��?���˖����ܘ J���V���C��q�@��� ��u��3��я<�:�4\�z`~�f�v"P㜺6���!r��)t�.ҧu�O����3���¬@?u��T=3�'=�V����:�d��I��/7�՟.����)������ ����p�b(E梙��tu(,���f��`�6�}�G����%��6�V搇����U�e��3m�-y���gp8��Y�Q_1�c	�&�S��8����9�F���j�jde��i�� ��$�Q��E�L��|,pm�pnߩ��"����uޱu|D�w��)qR��&?�#/'�G�p�b�Y좂aJǜbXv�N�H;�� YXt���s=�g��È1 �_��Z�S���g�����������e���g��>�Z1�v�S�9��ƜƋ�;��}�/~�@���J:���ezl�ӏ9��C���4Qz��i��q*LU^��	.|8&�vʓ���g�:�vN�)�q�^��2xJ����1�*ˏ�~JLgc>0�
7?Φ%�lxX��5-c����K�Г'�6�ҵ��[h��C�iV���m��T�^��L��b�J�$vA���,��4� ��q]���r[�-��Z9^ug������J<��p��ц�;{�m�i�M��軬݆�(^F�N�ӮꞖ���в�A~?�8;7�`���(�^f=�Ô��bg�
9*���+�t�ep��ģ�*f�� �:����Ō��І��d��	�pb>�{�kx҂�+��h)��C[$��	^��qlp,u�L�58{	Ό� c�1^��S�2MG.��t�����t?'�+��RX�`% l7�:�/.A�cU�̠V]P��k���"M�]!��v�Ԟ5���������Ӳs�VmAh����[�Xxp�j~Z�'Q@O��Mz����ڒ��ڴ��X%��|�P�.���XјA3�yF���A�>W�Z��r b���7��N���2L�cQa��hs� 9��\Z��q���qDY�iR��:�{�|#sR����>%97Tk��v�~)�i�mJ�Е3aJ�t���Z����.���z7�Y&�55���:r�L�˗����|mM�р������g�����Q���(d����Z�$?�P���^fB&�qdޘ����j:�,k,(O�{����њ�>��������w�r�}�6'�
|]�ʭ<_����c��1�z�x���@F�X�i��Y����-���&���j�'��*V�l����;��
[��l�A�\:N쓟�,�v�>97�2��rm�m(JS�X�!��:̢�W�K�#�#�w�O:Z0�{t��k-?�}EI�z�X���Ind�.'�hQ�J�Kxx�e>�x�Lc��F�c�n����D�F�U�X�x�9S����i��xq����#�okb��2%⌹7	���e�`�0��f`t���]��72&�)w4�<}D����P2\����䘔�c#/ڏ��0�`7�s9��n]���]J! ����<+���O#�J�]ո���;��]��bx/^4�H�7����[k����L����ߥb?%��	�A5ί!͌��Z�Ff���3�-�Ƹ���jc/�]��f��#a������@W�Av�3��z�@<i�ok�������㭧_�Y
�ή�;�x�@��`7�9���re�b
�H.��t����SZ��(q�t>(�]A�,�,����@�m9�!�)�"d�&z��|�@Ä?3̊��?��O	���0x��q[~�f8͗y=�����Z �[}��s���wvQ�+�A!*���������*8�}Pwx�Xy�#~�i
��s��WH�K |l��F?���zۑ�k�&czǹu����k���J�,ԭ�~?�"2(^�����x�׍�_���t@�.�1���2��<��2_3nw݉���b�NC�����~s��K��'C@� C�:?�6pQW���,u�����mbu��_}�m]Ђ2�nR{��mD5�6���i���Xg뜯�;����q@o�h�U>��d�Cs��];^�}�9Z�Y��{k�k
8=%�bZ�V�{�Z|:�"�Yt(�^�r��Ki��F�wټ���n4���~�lSƵ��&Q��O/�>]�� R���ɥ���jť����ei�ے�a����Эs����ނ9��m����y>��H�WA������-��zdt���f�r}�\�IU��!q/�BE�v��]�N7a�|R��I��Y��89�Ii�S>��B3M��DNkFO�s%�i�~J62�̖�a����4ɘ�`��U˗����$,:Mb�x,�Z>D ¹c*/�{������	kFLcmMk˘�ә�]2{d��ms=�7qcg�M��v8�gfMC� ���&Aα<5;ro��&(���1>��Jsr���F�y���xd5:�e{��2?��	��X�1|��?
Rmi0o,�	g�u�mq�#�dF�������i�w^�{^:E)Mr��p̂V������
g�Ww��PB~"H���&�4-;J�A���>��c��Sh��Ø�./Wf�����U9����&1��M����"��;���b��Z�YmkmmЌs�t��ơ-k7uE�g6���>ǃ>y��i���8R�|�kM�5�!����Q�|Mjm���1t���
Hc��ͫ�}�'�ѨӬ���s*��w���6�`y"�R�j���3a�L�;D�AA��c�ɾX.�S����B���=f1�~#4G^z��'�x���br�2��ɘ6��Ӽ9�2�~Jn����@fTd����I���J��=�]Z�98�K�o�S�l���߫��3�e͗���B�8��ba5���t�%}Z�"-�5���%�%�[
��t��p��� �Nݏ>1k8�6���l���v*� ����W�b�T�J�]Y�a�u�[�]�2Τ%���L�*��^�k�ǉ!w�i�fpᏹ����jQ���"���JKOkh�����?���T�BK������� $���e�Ν{sꬕ={]jszI[xd$=��F��Czn��"i��N��`S�i>��qqj��L�Ә.��
	3^.s��Κ&`�B���r���Q���Dh1M��F�t��Ƀ�L�=��i���F�����p��6�s�{y��nȦ���2�e��L ] C\T���l@���9�-kU�_>|�Q��r��I�D�AP�#
�q� O�#>�OE0 ��-jբnYK?�e��\*h���ۨ�i������Z�z�E�� �y2F���S��N��_�E��ZT+��0�~tt��.�ֺ��Oe���E�~��mYy�kU�8-�3d�@��a���D�X�.O	�+O�ٯ��-÷���(H3��9=�w淞�pɹ��к�y�~�`rݻ&q�m�/G�+���v��8spZC�Ke:���\1���� m�7�3�W_��nr�`�s���gm�%���b2&߭#��S6��Z�g3U�8��z�����T���m�6��A[�I>w'Ѻ�5������xv �u�J�&f5��e�Du.�˂������9Vus2��VNZb3�������g�w����>g3����N����l���w^=�7�^�1���7Wіe/ZC� ��X�{CϹ˕���?9��j��T���P�����!s�H'�7$���s�R��j'R�<&K��L�P���5nplÊ�i��AS+��9�>�T��蹆޷���r'P��+�-i׵�G��(xJ��u���0�)F�Y��lgMO�)��͍}#4��,�9���"��8b���b`Ǵ�p}h1���Z�o�:�t!c�9Ր~�ZOG|Ť4��2���O�����9�j��t���S�>#g��HzV+��Ҽ^�����c��8�!{Fϯx�%����u7��ׅI��|�>dzi���j6�ߞ��D]-Т��sܐ�H�H�P�(���?Ĭo_k��F� �q�nm�Wy<�`��{�u��0@}'�ؚ�^�R�)���"h_��dDZ��kR�ԩsa���D��z�&��ֵL���u�Yөl�%�S�S��g)d�Bc�5�l�9=�~��i-���g�-�5)W�8	:T��Z��X
(Wn���9�6����Q>Mu�H��@���(j��i5��,ke�tv��l����6��%�o/*�\3,:��`�UOR�h��U�e����1�<9O� �t�P����Y">^߄�=F����7+sLvi�|J�=�XՖ���@z"������ྜྷ#��R�e%Se^MA���
�m������E4�����9��b����o$��"�I�p��N;mo���Ӏ�7�hU�B���x}r����l�S��x�29�SB������}�8v����m��x��ȖvP(r����aW�I�XJD�M���6�ō�t[c�1I��m��K��k����Ssf%��NփS��}�OD���'���.�cI1��o|Uq����3�Qu[4��Zʯ�'�k�8�+)1/�]}���w~ڇ�R0w�+c�P�%�,Y[��\����Hs�]tȐc&\큟XF��lG ������iN��4~�
<�k6���|M�G�K\��H�#���|:�j�6��:+���a�:͊z�\�x��)
��qY&*m��]��/�as?AO\f@y�(=0:f��`żDٜ(1�u]ֹ������{K���}*��7���]��8�a���G��Q7(x��e�8:�2��ć��h�)Y��n3]I��q(ul�,'ә�gM�N�	����t�^k��(���	S�R|�j��_,�@��`�&�������'a�@�X�d�e%�A���Eγ�H�.u��l��m�� �S��]�5��=0���X�`��m��n�!m��6�`���]ڳ�.r����Ѩ�&��N�gU��ݢ��Ӹ�7n�v���:�t��!\3�ir'T��ci�Q^��9RN��I���N�81�ֱ �j��2�j�2u-f�1ū��U�P�[�mP;�w��k+����rH}?�_̨����KJ}S;������_��k�e��\5]=3:��ӱ�����N&�T��I��%hcDI����Ām'9�_�̋@cEh7c��d���%j||B=@���%�W�T[T,�1*�ge���7����-��,���`���ڪ��h��&�����u����m���ak��:�ll�U*M���M�2'�� 
�O�~n�{�&�s��uEN*�P� �O���E!�����zTL�V#Gh�0����a#?�ڈ�����q���5Q'�$qM�f��1y��A�2���TrG����i���'�ǝӌ�]VK�a�s��L@U�<���D/{̜�xh�K&�X�W5=V���ﮭ��ݔ����K�4�_�+[x�70�g��ԵhY}ǵ��,�,��GP�'(e��B�"@�(���=���&Z�����Y��p�3�˖�Tɷl���x*!&�ǐ1.S�2t������s�B�yE�#P�N�DH� uc�gIMl�!�u4��K��� ��H_p�}3K0�Om�ڑˣ�:v�ݑ 3���ծ�0��UM)����D
S�;/P�SZ����wa���A��S�n�b�C�'j?�`���Ģ�Q2�
J�uQ��ۏ���@�l�0��Ӭ	;�ߧ���l��mP�i��%�M��Hc �����\�E>2���疞u��d��8lP�l.q���Hk��,�؄�#i��s�1/�Ҵ�9�ֱBdCei�b�j:��$C>e;��$ �ԫ��X\�M��;v��Z-9{]
��5�B��NlX:�x��2��P����1|��#钾�΀%E�hm��L�c}~�y�wt�JOL7S|�¥/N�@�.��}�U������-� c7I�3�sJ�N�[>Ќ���9CF�d`������K����|�4���� �O�A e�Zc3�uHE�֖���ؾ�|o��R�D�h0��d�� �������B�x��@�QhlF��*��ԇ�[���}4��^Z�T��']�fVh����B�A͸�����L��9<����r݈��T):'�#z��z�̲���ui���ڕD�I<m���sLΟ��T�����&cH�cH`³w��`2�U;��"a���>��y �ӥpjJ?��1A8��	G��Hn�тAƋ��/,ՙ~��x��pm%V1���������tih�������Y�΃���d����`�� �0'�����o��vԣ]���3�^� m8gb�`��ؔc!S����2����2�߶A�~.K����N�{i�l���駔���@���^��m5�t�)0/���xF�`���ӯϚ-��I�U�?`N 7H��Kr�ă9��B�6t�:��5�^���4�g6/��=���~k;�d9���!F/)��*�g1�3�)^eKI>�|.��Q�CL��^6���>��^��;� [�΁�D�p=����*��53��=ȡ8V�@#���H��H���Z1�싉���W�Y�ʼ��J�ªcዱ����g�b!�J�_%+s5kӶ����J[Ϲ��>����C��n�(��������k����N�)�w�/=CO~Q�J;�$�t չE��ͣZ����-��Q�[C����Xi�xt;�9_r5��׋`/|�j|}\�(�!gA�ӓ�C�*�t������\��Q�,_*tcʡ��3鏦C�@�P(�25��/>K�?��UeU`���O[�L��g� ����3�������8jqk����/��~�Fۑ^$�L���SY�u�zhj���h���X/Sy�����ն�cM#Nes��o�n�	<�'�Y� t��j]�Xa�-��%d+R;�Y�b6��l��0-�*��s���K�c
�ag��{�pɀ�m���:Ȳ:_U������m/���[��~Y���V��hv����%О7is�'�6U��ld�q�(�7��+T���&��x���s�/&b��(s�0Y�==Byd^��Q�\�\U�
�.	�Yf�_	jN�����7h��
A�g��Z�Wn���P:�ju(� =�m�ϵcF����k�����/�]��;��(
ʂh�R~�Ҍ�Tp���(-��`����.��S���,���|���%�v�S�����Ys��h�Cv�9Xx����� KfU���
N،9��vB��x-���y���@� -��v��O��M/m�x[�h^&ܹ��.a�8�(*�Rr��_����>�{V�d�y\������<�\�隌9M �%��Ȑ��'D�L�Q1���H�A;,qTitb��VO��:�I�)H.z��IZ�,	ް���N�rA�G��E��*�p���ˣ��r�X��Җ\U[�����'��4�N�H�;}	0�/�j�/�+F�2�\WzHǺy�������5����_WG0�X�#�x-�����hM����O��_����/=lc�3?�`��HÃ��U��>����pD[��xI�̺��Rlј9�ʃK��e��С<T:�Ij;m�]=�B{�1{Y��*!33�f�F�]��z�1��F�ܱ���޵8��N�9���	/���� Cbٮm��sF���@7��%h�s��S#*�;���T��˵��7�n��fs���#~\��x�F0E�+�}t���	�]�qL��ZZ�>�s�y�B��Xɀs'L���2#���i������:>�`iڤ�i�&x奛7|�م}x6DL�{k�ޏ�"v�����e��j���\����kv�B\�E�#�Q���ԜGy~\o�:O�U��N#>�A�3���LT�� ��P��]�W:���[˧�����;�%�b"�Cu�N`�vpɶ��7o�����@��p6H9Eӣƌ�c맖n�٥��p}4 �M���9��͘���ԕ&��~�����o!���/*�?:���t�Yz���ޫ���v��qd��0Z6(h�P��tsm<|�\�gm�J#2�-��xz���˝'��M�&!�c����ӹ�BûA��}�;�]9?q�9�� �sF���5�{�ft�
MmJA!����.��e��a�V{���wp�Q4��^��v#�рx���-z�"�H�U=L���L:q�?��s��5��V΅�$������!5�z�% �o��a��kN����kOg�������-�����}c�0�L-0��M/hˉr����N��7�� őG�^7�[��t�9���6�Q��3�N	��]"X��� E��_��^�h���	l���E���Y-�?����BMט���������=m�_���9$)��Aՠ^��( -I�Ķf��� 3(X�)pk���$;-�K6���D[Qȑz`2j�6�)�ܹ���<nר�|8]8
tҘ!2N��%��(`�:j�u�����^� Q�ߦ�4(6���I�iLT��Z#*3�Km�TR�X���&QR�{��Y��ԕ�1u-hu@-.?��M`��W�����2L&i��?����i��e�
/�l�O�d �*8���$
�
Sv
d��>f���}%����u�_	��zfҌ��s�{ۙ�_0�����"e��7`z%��dᄜg���L�А����<�^^B���ߴt��3�\�����G
�}�1j:����I�!��Uc�����#��jT��2�H������B�������PoE{�l2����N��҈�>k���!��{6`9�Ge=�@f^����i�m+i�@��B�=���5*D��J���\@��/���ڧ�mMN>��0�t���bF�=���M�+x�!��?��/qĖ\7�x(p�_[�m�bM�5d��M�\!SkقϘgo�^n�9��]���KH��A��o�Y��n&��:]/e���45��k���`n	��`�K�5ϭ����ށ�-|~�B)��V��G
�Y��e��vL�a��Ig���Ѩ�e^q�{V���5c�T�jQ��9Zi)�&��[Ѳ��X�c�����Id���mZi�5Ҋd�J��������g�`���5�f�>�.hb֋����@���	��׭��ImW1j'��_��G2�����ޭx�|�V)�l,�,w�%����I錿�N�ڲUNE�Y�G���Xa�ab�Ƶ k��˶�O"O��ycy��%��+��VG#��r��^)Zk'���+��^�<����:��s><��n�a3Y���N:�uo1��?��tn��^c��5��e[�*-XZcC0ܹ�r�x+��?���� � �O��`�:MY�:�����H���ôkl��m�G>:#��m]ԏ݆鞅�s��jX�6�ǲ�y��9zΒ��`�+gl���hאW�?:�6��a�	;�=��h(}�	��¢ i���cZ���������N�)e��S<�ſveu��SU�[�v�IA���W�@��(��&���+�hFT�型4/�lG(��Km�"���h;
�%Z�N��QVLC����9��<
B�p�-�lN�f�bT�8A8V7�n�?�~v���j%��/���}���J/ќ���׵ ��\�"/i�Ḡ0�c�ш9��v�O95lFˑsT�1h��څiΚ�+��l�{���L�q��X&%BH�[��q��t�?М��c��HZ��8���Eqg�>������(��\���<|��%�'}^k�ɲ��\*�aI��v�=6�83�]�ܕ2[�1��J�1��>�l,a���*LЛRw��ϒ����\�)*f���}�NSK#�Qs?3v\�F�j�y4^�O�;�9a����)�4c��1�zH`3Q�^�<�Ȕϭ:�ίm
T�b�#�LF�v�e}N��}ny3�ޱ��"栗�:�#L�-ʮ$���d肚=8����ǣ+�`�64���K���t�bl����@Yޏ,��F�\!�"��<lz�����3�ݼ�6�3�o�j3~u���ѓs��尔���Q��|�2�}���/��i���'��������eЇ6��eW�Z�1��XS��9�ڈ�r�c�����9;�bXk]��蓾CȀ����/ *B���,�wI�u�S�\cXNLlqO.�\՞��L��f�cB���0��/���8jB�fP���������3A�}���fEq�ɟ�5Ch�7)�CC9�L������&{�v#����x{��s���� �|8�|di,�:�k8h�����M��g�V��ㄎ�>:J�X�)�_�>��G�����I�w�b�H��������﹁��!����k�nu��HM�̹1��*����yᲰV�DT��Sv{[��RjF$�f����M����T��b��E����bUQ��L�jjr�Q����i�+�VB�d9&��>�}?$���b[0�iGA8��N�]n@�a{��ؔ�;R&N�T$/�ݓ2���ŠA�$?�>�0��U!ټQ�
���9?�Q�QI�����%P���	�����y��m�+U�7i��:�Mr��׍�_����jզ+����1�_����4��u�21:-��ߩ�?F�k�|��a�]Z9-e�����>���S��S2_��ij>�i\ݗ��LYTYc�&��S�*s���\/��3l��Y.1_�����

i��W.2-�:"åV<��W�Q��:oI;�����U'��!�g"�t9!�`�Sx�ݜ�f�"��A�E�5�0B#�5��e�9s����tf��$�Ir ����>�_Y�Gc&1�dov���L6%��(����u�M�.k���L=��Zus��?�-��c�k�6|������kjn}cx\��Ǯ$k��vdje,�}��$1��i��/k��E'p��^P�\��.2�x�c/M8(x�e��ɤI@����J��	V7��;������b�xd%�j*�Nh�B�	�S �#<��b@�m��M���SC�l�י?`�m�r��sx��@�>@��!+t��0p+,3��c� ="�]Y�mK��ԇ'"���]�����ef��{c0�P7f��q�m屎��u���:s�a��p��>�ai�P�{zf�h��u�m1n��l��]X|1�Z�&~Xo}O4���j�G?�z�̄E�EGW��V�pi�i���I�R����u|�Iawpo`�IM,�e(��k)�s�1��\ԡ��:���Ō� �p�xQ�Fd��+�i��Ti&۩�N�c�	�6�{ G�2x��n7.����2�>e#T5P�p����@���<`���-��>��c��gR+�sy���3��||�<Tep��N�)F�i���4Z����،��p��s�EWsZ&C΁p�P���J�H_��c�,?1>�(����K�~���b݉�䉉[EQu^�آ/�֌\g�m���>���g�>Z��_��i����\�|�bQz`�}�18>�C�,�&�N`*2��d���Q����Cj��ͬS\+��&�V�mR�{�����{��9�r��a���Mx��N�0��c)��Q��i}��c�J'��;�B�����ږk!L�3�^��~��cP�!�8HtYRi;Y/Ok�����_��dͩ^N�.���|(SN�Z�˔~�����y)~G�P���B���O�4|�d���e�.K��� ���?��'{���6a�m:"������,����jWd��hCU6����k��[�WZ���k����9~���mc�fsm�-�Ȁ���H��7;Ȃn�;���O�S���jI��/L���W��1ڐeW��Y>��vY2k>y BQ�OL4�����2ؐ�ٳ�!:�Q���1��d�jr�g2\s��.E!��|/�	K��Z>�`�b$a�����/p`�f��f���Ȣ��&��&��O�I}�WYE�+��*���j�(��?{ߢ(��k����gɝ
����ѽ׬��7�I�梣���7i�vzB[�:����y�%-"e6���(�>fBw6)*�����W�W�3	�Ό�>����g@'�5��1��%�Vn�%��Q��u�>�k��z�6�÷cr���"F�f�ה]�+k���	����xm�_��tH�m��%�iS��{���g!u(9��R^Q#��Bf�k�K��K���阕F¦�%pF0D�՛���y��f����0��p�GF�т�>4#T�>I��Z�V�o���PD{���L&%y���c�h�xm��~�g	s �i>oFaV{	�y��I6V&�2|��躮F�3r�;�P�������Ʊz^�F�iz��,J�򚇸���er��WE�l6�F�\�Am����aB$-�~9����C.�yd,��\����8ᯔ	�2~I�>i"}YS�z���a����121����k����~��}2��R�ˇc����&�X^���S���;�2��?����I�g����~oh*u&��@_�a[!��;����P+�t��!�5����%��^��
�9p #���NNS��hS$Z>#u9|��_�@��.=� ��YϮ�d��xq:���n��u^�>�.�?�JB��
���俢���e{p����}q�8��U��˦Qq�������aԹI�e&�|�t��3�D�pG����z0�Z��=�I��a/�����mZ��>-�T���\��N�(/�b-R�xΞ%��~��FW��/%��Q���A{�N�X�����M�(�yl�G��ؑ3�^��X�i��Ŗ�A�m{��@�C'�JmB���h��g�>oZV�^����}ޤ����mT=@���탃zjo�,9��}'\Ҡ>/���E_�#kaS�r�sŖ��˕�O��:6U1�K�����l*=J�d|��_�䍪�m��pQ��Ԕk��݆<��&#��#�)WnA��������<�w7�5�FV0�w)�DY_+ߺ>�Q!I�NEe���6���Uo�eZ&8��qc�	�h��Cu�C	����0�
�XW0N�B)T�0�C�!�T�7љ�8G�z
^�C�ܢY����L�G(���r|���Z���L����ޢwn���]��֞շ�j%r
��<�W��r�m�g�@����{�����~|k�]Y�>���w�-'+������>���{118@g`�-��}��"4�o����ؘm�z��@���~Ļ���MauJ5j��N$�$
*�ĎOf����׵hІ�[I+Ҕ�
$Y�i�R9�1t�Un�b���u���~��5n��	��A/A��4:͐1��Hq���L�q}�\|�쯸n=�:�`��t\�WH2��M�����5+*�?I��a+jaڿ�h��|�Ӿ������Ss�����s�ͯ�tu{�z�����v��@3����6x���ظ��῱���m0@a$k�8"���7������w���r�؋.�f-���)���v�O��������[�\�����I�^������.�v�
N�Z�(��\N��>���4/d���]��]]u���Ø��ϙ1�0��Qx7Pm����r� 00���y��𜑃ܔUܴk5��8<�;���4�&GF��#/��y�0@Y~I"��yP�{;����>�����3�4��e�H�:��[��g�H�
%��b���n�N�-��o}zvov	�������`5bAӾR��I{p>�L�G��Zg�w����ɿ�f�v�5��X6���5�K��X3'���d8��g4bJB�0��:�2�42�\�mZ垙�J�Ə���wwI����������d����W��Ll��K^P��̨9ݛO�{T�j�_y�����`���;�`9�C;O��qUF��H���1"_�q�!�U��0/��F�g�(�%Ώ��l_m�Eх�j��~�vu�U�K6���8�c/n��Dxkp���2W����(���{37#����+3B���G�|@�� P�eyJ�A�:��n	W��؃�`�m��k�0��^0�`���g�+��'��v�����X��H���]�˱B2h����*�Q1�b���c)D*��F�p��ӈ��j��� s<�����NTiˮk�x	#�9O8s
̨Z!']W�S(E����c���>��:�hgw�;Z;P��v��B�c�C���~w��/���N�1�ePôa_vZ]dK�72�Ս�&��|���m�)nN��8���~88�����ٟ�2B]|��������G�7O�Ǝ4�\(���!�k���rBhܻ7aT���;y��82p�8u��ߚwx����u�Eo�õ˃��щ�z��l5������p>�O��"{5v�a�-�	�.?	�>�O=�?c��0��~{c�}n���K�T� �� ��}X��o�݄�,���Q�[��O�i�}���+:�"wx��_�t��7�!�*��?�*D�"2�f�%|%�z�2hN�QZ�9c4�O�oF�Z��4�|r؎�� �$|����3�JE����^~����������z��Ѽ��8�J"O�~���G@�̆e&�</���������Ag�	����`�.6N0�k3�\܎�o,�E툸B�ʢ�cr�|���k�)���:��_�W�s��%q�P �$�������h��������������r��H;)G2�q�/t��F�W��W�]G���Ψ�l�Z�+K/��%��u�;�E�Z�~�����������u����S���V]N�ނϩ��������&ʯ����ϏoAvQn��_Dy��[�2�gZM�y�q1*B��|�zU�Jt�To7��������<^�W^${�~U�bd�}��jiu��%�����?,��Xzp�.��g���`�a�~�F�F��¼��,��W��X�x�Q�%��g�s���<��p��@�	�9��8v��&��7�D�&9�,+_���Y���~��l!���J�PrK�f{X��.�b{�ƾ����X��
m���y����.���唁Kf���i�
����q�� @<h�3U�wm��XHp�S��77�F�Y�͓���+����Nڷ-G�J�Dq�k��aU0/����)��Ω�Yg�����i6r�oK�*n�����xP��P�Z�Em٧z`�9>�WQ�,�Sop� v��U؇���Yn����q��?@��i�_��Qͥ�?J�`1�6h<F���{�}�g ޱ�zW&m�.���o��{�/F��OG��s����|.�)&![SֵN����Y���n�u��\��8=�8_&�S��9~���GX����;�LI�T��F��EΑ(/��N�Ȝ��e����ߢ#	색���_p�s�,��*�b�����u�y@��9�62�o���s蘬(i�����ۜL�[Kt�Y�V9�6r�	�%zx)�=
��KL�����_ǖ��V� �Vg����E�@
�&M�kVXcށJ3��qr9�۽�Z��l�}8�������쏙������>�����2O}��S���ˇr���(�ߒG�X��+~tk?��]�	���9���ɤ�?�����~�x�i���y%xr�d��^.�����kR���_�5���k��`;NΩ��?#|!�ڒ��@<=b_3'��m�e�M���]E<a~�g� ����/N6��+�v�&Zv��U��2�y�#��d�PC�_��I�	4��(�t3|T�܉.\��3􃫟R��� +�Q��r}��0�ƺ�ۻ^s�D
@���926����0
P�k����Je�U�8�#�����=lt0A����2�X�s&����R�@	\�g�C�860n:��B��HQ\"��TY��[7\}�������܉�hX��Lb=ܕ�3���\�M�S�E(+�_�}�g	�����NC��ƕ��}�x!n��<�RḸ��O��:��'�Zy��2o�[��$?a�*�X�<�>x#kɹkg��BzV�W�s��$�]�LU?1��d�̕�����7���wFP(�˗�����z�7;�L[��\#�|��Z�{%����t��W�O3r� ��F�tR7O���u���'�y��N�@ 8D��o�F��#�-�7B��,���a �����s�`Fܩ���'�����l��˵ڡ_M��R[s�t���/������i�)���ia�50����_kd�ui�{��]���3j�W��`6ŧ+U���H�a��p"�zd�kHHYL~�V��8�#�>���]�s�	Q)p>��ޑ1�3�h����*��	�a��(�Ib8 R^���>�I!l:�H�m�q��DEy��4V��xӍ���7R�S�c�E����@rWlo��}Vz�:r�G�O��Ԟ&#ƾ������H>��vel���zjD1~���̯t_���G��wt�wn_��{9�87�J�4�o��w�ޮ*?�G�0����j�{�l���C4�[�h�>�Fv��M���Z�s�E��P�d��8����[G^�\��=�};�է+g�zsM̧��9Kǧ�Q�&y���d�ƚ�^���� ���x���sT2�k������Nv��/��l��s����mu�����Z�0O���=C�6j�'�"�Ʌ��LYx��}J���-ʠ�{�)��nl9�����ͫ�Ki��ٺn��w�"��œ�q���Z� ����F4>��͗�ox����
/o���[�����I�q�9}�f}q�{��se��ds�7T*Ց	�ѹRى��ٵ��њ�L|�7h1�]i?�G��P�rţ30��n�@^�'�X�e�|<��:��w����e�֑sec�Ú�̩����1�n�;5RmZ�X��m�<@�����2�z8!Ԡ	4��L�&���Pc�X�ƈ��eMl�0J��h��zg���X�}Ǩ8X�V���i�NT��z:����iY��w�zØ��]t{�������n<`�u�9�+���)�$�(y(F�fz��e�Wj�MY�$;����E�c�A�2ve����g���Hq�E 8�X�j*÷Ko���M���z�W�����ʣw�}��H	�J�h+�+����g�>`d�P�gM8�H�BU�h�rsާ�6RHU�uOA���,���F�x��6��m`yj���'҆"��7�C�W�������>�\�s�l�c�I��~
�O��F��&���-��BRn��<mD��+��r�4J��JI�v�3����z�=陵��ݡ���q�BY�?.�6'�`�����W,-�����U�w����Xf!d�8o�?_�z���5��15�_+����ۍ�+���	��#Ɖ��{}@v����2ƥݕ�H�����c��3���М
6�؅&z�6��uW���-M��G]-��B���5~��Uk5NkwUR�b�Cj`�&F��1w5�Uc���5<{�� �Wٝ�� ��d�tucN^�y�0O�� ��G�D�a� mC0:jv/�s���0��n���N���-�5��g"e� �u�t�(�H�l�JG���1�]��q���FNr'�Ү�|_̋�|���Ї�'���/0����	�)k����Bm�����Ţф���6a���8�EX�8��R�~Ҡ=�� �ao��(j�d�Wa��2}.���2�lH����л�L��F=O�e���l�S��-��>��bU�|���ظ�G�p�+hB՚v���ݑqcu�s;�AyX� D��}��!�{��jleT�ww���ٹ���זg�͆�"���Ҹ�����"�:J5�5�����<���_wҲ@�/ۦYf湉�u¯���T2h'��Se���3��Dx|�m��q�^��Soy�e�Ϲ�L�ٮ�2�r�B?��]9��D�%2�@��\�
�/��	C����>v�{㍩n#>YӤ�C�~§Ć3��N�[//f�D
)�Vy&T;�$�<pq�o� �{��
��� !��煕zԨ�	��aիbE[+��Aq���F��w��
°uv���^�:b�o��[Qŝxn˲Ҙ��GѡN�9���/�ַ��N�5�)4j�B�1������f�6r���ٌC����K�=��:��M�2A�l�F}���a ��:bp�^���ښM)�	)���m�����(�`��1;:�eצ��p˸Z�I����)��\��uI�c����{R(ڊ�҉Hg�f���*����m�4sa˗Uy��w@�������r� �H~���2)�,����V�f�]=�����WXc��/XY��B�H�ǉ>�gu�����6�D�=o�����!AE�Js$����uQI�j�'��X��͚������]e]��Θ��J�'�7ԭ�~�4&yF�P��S��v���)�N+��o�˸,��^����0�C�B '���������V���@�y^7]�b�M����f��}�s�mΖ�F�#G��������c������]~`�T�7
�0{|�8����x~&�R 7��X���N�q!�_J�P��@��N:I�]��AT�%60��a�����h�ߵDH{�R������~�U"�Ey�ۮn+��z��T�Ǎ�rtW��>����j�<V��1y~��a~a��P?�adD ��\�J޻ZV�Q|ơ�\E��D+��Nk�y�@0��W���.�\��~�O�w�o���-��֐ȓ� ��ﮰZ\ҿA��?�6YH����\��Y��wmy�m���m���~Mq����\!�h0^�����q�]�i�~� �����j���UჂ�r�+x��j��|s�0�������}{��$�;��9ⲡ�m�G����
r �]	]W*Z�21��q߳5�����j���t�> �����%*��|i�o�NA.$��V�7�y��H=���Z�4�u�L�<p����o��sw�צS��W�8=N v��[i ��,�߻��d��&¡?W<�����fl���%.����)T��y���.v,�E��cgK3
�V�4��b���~�׍r�?tC���F����,��]�s�]S��ѴM5OX��,�������P��u K�/��Lx
)@����yd��Oz�~+���~kٳ�������3cT�Gg'_n.��`s��go���5��9�d�AU����HY�#p����yQ�y��N�+O�t�3�5�JmF�S���i&g�z�=e6[�[^�{M�ӏ�1�n)��T�M̠�q0�W�{�:z��qK���{�i������3ǸZX%-ٛ�'9�Vt��ў����5~΍Wb�ä�p(�<>6�iu�O�0'COk��x.�w�<��t��e��6�
��ru��qe$�:�d�V��'G
NT��w&g��7M���]+k
:�Gm���X����zYc<Y�.��h$蛐�*���R=�:�y� []��2�!I3��s����YN�������(y?r��9�`���%���ՅMuɱ�W����s��t����/:y��z�+�+F�T�Rn��7dp�uba�|^T�׌��g�� ��}�o9g��|8�/
�:�*�"�R��kX?����"R�cG �..�S�\<�Qg��
4�,�Sr��I�X�f�*�&���H��Y��ay�mY�Y}*�m;PZ�X���9v� ҬOo�q�����w�G��=��/����c�6�wƲ����*@+�ꀼ�j�7�;^AG�K`�c���e �]�	���]�h۹9Lo�k��%0�6y��� ��&���/��>M>�gv�W$9�dn���ʫ��.vtE������U�>D�\�b�\��UqČ��s����G-{��,z<�#�Fx�I��Y�d�R�]<�|�N��~�8��}��_G�+�E�xN�<l����y\׸�S�.��t�f���?�Y�{NA%D�9>ƳbU.�q>��^��|��Rkc�=/8��VL�~� CO^��ф�^�i�*�g�eo���r˻X��y��`5���X�j�<k*�M%��B�~���LV~2�~T���v�| у��0`�oJ(=N�m�=(���\�A�N]��4���-�&���b������c�-0�_h|�	��#|��#�yO�WGvr��S2��_����r~���Z'Z!�a��d[�͟9d\��F�M�9R�mW�� hT5�2,X�w��k�,Oi�$Jr���� �c(r����B���L#Q���G�O�։�$o��xO���N�Z����j8}����x���Em���{�W�Z��>7q#�B��P�2]{��`�4���I��F��ג2��1<[|}�w����	�y��D�ȶC���w$'��'��:�L�3���;T��8���\(2����ԖGϸ���5��Ӊ�b$��p��2g��B��X�>�)����;P;��4����2�6:�猲�j�s�B���y�:r�UF���1�Nb�4�>I~�M]x^+S��,z������.�-�n�N�#���p�'}�����0�"ԋ�]Z�����iOR6wb1��mNI9���u�> ;ܙ҃2���i�Rt\�p*,�v$�J�i�#v��I������;���5����dɸf�"�w���k�۫��M�<[���`KT������HpVe枎ٽ��
�o�3!���h�y��S��ȞO��,<�J�?;g��;���Y�bu�)
]�»f_�┻n�Tٳ"��"l��G�����kqă&�/WrN$�~bg]����]�w�
�*Q꣜�� ����*(���^�Ჵ�1�d�9�y�Jك�;��|�t�281�w.�p���2v��[C�g��cZ�[N�eK�� ̆p�&��{�ּP~x)����4r_S���b������B)��}��i	4��,��a��M�0i��;��ID�4A�5ٯۋ܌�7G8ļia9��`�����Et���S㽚�d��#�o0pjZ�ʮ����<���������hO.��溈Y�V�� G�E���Uc����"b!�]�%��`�i._�&����M�A$'wD�-����ѷS���>7�cL�M�����m�W��OfoL�1&��D��Ȧ�(�8�S3Ή�	��Ki)r�S��rk
}g�9�qu�jQ��-�sȸO'��4���O������\��*�>���̀ �؍Ѵ<]�O�!�[܋#^@��Ou���F
�k�ASc7Jc��b�Ft7��=�]p`��W6���*~�EFS��֍�T��oT���l�t^��t�*�uթ �c h�����erޣ�|�@t,��\���8��e�n�5�O]*;a��w&?���_5a���t����:����P��;�NN�`������S���5��U��kW`<�<^������|}��@����5U�^;d���	�K�yjt��T�ڪ�}��O�#%�%���?��IhD��� �/r+�6�X'"����}R��5�ЂEk���,����&����Y ����e��>dy�%懁�]]@�s�
����va���'����5�Mm{bdY�[��������0��㿝��? ;�W������kֈ�w�N�I�{�jd�^��A^ؑa����߃�Z����x Fw�7.��8���{���I�ڐ�e�^�b��m�W��1�YD�4��5�L���pJ��*b���]��I�K�'\}����NTiz�`����;��m��{��1�:���:bO���s
���W��'چ��m���?��{�C?��ڽ~��x��m2���ʙ/��\��*�l]����ҭl��0ϗ�t��>��.�#�C\uw���_ڳ�sԏ�I�2�q)�3�5r�j�U��.,R� J����Ģ�q�:�\7L(�F�-���<Ad��<�!�rK|Â��>�{�>�*�?&MV���k{s�q���%�oqF��#�<�Q��5ܢ{���`�sp��S}~��3�tK�5��;�5Qf������Yc'����
��K�+�CN�M��l}LX|��01�L�A�T�H�N�7@w�xg�R�4�����,}۴�Q�zn��i����C�nE���#�x����k���A��tdK�x(�����΁�s�Ҽb������rv,v�t����B�L��!��V^�7q�M�ͅ�s;�]g��:a��.Zj��#��S��#�:�'�Y�f�'�����i��GF]@��Q�a�kLDT\�W���#͢82��F���2-
�L��JU��\_��kaRs�~�I}��"���{��G�?�V�А���U2�o9���8p������AU�ם2�su]'�Ӓu�"�� �n��o_�1�L=Ss�d-���i'�ۗ���6����U�}�|�~6���E�*2��y��?�a�����U�x)0?�t!/�����-�Wl�N���L�HC�r�ۍF��ن��4� 7���$�(����_$�z%���f�8��#��]XN2�;�4ܕ��Ym��0�^�%-)+��;�d�u<�W��5����5Dn��쁏C���=k�<����&��A�0Aa��jՂEz��������Ԅ虰��6�y��(��<�m�kRP�h��Z��Dc�/���s�{��ފ#��~du��FN/�M��O�7���c�rWm�*�Z��~�ڜ�ש�=&��u���̇���O�PRSO���Έ�u��z����^5l��hh�����UQ����$�Xƴ�:\�' ��>�6Ks����|�e�t"Yg�
DUjT�����9&z�"o��t����ۢٵ�j���q���ڑ��x��^V�QHl�/�5��O缑�7���$�LY��k���[k�-�6;pc/y�u��y��W t`���_�|� :����1>>��^p��w�y��F���7��,1H��Qَ���}P&�&�ʍM�9n���y:�"�p��'��>D�jJ�==y̆h/RN�T�t�=@�3H��][����X��kX{�E�cώV���ӯw+>����Y:}��p4�x�UH�����'Ef�W��w�+���?Pꮽr�~�q  \�U����Hm��نj�X�9����lAW�5/S�d˒̶�^��Շ�.W�#������9% �K��|b|
NYल2]<�7�$�m�=ߖ��֩��:�Les�s���aK�Q�S�C�IӃ� OAO,�g֔&7����1�L��q�I����deZA�+�&��gr�Í��N5�}K�9=�W��OÄ�4�1a�7`tS�/��){��S�Wߧ�d�*��;��Α n�l�
����A�$5�{'�nð�0l�3��湲󙪩pUu��D�b�!�ܑ˯�J_�	��fL�F���yx� ���1��6-���_���ަ.q��d+�g��J~?<!���_W�&�L�?l�@s�?����|\G���alO�$�sFƷ?��\���!�"���2*�,�
��-�Qt�z�>,���M��f�~~��+5���n��}���%9X;T��Zv:?��XY��U;Ŧ�
�2�k�S䏫3��:�w��E����?ut+/_��jE*ұ�1I/CIG�����޶%(֏�Ҙ�]�*�Za�_9�zk��Cl�@ ��`��3|�5��a��k�<p�(��Ļ\L�ϫŢב^V{�`r��15�}���F����b`�
���!�8
N��K�q���t�>��(hvǍ�����Q�"]��vQ�#8�'[���T]����G8����(͕�}NsH���6�;�P	;��ǹcpJ����gP�GűE���NB��M�d��� ��$��抈�?񠃲�1c��%�A9��e���wl(��!���)�?6�n���>�Q��ur3L*t�Է=�/x�3Ɛ�㹜��0�:����1�~V_L�E�5���
���oM���DE)3��K�/�<�w���-�����nBf�m�V7��w�#�'�	__���;�Sb�r@̀��i���ȩ��>��[	������8 ]��{��G���QG��4��d�#���{�n}�b
~ܞ���?Z���~�؞Ci�~�p�!)��v6U�������ˢ=���<��mW)?a�3�]B��r")��ނ�#����Zb��Rʍ�+M��iq�u�q���U�P9�knK���3bʏ�V�ESI,�Z�~�{�)�᧎����7 a��>=�o�v.n�KxlЛH���ϡ�4jc$�e��2h}�\����}��W�<�F�9��L��`��M���7}ˎ�g���l��¸���p�����e�@0%6Yf�Bs2��*����YgA5ro�r��]�b���.+�w�ۢ	�����Q>I�B��|�(��cǨP�E��\;��H�SC�Ք��3�s�}����?De��a��1���� 8�I~�Ξ52����Mڥ�y��_����#j| �
u�堜��緑��u�N?�j὚�>�v�GF�Y�z�~7�|�B�)��-��褞A_����{':��Bc��9����^����q�$\G嚁�+g��٣��s��џY���	�_�dbj��~˂F"�~��������8���,v��7�0D�[H�|ga���8��WG��o�����Yon��8��6�Ā)TD����}�=>�A�f��+f�WX)�����d�fE�#�	w��1^��/co��������/!L����9�즈߷�:四>� ��#�]~}B���[Q��~U�!�֬�>o��)_��;�u�� >���ygn���qb��)��#8m���b�	#��H)���kP_���F���!L�#��\*��ys�-{�kܗ���
{&x�"��������+R����"��ur�	�ͧut��~�3��,��@ۿ��P��nO��^�xʿ/��'�������`_o��n���.1�l1��Zp6��Q�5e«����y #�ؠi���i�H��[��6�+������&8c^�^F$1
ٍ�[6uu�j]d����o${�cS������J_T�r
Ne;
���YHS���t���Q4	���Ct���|4
�Pq�ܨNKp�2��ō*�5��qC�`�Yɜfea���3�x/iE����]H��'�������%
u�oT�6�Y\���3j|��[�n+�=z�u�	��d���� ��\M�[�����>ro��P_<� qi��8��)Qf.��AH��+�T�����7,H�u�7�{�n�	���V*�m�Va~�&4�@�s�&�e����h���7߫�m"������U@Mz�,�Ԉ��Omۤ?����62�=Mݷ�}S���������1ϟ��p-{{�'�)��,5O;�a�?�Ù�_:
�΀�cU�o�h9~�D5��0���׸��ͩĖ��sz���6��WS�s�+���WE��W�{�÷�+�vp�(`�Y���aëN?aS��"�7�_0 ϏۥR�Ax��vY~���;ϡ#���)�.*#c��괵
�5���wY�:����~���.,��o^DAk�<چ�/�W�-mqe�.9n�x���i؛��1l(�Dl��[h(K+�����{<f�dܿL?������~Fǫ�����V4J-	5�����=s��/�jvGţ~;K�a��G��k�QJU�u"�&�j]4�h�͟�)CS��)�b�&=����<S���`4�RK�A��H���{��տE���v8B�Q$���WZ���I�I�B��v�3\��ԏbq��{Q����K�����e�Bf��m(�!$)̏�|ɧ��Ө�0S��ȔU��LE���M �D��"Kk�2��1y����*�L��o�#A/���c ���,ק��!a Pf^I�����w�Xc��,)��'}�e#c��q�,}���3�r}�Eu�e�o����k����o72�'�֕�骧��rr���҇�qĳO4��ZЇ�G}���:�*g0Oe�<��O���2�{�H(E;>�%��>'e�[�'MVN.�pn!{mMO���E�1��u�(�ٖ��tfS4�Ν�H�-�:v��pE��".�C��CV�x�|�>�N��n�0��?-�Q�<ҕ+�D|��k7]����@���a`ن��+9�����F�sMY*���W�|F����9L��Ar�.8WY+o������ۭ��s$1����'$�4*T����C)4��C�Y?*Sӌ2�(�gR�r���,]7s3y��?R�h�G=���!J��������ٻ/�.�u7�%���Qz-�[���\����^��J�H�cd�ysN��xw��V=y1�D��X��lGu���l;�0����ç�!�N3�n����5�����6����F�٣��p�B������(J�ɟ�qy��%I��)rոk�����C���9ݾ�-�ă���1��S����p��sG�y�����w��N������3ڿ�����(�e�޲ԥ:�|�Gs�@?�"��T	@�<0ҋ�Ҝ�f�fG(�*6E ܉��QcǸ�����*����jC�Q�M���Ӏ!z�O�1��������{�R�Y�s�cpbpf�-�e�8�mg��[�[N���q�̧;�r�_�O�
���v������h��4�SP�#@��7����Az���ҟ#p�f(���B���nu�K�/���^��������bs� e�9A7c��bȼ3"(�@0��ya�}����Lo����6��vd�j.��������ux+�-��F���1Tn���������i�M����y�� �1ڮ�\}�(��8���8P�,�&
'[��{�ή7�X�S�����jo���eM�'-�O3ܭm?i���k�����C.މ~�|ac��"��=i�$*�YuB���F�P19KR��y��C�9��y�[�����4���>��]���Oć�82m=�:1:G���חaVS%�u9pr�{'�/Ȅ@��{�?��-$�;DֈyH��wr��(ju�FL�۸�w���1�t��u�Ɔ�JǬ����,�^c�t�_����8�R�J�g�����6o��X��[��r��I�ý��6|� �Θ�=����FF��`���L{����n��{�t�@ �ٱ���W��G���(%�QJ�wF��zJoq[�"���9�}M3�s�ۋY�ԬHd�r4amw�GG~���x�~��@p��sɎ��^���+�b^���Oћ*&J<�G�ޢ\���N&��9�A�M�ɸ;�]D���+��P9=pl�	U��P�-���O�y5ҷ��y�֣(+�����o�z�:a�=:��4O(/��f���A]b�[�h��c���9���k>%�Sw�I����hor{6���7�k�H^*l���=t�)W�}sr+ ǻ��ժ�tc?���ҾG��|�)C���x����8yr�dx���#��	���%(���O���<]��6W_Ά49G���ƾ4w�]Nv��Nm~8O���u G6N���z�Q�S}E��㴭v*:f-2h�޸ܒ͎�{>hPf�� �=3��w9pX�SX0V �q@���3��M��C	jn�ʢ�K�ZP�.��,�3�#��8�8�]}<�馶,\���9�Ʊ�~�k�o{x�`]��9"��O:ԋ:��P�=�(�͹HP�C�>��7�-���2=���.Z�_A��6)�r��gUV���$�Rko0���Cs�z�MoT��3�:� ���rs�;N�B�ss'�4�R?�a�Zy���G�u1d3�B=��Ln>,e��=뜸͍�8H�����n��@ �u�����?����򕾈4��G�R�3��N�]�3��*hp����ЖO��'�'Kp��9�s��ҧS�V��u-f㯱�uM�r�7��m-z��� AӔ�j�)ճ$����E�t�9Ώ���Bˣ���9Ӝ�C�Eݕq�
���8�;ӂ�Eh��d �Q������Mܽ��<�_9%�09�iAe(�R
�`�D�6�uI�M�@�Mj]1�W�AE ��[�c�2��T����w�{����X�s��
��Bˠ���Lg�.��q����9y�sC�<�h"���]YI�:�LW�@ �	�k w=�7�[���d��p���;)�G��c�5�E�ʻ��E-����3spԡ��y�ǉ�8rث���c4,-J��qUH+���t�6���#&���aH��BE+w՘������um���]�@ ������";r�i��%`�t����<��&A���*�r�q[N�8H�̾Qʛ�d�B��(�%|�[�~C�y��7rH�@ x14u��d�<������Л����^��7f����EK�S�.缠?f�9jי98���Ũ���fEŚ,v��+T\V�GrX���`^p8�בl�����h�&$}~�+Wƙ4�2�Pɓmعy�/!.w֓�G��a�u�Ԅʛa,'��=��Wk|O��12�a���,\���1k�^� ?������I�(;-X�:E.��pMr�3V8�'�r��@��8�U.�B���F5�V�@O��N��:�g���?�&��Zƞ:�V�e�o�0Si�Յ_��ZW�b5�=�$w]ε58D��U���.���|0�;z����x��k�5.~9]�9ܨD�M��EUgߘ�7����U~@M�YY/��9�G��ߢ�3��5���8�_B����K�'K���/�e+�����g�8��	W�e�ťs���GO)� -w{����f��.��m��2qs���>���HAZR�~#7��[����gpM������������΃Sf����m\s�Ԧ���b;�����AN���N��~��Ƭ��qz��<�[����^��~��Z�i��9�ԅ(4��f�O�;<�f������Qh�h�@ x!���{�6����<�`iGs����[��GR�&�-�tږ��њ������)��/��.'f��VY�I����4��F�#\��%�?6�)E�G�/W�/�I�ޡ~�gŷ+��χ]l�b��2m�6�����</7� _���H�X���dj*���m����_����QT�G�漟�����n��"�s��ԡ����D��3@��-��A^��0��.J�8�<������y}��[���1���z�ov#F���������������Cϋ�?ﰡ�:�?�S0?5J~�%����u��j�� �gτ�v�9]�Cq����S;o����m�U6�{�H��s�ؽ��r���9��NDv�>;B���$@.'{kas^�n|�8ՂSdQ�I��5��f�#���4���mn[a�:;��U��[?s�`�
�+�(����0 N���� ��S&ټcM�gp信�q;�������nT�<&����/��s.MM>��c�� ������9@����gP�B��&y)��ĘY�;���F����Ɓ�#?�ku�G��p�}�넬����;*W|�o��H�����g-y|a.��@���B�y�I��p~}��b�
�wq�pr�.ހ\;dMg1�]9�e�&�Y����c�>��Q�|e�RJ ބ<�~�:V��S6�@8���3 ���n�ڡ�6�E	\d�Z�R��N�{d�̈�m��ǅF�x�n2o�oo�[��m�O��V�����@0)b�j�7�ɶȷ@7lĴ��A���Vݾ�]0/��p�@�ؑ^��+Tvr�;��%c~牧��%hؠ"Q�*���Y5�`$z�,�P�U���ʅ~K���^���̭���X?��&�F{׊a{5�>U�D([���V�o�@�n��>�o|��������z�	��	^�ʍ��r|���4=��ă�~YX�{}��\�:�FÎ��&��^�8�D9�U~������m������G�R�~���_3Q��]�^g���^�z�Ȇ�C�oEN�4F8�Z��)zmF3�3��p���r�د�D���ɘ߹��d���B�����9�9�(�[�9JG�97����x�ρR��B7Ӱ�3�&$\���/z+[��b������O�&�﵉!r�R��zi�ՄfjT��]7�Ƶg  ��}��S�~c��ّ�wޭ5"KI�$���A<��&��x[9��~/�N�ؓ�Ϗ��wW���iiv.�F�҆�&%�kR���A�)9+����?E���e�N��1��Y������P��H>�#��,�<��=j�qv�����<�����]�oM��ukݠu��N�t������"����`r����z̶�{T���;_�������[Ki��
ڐ��J����/y���Ӧ����!�u���CE�S8��<��x�(�)���H��+��<�J`��pf^�*�h�F�ߛ�S�9�����Y��F�~�N�.�{p��*��)��O,�F��^t�n7Ƭi4��`Yb-g��V+�<�S��j�h^���ke��6�����fq@ϝ�����pJ�p~dL�Ex(�_����롈�� ����� ��Zt6O��t�'J~M�|�������׫������ ��Ag:,���e��C ��pϧ��{*���E�&\M��u��E������p8�{h����'�q��<v�ͤ��`�����!k0r\�\�k�5E�!����+P��������Z+6����y_\�]>4-�[�|2���EI��x���6@�@09�k�C�����of��(�wO��d��R(�3��q�:���-�]�� `����	 :s�N >�ixӚ����.�:�^��"�4&����|��s~o�EG�4����c�O6�Y�,�.�`�c�|`��Ǚ�hu�����`�o{�B7=~���y��z��_5y`�	GTA��v1�F��C�L8ۿ-c�#W���q�}�~���C�w�Jt��=��joe{G}Gy�2�z����E#�7��1��&�718��C�/�s�0�dw�g2O}�J�op2�'j��L�~�x�	�7�V����d�
�HLMTG��f�jVL���r���B�l��9���\~�3W�Zg�$���9Բ�3���rt��؈��<����Zr�����F�LY3�E�>��y�LPt�R��xuQ�@0;��3�	�G�u�&��ݞ���PP�U�u�t����l�GM�k��0��;��g|��w�*>|���������؈���ix]�dW��[�C8���^Q�����kr�I����6�{��7��L���s�M{u".�L��_�<�&;p�%ޖq�:�\Cs�4�7a���8��8���}^T��
�k���i�F/��*��P񎿲#"����0}4��_��&8w�o��3_���О�����')���|.��i��Pu�K��TkH�5.ڙQa�4i�?r�G+s���F!9���U|rJ��!w�lT���SkT�r%4��(�S�7m���A3O(pGg�3�qe)S�:�[�%v��%�w�!)L+.����b��o����y����ѕ�C��_����B_���h��ql��;�����$W�>`�yʮtf'���p{$���8@1aJ݄1�!�f���nL��P�)d�^W��?�>�������F��P{�����N��g��Q��f7�����C�F�{��P:��{����g	4,�<sf���?��i�>=`�9t�ހ�l��5s���t�Q?H2�k��a���a�+2ؐ�G͞D�5Tf޽R����F2؞l{�{n>�N~�h���q���:(k����kcxM� �������<�K��.q��q_�Q���9�6�&�:����q�C�P���5���8����:�O��҃%H��@]V��J5?.�3�H�ӂ�rm��s�]�令i_O�gg�L��d_ͯS��.� d`NI\j{�S+��ue?��l��ؙ�	�����g�ې������U��N|a�!D ���U�8�n,�/��%r~�j,�+�������?�ƬvZ���-/�?坖ɡ=��_��<_J/����>X� ��ir}��(٦��+�k�vyf�e�����i]ނ�vp}<4ͻ-}� �u�l/X����ךC=z�j�3�#�aO�GOSt�6���q���w]����U̴+G�eo�Sn6��@sNw�G���3	G��FzY�Z�V;��W�3H�F�"pD��_�(GW��hc�QlWqJK���4��l^����E��H�zpeM���^U	�`
B,�'�[���>������G$���u�y�X��Y~2��ܥ�.�d�O�7�?��B�^� R���;U�xƲC��2?��$��ݢ�<cP����8J�����#�kX�ˍ�7}�] ~�YB�1Д�)����<�9�J����Cq����n�5�v��o̦W�u��u68S~kY%����_gW=S���~�-�N�qd�r]���0�.�눴~��އT����	�s���sx������.3l|�<��0�"�#������x����>I2��2�7�<D� �D'@��TVVKc�@ ��~)ObO���C�B�.��:!p�>�t+9�ĝ
�J��tOS����Ǫ0���o���T�
�`~U�ڠE�`T.�c��$�T���A���}z� �"^:�P<<�7�G���;���z�>j��Edy;J�f0J�!�Z�oit�pJ/B��������+��H����1��8ku���fD'�8�`#D�t��v������Fg�������6J��NY��Lq�	�@ |���@��'K@��y��c��:�u�8Ѧ����p���U9�Y⻰�d��b{>3"rF��tRKk��q�,�sRml}�Z�Ҝ��?�A��E�@ �8v>5�O��F���3��WlohG.�g3��ܶ�B��\��yw �3����L��J]~Q���������UPf����M�f9"v�����\��'jjt�o۠K�s@8�kC�aa��XGȅ��6��#�8�pg�� �Ƴ��IӮ�ȴ�35:�k�����2�)�È�0�&��@ |��g'���i�ϻ���+T�:x"68Bc^�m�`�!���T�QG�p��M|9�N�T�k�'���q�0�����#}��?�qm/�>�I��� N?�h'	�3Wˑ��}�_}6}�QhV��XW9����=mgN�*Z6�{�<��r�.fFi��ɺ�%�ڣ>�@`�6�+�������@ x@����v����ǂ�jы�-�c �|~�k��Qy��4*K��2r[����<�e|e�flÐ��F�AOt��<q~��2%�l�,<��e�*б���ƷρCk��8Ø�oM�x���8���?�];&ls�X.a���y��Ý���oqJ�P�T�2�\^o�?%�O� cA��=�m�~�b����;��Q��#A�ڟ�!�0-�����Њ'�'���Z�Ye�i�o�%k0��Q"L���I'�`�JlQ�)�X�r����A�o-��w����ѻj��g�"&bC���֑s�/E�8䉱�I�%�>Ǜ�Bq�3�K��7C�?�;'�6P�=}v���Q�{�v��YҊ�Zh'��>P,�я��m��@ ��^v�����ƒ[_ksr���xW�V\����s��sߔ���=�:�+���3C9ǅ\��r���� w�x�|���a�������9�r
t&��8��;�u��9p�B���`�vޒ�s�K�"xdL;�ֵ_#�7�j�)�O8�5|z`��ik�x��,�iY�ޣB�^�@ �Dzj��^�`�JS��o�s�LQ�'Wv���(&�6��Uȶ�<�@09g#�V����"�[k���3�Ę����5�P�cTT �]P�QmN�42Ӡu,����[�3%\}���2N��Wt���{�P=D�Xw9p�,֍'�>	��H6 �aL��n�NP�̏:Dk�y^��!��]�4���p, �~0A��F�����&b:zz�pB{�Y85<�Y��@@���>ғr���j�H���+$2�7��Oz�W0�<�����gyң�h��T�S��qu0�5�"J2J��E.�>w����sy*�J�=t����@0%r;t���CQ:Ǆ_��r���Zx�@�$ު_�f�P���혥��8��_�1;���x�������н���1|g	ѨE��M��_�3�]G�$�a�iw.L�1��_��\�Ծ��(;q�j�>G�BV��~r��.���@�5��-"�0������?ݐ���TpL����{�5�=0��}��4���v��H�x;�H��ǥ�!:��b���ߕ�U���=Х��J*�I[Ո#^���A�c��ڦ��י����)�@׾�,�8O�7��~1��� v0ޖ�Ϸ�&��R[���%�����5�?eό3�գ��e�}cӤ"Wq��퀭�=�A ���V'2�T#�!��.���DQY`Z����yG�>zJ��U�X�6�Y�F�K/���Ȁ�FV=�V���(��B�Q3���U0�/_�i�]II�̻�8��7!��i��Vz��W �7UV9R�&N�)�{Ӝ��+c��lz��տ�Ռ�,��q3��:0<X�u�%�0�1e���<������p��,��vȡpݭ���h�a;��[���ED�=��a��h���7�O�.M����[\۴~��ON;m�0>�Ӌ�w���_S�3*��)�WT/9�l�ڮЁ��(���
nW�R��A��.?�Tc}W|#t47�ǐB�~���5C��Kuΰ��Hx'�+��I�l�+�m�F��>���F�#�gk�78X��n>b`���JOqY�%� ��������i%��
"�9ީu�6z��Ι����؀����sǭ��H�4�+tF^ �{���P[��95���<p.�#g���\�VY��@�U������w�anr�)��'�,(�wi����9]�F�e
l��<�>è`�n�z���1�Ӗ����+���/���J�F���g�p�M��(1Z�ؐs'�Ju�id~� ���39�؛{��Yg&�����6�-G�[gl� ˑ��� ���@ |M�>��*,�
4���/�\��7`���"�A�|��Q�s���iis��2��w��?D+�A��3m�ܣ2�����ǻp�CVk^����tb�5��$�	�;�עECu�)`/�⍌��mi��g�G�}g;�]����������=��w�y~9Oy{�cQF�Q�b�C��tc�5�������Oݸ�^Ϸ���N3�y)��sw.����vξ�	�C�7z�^q��iԝZk���?>.��/g���jId�Rh���Y &��wD�/�8b��8q�� d ��N��Y=}�w��'�@ ���E�hnݧ��#py]��Yo>l;�i��!�I���H7,Q4Ϣ=�ڣ}*��Ȳ�<��뢩��
g�A�Zf�O}wP)��E�wg��W��L��	B�p����_W q�y�T���糁,��?�|}�}�.g��81�~�@ � ��y���>�5�W����M]/������8?��>�?�0��6��[��@p%ZB������_s���(I�@ ��
�E�3TJ���l�Q�s襑�&{A�/˶g�1!w�  ��IDAT�lj�����=;����] �y�^3}N��D�r�����U|_Z��������>�;�O��ՙ��[o��\5�|	#��7�3\)�<wE��?����ӓ��V�����&P*{a c.�}���W&<YG�3����iZ8l�@��z^��0�re򟳠�贄3z���l����Z))���ަ��W��Z޵�gk����^�7#�q$\��W��lm��>G��v��ᄹ=cul�?�iS>��5C+�{�G ��H�fй)A��m�mT�ϥa�`��F�tUJ��O]�!�G�sx	o_{u���C���s�0�ϦC ���DD.Ft݀M���J>������4�-��:��-�w��{u�����a&V�be��z�X�-����k�	�n��XcO!#�1\�w6M�Uc��s8�w��X)_��O��(`�s�3����`P��_�w�������Ԯ��a]�2O�r��8�xڧ�sQkd��4�C8��Fj���ʇ��#p��l��������O�/�>�����{��%�Ǘ��ZTx,�b�J /�"Z/nc����oc^���/�m����_.k�,3��G�b�ou�.ፎ�o���1'�P>�vlۻ}�A�5��p�PS��ߛ�kT�+G�s$]�$�B�)�e�uF�����,���=U�M��z"��p�;v܍��i�ܣ����Ǖ5�!��}b̏-h�ZT��Ր�'��~�qc�J� �&b6v$E�*��k@ ��M�J��r!|��q�Q��3�ZzV����=���2�/��{����k<��yQ�Z����A7?�rf_D��(>��}�cg	�'`D����t�#_8��.��og4�*�Cf�k��{�;���'���_,S�x�̀�8W̱�}n&&�z�4ܳ��ue��1��S��f�wпZ�xst�*TL���	 痣��g�ۯ�4��^�����$0���G�]u�C�7狜���i��?��{kxXZ�p�'y���?��Ȉ_��Ku��2�@ �{h{W���"���"N"���1���B#5�(S�c��d5h��?�8��Ufͳ���{�O�E������g�n��(��{Q/��h�HN�1y?�����ot~��Ԁ#^9�/��f�C~Q<��ǔ^$VB�n�K�=��RR?mi��{��h�d���u#ʻƬ�C�B�8h�&{�r�FR�ֻ@ �}/���z�S:C�լ���ͽL��3d��AΛ�`i��G�(�v��+P8~GUx�u��k��ɕW��"f�+Z�5r����\�+�˛��L$z�^<���w#R�@ ���=��6l��w;M�ȶ�7y�j��c���`ZE\�=�#j�����j˿
�]f���;�����F��m
#������X�2�7ήdnos�m�#6oMe6��s��^��{��J�9]�`Ĺ�6������*#9�3�"w�%"��eN�z�ލ���}��-��D�su�!��U�y�C����PJ!�k�>����#p��2U�Y:�O%��5	�#���h�C=���?��B��N][�y��g!�@ h��}�ь�t7hp��;�q�&��չ����芉Tj��or�?��^\��ؾ����яu7�հ������Vl��U0��D_��,8@[k�rHI!�#��O� ��-swĸ�5��Y̮��lP�R�r���ˢz�Sp|�9�`�s2��K{������I9otw���a�OF����=�S�
��	�{=�����E4.�(ݼ�N6a|��n3`�鱱q��]��YOېfGI??�G�|��s�b	G����X�ּ��	��p�ȧ�]��ʂL;@o6�cwn�y�������8g�������i�2��vQ��|G�ѻ��w�g9S%���U�[��Q=��6�|���*Ӯ��|9g4=A��;e���ґA��ꔐ�k����[v�u?	jX���#�Я�8ju�n���p��#J�f��*/']U��S��p�<j�ߩ"�t�-	Ϟ��p� C�Z�@ �.��#�p�[\��2ܹ��F�$�$w^��fq�8������ow��e�w"�	��k���K�x��m��r#a�,���q|�G0'ΞdzZ�iA;L,.��>���u�Z�l��q����u��'�����[[�wkE�%�wv��l�w�F ��N���;���	��@��0�7��Ǻ���m�>��L����@p~���ߜk�ݭh�7�Xҏ��pt�FM�!n���l�}�JMY9�\HVA���Py���0�$������}��oc��ҙq�|c���Sǐ�O�~���2�8��aC<��O�c�E�������������;;�k%}-?���#��2�Ͽ���1x6c��/�O\S#����5�5��|��,�~,:8�*�h���3��;ḱѹ�!��s>Bn��}ɝw���q7ww��`�ј��� ����oa���� ��R\��
���Q9gUK`m��6�7u��
���-|�s��k�m�@ ��I�gα�M���9JE�me�^���2J�L��]#�lm��a�-|��9R�L���}=�z`~���N�V�������MO�<��_������s��#}���";�;|z<�_Ԗ�e>�:4��/`�v���Ls�;�}��2�üh^�m���	%�<T�����f��_�������~7�����k���;�j��֯Z`��-�W����� ��[H��c"AH�w��2�g��a-�������$뚬��[���%��N��

�,{��
t�KD�us�������%DĻ{I+����vɹ�Jސ�[�sv6^������C�m�C*O�;.{&t�{��q�V�٘Q�zc"�������(?p�{9P�g��R�ȗA84�*t����c�梤�/jpH�g��eY�9��)�6���52u
�=��8�^�:h��;ui�8^0�c�.����A?��fa
���p����xz~�S�|�;�f����PdWx"�u���o��{�D ��=�ܳ����U�\���U<�H\��L|ٗdů*�FB���S0�]��?3�⨽�@�
}��] p��;�CG��euz����ڗ���'�\_�t�o;|9s[�Fǃ���z�>���+� �k���< -�5�Gu5>̱:+�N�H�߃��o�|m"b ���75GV���> ������9�[<=y����������,�шé��P5�N��xY�s �ʘxw����s[ x-Jqxo���S�@ �{|L�g�{Q��Z�@p'f�������r� �}]�Z�SӣF��'�S�LLH[&<���ӐGOߌ�|�WI1I����
b|�y�aq�W�q|Wz�G���屾��u�?�2�dK��Z�q�:�kT�#�OQ_/��g�@ ����N-�������	8<�0h��RT���B�$�(�L����q4���~	=ОԔ����N#�gO�d��_>��UU*§ף��	�"��9{�S��O�+ǧd;�eN̶^zP%O�����}�W�D�]j��'V \n�^����Y��4�L��>M����p0��Uw7�GQ��>��Ֆ�ˢ�_zFcX*��]��s��O���+�W���{WCX����:�����t��q�#�.��G�:�_��X��\
L#UXg�/������+��r3����p���y��s*�|7���;���\�#I��g܇n>������<si4�Dy$�p$OGY��g�f'K��Yi<� �99�%9��M��s �5}q��Ho���b	���5Vic��h�'�N%6�_�cӮ�[�Xl�AG�X�,�!�MH�q���J�]������Ҹ/ωC�`�A*@O���!�/�yr�<�.���㡱쉟����֓s6���amN��~��P;�9���<f\�����[tM��+��#N����[�(�	O+е��Ӎv����ZզN����?&�p�v^���9���qb��%W��%�5���(�7WV/8�++��)�km��(�w��������(W��|!��80v�x�Eϵd��H�zS�Ц�`�:��y��D�VqE �ë7�?�ʵ؁N�?n��N�`�e��!Gu�<�F^��:�
�'�J�7!�0�mG�7�ɓ9��\���ct�w����h�i��)�@ ��~Ͷrͺ��:��Qyq:F/Oh��|�X\�2֙<8��<�F��2#��s|: ;��6W�ݣ����v\�Q��VY����[l<g����7[�SI����p47�Us��:|�������2�8v��s>��t�-�<�J(� ��x�,�Q��ec�y�῭�=�x��g��7��7����3�������s�) mCN�V9��i��P�cW�(p�h��Q�7��Mp�����W�~z�?��	��k�T`��S�Ț�Ǽ}�����dF$s
��w���|˧�@~����m�zy���˳�;x�Y������i��j�<h��7�Mp��m�O(��}86O�m��1m�n=QB�϶hg���8����_�G���B�!\i���B=9C=�:`\<.�،��ur�LkYNo���=Lʜ�-oA���~���T�^<���#���A�)�_#�܁7�?��(vR�h�Z��D ��S����Y�*>!�9�t�~�����=��G��?WG.�CM��44�R�Z~�E�x;�d��ը�+�6d1AD�����a)�N���ē�FPe׬�۠�x��7n�<��˱��Y�5���� ����R���%0�'��NS[����>[�s�P�����'��@ ���=�C�:[��#�0.�Ke�7������ig���	o
;|Uf��(hLl�,u2S��D������qY�"p|X���;�����+xD.��<��Ps%��o\=s�;Z�����|g�Hۈ��+�G���M.�Q�gu���!�z ;9�� �CX���қt^�<>�&}8��p�xQ� F�V�-#8�n8���/!G�K�J�J�� ���%|e�k�n�q㞟&�nl�>�C�g
sm�4�G�����2 pm���;r�IQ
�D�Z����@0�(�Y w�J��8��Vm�o������?0~�v��ڏ��$�:��)4Z�w�No�i?.<�]u/�w�cN��$�h3�^z�Z#?���)���M崫�:n_7��_G��9���Uw��g�i��1�d�i�N/c'�˰�hL��]�C;�x�~!����\�5��?t�W8�7��a=��l+4?�M(��9��k��RY8ͺ�I�w�r�<r|)�-礂(p��D��1���Ҿ��Jr(ԉ�x~���>�ܼހǣ��� p������[��ͩA�������a��
Y')�G��F�Y@������̙A�.zp�|�F�[Z�h�EL>JD���q�ϣ����\���M(>�M��\c��W�*BM���
Y:�-=�^�l�$yX���Ԃ�y{X����1�y\ݗ��d��#�N}E���ƃ��.F@<��`:xZ�����k��\s͛�\��������j���_�����N$GN%9��}V�H"hǷ��-q��R������r�؃nh��NS@?E�tv���6]c��iE�8�ů��U�bþI���ت<�V����x|��͝��E�D9���b6�S`�gp�Z�e��k��W��A����;ͭo6ˉ#�@ ����&7���q�(��hvd<�C������
4Jpd�/�>�={A��`8�~�<�?��8���_��u'zy��"��\�H����� ���8�B��v�'�4���">zV�����s�4�x���=��W��j�>����c�Ym�������2{�U��^�H��=�sr��J����?Ӷ���h����g�1����)����sz���*<	��0��
b�h_�yGZ ��tZ��˽8��bR�ȫ����$��1�4}-�P&r2ә�K�圧k�̈́Y���8��/}���
#�ELK�
��@����K7 �D-߃�k�H�sb�w�|�AOd�� *���fR�7�Ö�/�O��]�s8W����y��
��D�8��}8H��
�KC�O%��V�P����ɞ�~�".M���jh��M GLk�R5�ؒ���(1�.�Rņ�r[A�D��0nG�r�ƿ��\:�,�/G�hW�3�ˑ�K�{�
D�ц����{��(͡YQ��c�A�dɘ#)!�E��3��Ƕjl�3
|C�����5����/h#f��}�@�Ex���-ۃ[6!���!nmX��e���ˮJV�_����~ߤ�>�pi�6��[^p�0�ߛ;�|08^|_�+;R��~�=�%���G2o�\8���#�����(�Rߗ��Z�}�����>H�D����-*Ю�%q�'y'�������2�^Pm�@0`��O�����
)�06]բ����ns��M?,�<�Ҫ{�Y�]���@s<�dq��̓ʏ��E�,���gAH������)��]V�)>��D�Ɔ�Ӭs�:�o{�fYU��wQΫ�h�ʴ}8���������
C�g0k3N ��K�e��Q� F)��T<�:��J�9"�K���HE&.���-s�cN+rs���Jk���j�j�����l:�z9��2fD��ռ�j��(��m���_��F�9N)S?�w>'K����gs��@ �Xzc�3dgL��Ky�JX��
�ݽKMuX�	~���ͯ����9��:w���|�8R̞�gē��#���2/gT�1� UE�?s�`�	j�0�a	�qQ9���K�x���\��j���t�|'�YxE�9g�ZG�v�」�-9􂓥j��s���s��(��k#���;G�/�	���w�1h����Qs�����џ�PK�~��خ4��J�+�ZuF�0ޝo��N@�����+��s���q�m5^�@9��:�(���`DPĘr���ո��(�9���F���5�hq��S�@�t'"�%x<W�P>��.ʮƟ�/|�JS�Z�� �=T����@ �GP��B�	�G�0�TD h������~�ǐ��z�B��.��z�>`���Й�/@�&D��n��/���.K�%�޿æt���-<j��\ږ�z�]�a�v��L���<f�k3ȫW:���|T+��!xjp��Ĵn�=fJ.�0xg ���c���y��Q����g ��#r��{���"9���#$i��a�{:i�h����Vs���sl ��Q��!"=�>|�;	���Q �����H�-ʣ+AO��S}��rt�U���lz�a�@�Vc.Qy^b�����\	酌��0`_����Q���f���ȥ���;�G�d�����lc4�BE��jЩ�
�.���}�'�\�\#e½�=�����x����Fe��%�܏{��^^�u{�;��=Lǈ
(tM��Z[,f��o���զ��#�@ �:fT���d#ց<{���|��e�R0� ��FxX���uf^ #`�x�R��$�U�r�X)�F+�i=�:���F��:�/D��\Գ'W�9$/D��j�}�Js�Мm�����M��l��S��ۜ7f�Cs��h W��Q]� b��E[G�G�\���f̽VT�8���xv�"p�C��U.�ټ-�N1�8�$�(E�ȁ�����K����xz=���u��ǉ݉��z���'��OH/VY�O^����=s�xH}�@�[0�O�Ȭ�e)�1�ڰZ�(��(�_��Kr�~����泡�'?:�uϽ�:+��߫�ꍒ�{䲷#׾�yE�5#��ΗM1���C,�<.�p�Y|{�
�����S�����В�����A�\�܃�����e#yq���s$�ն]��\�Ým�9�ɳ%�i�So#,iԑ)�]W�D:S=sϵF��&r8�'_>p��T�'wu���s�ɽw��c/el��ְW&��������u�� 2G���c�֭���u�Q8�<{��=�56��_T�@ x=���;��ٻ5�/������1J
?��(��|Sh�_~T���u���e	�@�%T�u�`
���9���������u�\�D��'x?>�`#ӶՁԎ�n%��V�SL����.�"z�G���7\8"���:H��i����i|��:r�  �ݠ=c�;�&L�l���W�n/�yCu7�7A>���@ x��+�Ow����d���s+���!���"pht�s0H	y~-�����Ui�#�2.1��-_U�QT�p�½*�ޯ�ÌA߄�D��-j�wj���*���~{����錣'΄��d(�TxOk���"����O�����%�l={���8�b�u2�kk~�|�����2�f	�;p���.���]�e���r�g�3�|�5��k������U[F�x����]�J�\��s=�/b6�g��^w�Ǭ!��a�oF��۰�o!��ن��ɳ���b2?1�t#1F��W��mM_sij���8r��*'�4�������s�ݳ���~K����gW)��8r1���>�rP
�D�p�z��e�+o�����3�t�N�s����4o	��,|bN����9ߝ��~�_>��a�Q86z���l�߅���9�@ �A�CC4��Cz��镟rih���.�����˹��5m��h�!bE�AMɑ�����D@�0�W�v��48m�i��D�x�"D�c-�>s�Jfɡ/���E��gzx�'�Ս� je�\>WֹF6����U�]opd�j�	�:g��M3V����<D.,��53�Ɂc��1��y1O����Z�讱p]�:�.t�h�=Ӯ@p
�� �Yڿ+p����1���%
�������HS|=����4h�����G�wf�6#�Zs�
��K>3)j�l;}�f��y�23·��y�����'t��zт��eYN��³�:5h�s�I�V�zݼk��@�`x�T�����կ�r��i��h��>�!)-��f��.�ņ��_�Ao;����������m�����I��o�����1'�����5�J_�/�q��W��b�ƚR��P��:��g��G�/��Y�S����g�J]Uy5q������]
�äآ�w�^me
�@��Q���a��\�\ފ�!�Dc�-D�DRW�cI�GIYS(.���b�ͳδ�lİ� κ���-+ـ�]�Q
�B1�� �g�AZo���y�{P� ��w��yG�[���Kq��x�<De-
�B�xr�gE�k/�{��b]�7c�}��x���ἳ}������V;�ۀc�����V4s�M�B���P�q����[S���E��u�b��.�#�<3*��&�0���%����/��a�9�KC�<�*
��ឱ���'֟`뚿}5ѓ`�в/�J��%�H���DHh-'w�Y^�_�Qʷ���I�KL����8io�P(���n�a�ӹ�e\ |���V�P(�	Χ���B^虌 T����6��Q@�F�woN"W�rRK����	��!	�T����l�P2���kw��=�3K�4��#I�Wk�Q��2F�]m0� t#iQ�W^C�.��%V(����<���<&wMW��y*��f��uYM沭�@�*5v�ěq�3�0�f �[�t�H-����%׵9#Z/^���韀��u���8Z7����&���*
�g��>�@e���Q(ވ;� ���]Y��Jq���6
Wˠm�s�� ���MKOtp�
.`������e(�p�<T���?A
����3�l��;����ou���Y"�_7o�s�/nK�s3�s<uƓJ��>%��k�+�(�6KW���B+���_�6��U0���S(��y8P��?6�i����WQ��˸��h�<p�S�e+ט�dq�P��+��O�uTY������]��7���b��3���V)
��΋���m��Q��j��}����� �n��۸��D�8~���{@�%F�[7-��l�������xΕ�zH�m�ܾր���a�����16��-W�d�4�Z��j�#�^7��
��fx��3����7�����9f1�Z������y�B`��U
�B1!R��p������a��`����Y���g��t�+��v�)�_G����:qמ���is?%,9��mp�rge�z���(�Ӈ7^�� .H�m�6� �_~E���9nW� �/@�7�-�.�O�^���%Ѝ������#y��f.a������9�枆c.�Ւ�	�؊�����͉B�P<�$��a�s9��z�P�"�Z�i�ʳ�]�
�G*�_��B���V'ǋ8��O�QJ_݋)�w�]� �4�wp8�`�w�L��8�M���{ -�����t�p�:O�<�D�5ri��&Cg��\9o_�7��}�����J$��E�t�cd
�ۛ��xu��ڮs�ҳG�B�P�ūL����ᴾ���&��*���o�G�U&WO
^Ai�q�C�]���
r<�7N����X�W㷤�
��ӘW6y�iݯPq���� ���3㺤�Q(m��_����:��^�@mβ��s����̲uBH�f��Y���`�w��ڒ����q��Q��BF{k�;�O
Q��&wW}��'E7&�1xj��ܦ���4������?��h���]����p��1�+���L0���o1�m곋����͝�����B?d��%�c�����D�_gC�B1�?
��*RP��a�`���u y�5����a[����wn��}��{���Rgi_״�����'@��S~�1~����6),g,��Y�s��N���s�,�o2*�$r�o	)�� ��Y>ܒ�m���_ɀ_�V�B1
��:l���h�dYh�>
6�by��ά��_2t�a��l�\�0�^� �y�����K��ГຯG�M�h��d����>j#�ۀ��̈́�²�	Ԯ����g��_����3�6�t{:rd�������&��;,7�@�)��?{���X�i<�B%d��W���&�[�Y����s_�a���YB�k4��ʻ@O���H���8F�P(��h2�U*�~:�0�����3�kL0Dw���=�HJ�I�V�x�;�o�д�u�øZ���)�y�h��{_�����}�,�Ó!�� w�05�u��k�
D���[k��Q(o����}m���M����oӫ���eg��܏κY��Y��?ۻ餁p��[���7���K�pLO��hsF�����q���sO�Ǘ0�r�ǆ �Jy��F�WY���K�1qT�K+�^�3G|�8��V�����J�G8��m;��g��lֶI��pe9ɋ{�i�y��(�a��6-s�7Gf *��4G'{�
Z�0г:�v؄~�_b�(
�Mp�}�;�ם�!{��-��FS�q3�,w�ߒ�8
���KU4�Z!�B�P���$��V����m�0�է��Iz0=�;78o���u�g�����Ne�o��.�����%^��	���������W�$;�d�\�".en����U(ނY�K��wX�Ύ�����m�����xZ �����+���d�z�P(��q��t�3����	�$�h�׿�-�
�B�C��)
�⡈���oM�<|*��BW�f��A�Q�+d��F�<p|Z؇��A|���U�)�}�;���L�^<�A
�Y�76�\M�goG�]H��:�c��3r��&��4t7�+�G���}�}�����
�����������)�
��쁃,�_�D�Ն���Ue�eHWh��{#��}��V ]f�ՄU�fR(O�����B('E[���X]'GE3�Zhj��_�Қ�,x�-e�I��j��y_)�WxN�|u����p����=0���N����&P��]u�w�,�n�bJ3��ߒ�=p���=�-kW	���c'���-/d���n1������_\Ws�)Q(��"�qLg�s9Yj�k��9j��o���9N#���h�f%)o�������7�k��V�>����	!��g�����y�Q��C�ބ�Xj=i&��������IyF�����(
�X$W ��GhW��QxU�x�:�:�_X� ]�R۳��%�ͣD��1���^�9]9ވ�S���c��ךO.~������/�)�#�R��_�>�a��y�4���?�W��'T��h�<	��,��%\-�ۀc5kZ(��z��^N��N�<�%哱s��YZ
�g1�u�'���ކrOg4��Mτ��9Z��S��,S
�B1!�q;ow^�	��'��<��!�����#r
��n�y^�X�i+)�?������<oʣ�(���x�M��xZ��co��m�`Pi��`
��\]�n4{��:(�O��:?*r�x����N�}or�u���-�hͧ���m��kIa��(�S�G/zx�Z]�������dx�E���#���.��hIOE���������}BX��ee������{�*�[/(*R�%�S(ގ�f"g��sH�Éh�B��N�|*
��7����0��+��]�⹐�����������pG�����nP��pr�_]���S(�A�@���ہ���3�[PPt��j�����1���,+��Gi_-�;c�}Š����:��9`�4<�1by���u��x�b�Z�@����c���zK���RNz�iZ t�(�{�;�줵E^g�?�G"҄��Ne,̟�*>U(
gȰ{���	��@�"�05�1�W�I+���ɯ<a<-.����Da.��:��
���?���F����m�\�(zS���)�	!3f��{�^���ֽ���wx���4�����zwp��-Tƿc0;�+E^�J��~�O`�#9w��B�hG�b��>�7#��m����:Ѕ[v�4�Y��=����ڜ��TǷ}?̣�Q�X�P�v��՝���2���,�ݻ;��~z_WֿuEZ�;C~ �r������l�����>H.�K�CP{��5�}J�ۻ�8(/7:�*
E	�ٿ�Z"�^86攲� t�o�U�����c8�W��Y6>/=�[U�z'Xy}Υ��}��R�3���=�w���	u`<����rG�1|��������ͯ�xZ��縯�HQ|n�f����G,z�%:��}�fmR�M:��O�B�\H3�tG�8�E��l�!�8�cq�8�፩��'+�v�V ��O�'����>�iU(���4Tc�r�݄�1N�`�ӻ�@7�䡢���F�(��
e�wI�+�t�j�~�W��� z��w�R��
EX��4c�rF�g�
���kv���|��� �\-�������)/ 2N��c��8�N\I������+���(c�Q8COˁ�;̿�}��3&ߨ;"J�6�׀��� ��~!��]�P<�bcu�#i��%�pm
�XpYx��X4��n�t0]�����2�P(~�Y���>ܜ��w�Ԇ?Fq��?�vw޼�R�R�'+#�f��%�B�P(�p�|�q�A%���P2.�\�7n���B��|��p�۫�5+�_M��翷��BI��Ө K�xJ�v~eq>(b�u%C�[����WG��P�|_�?uM�R(
ųpv��F�>�`%8vo���*�P܌;��(���?6�Q(
�l���3*�����o�+ҽI��5q�5
�������ܪ��Q�Bee'�7<���� �u���	@�Bя��YoG��=د-Y8C�I�qD�����_DfM88݉=��N\/F�d�B���p�:����j<-��-�oc�ĈBӪ�����ʹ)��~#�hx�@�1��
�b|hN�b`�NA9Ϸ�#�շ./�p�q/�^/>޾�+i����*Z7�ɕ�Z�d$4C��x�����e��FR:���큃�q�n���D�y#�K�/�B1gջ���쏾�ѵ`�LDt�1� ��A6��(�Ub�iO����P(~Λ�fǞ[�bf�$xK
6xpj�	k;5 �D���>��^�eӌ���O�hw��Z�)����B�X���O�af.н��-�
�B1 o���5�A��eovq�n�� ��4�$Z��<��ޔ^�C�d�h���	��_mU�o"¡��>ô�{�RZ>���i��0����㉖2Z��۵��Z;��s�W(M�6��|O�ܪ`�x�������Z-z|*D������ �/E�p���8(�����_P�X
�u�b0��t��F0QvE8�
bM=� �W���y�S(
E?<�
���+!�0��p��P���'��.��lD9���~M��d�W(
���a�H��>���+��̎�1{�A�~����z�h���@oٳ��Hz��?��_�w)�+Gkzh��yޙ6�b�f��t�\��#�h��M~R}Fr��b(�CΚ4��p���<���x:�+Ɓ�y�+%k�3��7�����O�)K�B�P�,�Sc�hD~f��20g�B�P(
�B��,6NdSXS��� ��S��q2L�Q�n�_3�YOPC`Ť���Yж`vpl�b ��9+�%N��	<���7�j8�P�Ar=��x�~�K,�i;w�I��u���P���,NůPqf"�Ի
�B�@�͎� �a�I��������+T�_�sީ�V(
�Ga��ǳQ۲���hD~O��\�ǐ�˿�5�<槯ϕ'y:<K�ȫ4z���L��\^��K���c������[)��l����<Yn�}��?C�+��s�W4[����?�;EңW|��x�D�x,�8�Jw�a8^ou��<3������[('��B�fx�X�������ۋ��Ib����D���R( ��OX�pHY'��F�V��}_�n��D���[u|�
���^X�Ɇ@�q�ށ�>*�~w����q��D(�P(S!��<IɄ+�F󲯡�׿����Z�ӹ���5ȭ٫y:�"�?��H�`ZTT�m�p��w'r�,=F�9:K�5O�b��@���i��s��\�y��B���x�\:i������_˘�y�=�y2�������g^�eͶ�,�h����"�אp��th;��m�2��Ig�<*�g��:>5w�B�=\�S��4���:�y-�˄y=���6Fӌ# =p�͵��PVg��W�Nq߇2
�� ��zs�"^�qd�y=xm*͸n-�wL�������F1��R(���g;5x8+�����B�~�ֻ&n1������H�P(΀L����yΰ|5xm�1�õkr��ɦ8�E����L^��.���aj�������=*y��y&�ϤtܸA���t�?�(]�*���gK=����Eˡ홣IBk?p:Ό���j�1�D���z����l㬔n���2$j9���΂������m���u���z�L�ap>�n=p��Н5.mN�;q�������o����~ m8���*��ǚ��n8���e@%H��=�#G�P<	��{tg�a��3���ǂ�՝0�Y�u�}���ʗ�G�	�O�!�v����o]
�b���Y�V��hTp鷠�x��3��r��IO���[���Ǜ�E�X���O����j�h:)�eYĸR�\-�>K�7�Xٹ2sm[+��7�����;H}*A2�y>���>q���Ēzã���]R�}y���r���~�*V(n������G�oa����3z��,�	6c����<n�$x2��t�wK<���mV�P(������%O���?_��P(
�B�P(>�Ԩ>bd���,�� F�h$e���x��R�r^)�|r��[��}��/a���$��o����@�=#�S�吠ۀc�,��&���[�,�p�R[C�eR����?9�6+�[��
�bG�C�b��8,�ֆ{9\�l�`���K>�)�G3��I���9�oZjX�y0
�B��nM�Nkr�ޘ����Gz�p�)�B�P(~ �WT(
��<�#�%��+��`w.Y�P~K��935d���WlH�P��UM~�i�e<�T�)�j��e��O7ȁ��^U33��8�.�94���lyU'�n�ůΡ�Ɵ~R�S�u?�]p��E�z�P(��^K�	�ߍ鞊dA�ud�J�W��Dȟ���9
De\�6��E�P(�	�7iZ�F|���#'aOq��eN�=�X�[V�R��!	����/�ρkj�=��OG���P(��H�˭�B�[�辂�I�kM>�/|ғ�h��򠟹t��FJ��g��ɕU��v�J)���r�=j8�lY4��u��A�x��U5#���!��ۢ�s��[y��Wُ1��v����o��z,��k�c2���osu�w�?������|aU��P�CMxO�2z�.t*p�Fz��\=�����vr�L���n�)
���M㟎�\u���!�"/��Q(
�B�P|�t��s����po�����
������8ϴ)Ig��eT���V��G�=��Z���I�ٟ C؍���`,u]�������Y*;W�7z�X�{�'�7,~�pJ�}�
��l�J��e>j��A�ק(�q�q�Ǹ��"<e��Gv��c��Ӹ�X�"�#�{�*���XV �A�~}Kf*��T�V�P(��ɞ��痕�A���������i�g
�B�P(��Ҍ�mE����M;�^�5ܩ��
��Bx6�xF�]�G��(�g�^��'��1�|r�Z��n;@��tR]���+T�o�4��w����;�:�����/�h�R��W!Y:��D/��j�r����N�5�_F4��u�Y�vK�0�W��o�i}�(R(�q��.�[�&4�^���צ_ǯ)��k�,PU(�C��W}W
�B1��װ�5jpm<ʿ�!h����`,�=���m�[��#h�����~	\N��w��'��<��^;�=p�p��7����Ud�㿩���[�vK§�F?ne�-�l��$��[&f�w!�o�y.~�;)	�1��jg��R���w'��$���+ 2���E욓m���{,,E��*y��1
��9x�>ׄ��of+�3������24�X��0�Vc�kl���@�g]���*�[�7w�t��|�L�@�6k�/<}*�
�B�@�N��nŘK�+��vf�i�84�a�q�ڑ!{�_&�Ps�:={���wkU�3+r<o����c\g���MF����:��6��k�
�>�-�p��(vι3�U�G�f��rvc'|��(�ʩށܤ�i!�''���й6�N4r�_���#ǧ��d�)�2;{g`��«<p��x��l���qN2�|2���]�y�z)|�}���n�tvT(�D!��	4�V�:��1Q�f�}�g����|?����,�Q����X��	.^�6g����������+�?�W*
��������̶��|7� ^��}#�����7�7�!s
�3;��0�Q��Z�T�g��Nt��с^�K$��%�ַw�x����Pl��Ovv���i��خg��y������G���0z�_Jni���7�t"Mڴ�ɵ���ⓐ��6��������(8=\=B�]�hvh��8��h7�L�/+��ǖ�� ���_9�Q(
œpb�o���e�:�bF����@�P�Q�Uf�tS(
���*�{��e$pCO�7n�t��m��x�xx���pG��vE�Ytpx[��;X�d����oT���z�t���@7�~5��\�:�)�{ո��՛���,k5_���muAo�(���p� �߉d'��n�����ѾW(��aѕ�I�����1P��Bq3��@ye�B�P(�ڤ:��<��SiQ��L�ԃ�l�+
�B1N^�BNTʋ��� TmAО�]��p��`�Q�BE��$��O�C��m1���*��UT����yGˈ���TJ�P(̜º�����	5oT�K}0? �J�$���'`U��� ��Ɠx��ͷ�^W(
ŋpy�o�T��K6j^ ��?+�������fk~Q^̍d@�DSC��Hc�v�+[���+Tl�޾���+Iv��_���}�+w��_���ƐM���sA��dd^:�(>�o�m��{[ᏡMF��m�_x�G�<�B�P�﯄���4ȴ����?�q�^��
<,"�,��b��<ܳ}�+���`6A7�g]�÷+��_�}���m�_�m#�
�B��l��ů���p�%jR@�ʞ/��'��+N6o�۳n�;(v�����k����= ��sT��6jc�[tpЃ����Woʍ��|�G�~'��u_�W#��ߑZ�{�1�恃�ٯP��E
�����k�o�&�d ��=�v�C��$+T�l��ۜ��	����}��B�P|�����,�J!n��<^	̻�7�ו�ِ��oy{S(��e3����:
�B�<�i]�rʔ���e�5�ݕc�����̳wL:&'9��@<mO��I9�rķ���!�bn�9���[
=n8/�K�����m�iF�}�7����z1@-�$ț��h�S^�xHF��∩��!���Nt�	yT%��^�Pˢ�	6�aMh�3��{g(�Y����S�nI ���h0g���������<���jms7��Y�
i
�br����Sz�m'̝���}������o�={��{�R��}oK��˸ʳI�����}O�P��vD�[�P(���%��X���	�]�Uzv�Gb�v+��x�A�G��Z�d.~������<����m���1 ��h~��*���Dzl�0�m`�e�Ɉ�f5�IH�jxg��)���R;��Qʯ5��^5�,���>$�`3n<=b�7�^��$o,:�71;C����a-��m��jN�P(���ޘ�]IX/m����f���}����7;�L\�p]p+��qu���ǌ*C�ݒOr6�����޹W��x���� ������P�*��z��w&i�YR����?��- �q���|� ����c�O�0��?�ԕ�����q`5W��C�W�����h�>����9G�x�'A��y3�9�{��[����o���Zf�t�~���/(�Vf��l�����B_�o&��	�ya�p��'�� �O�����VF���օ��3��h�ϖ���T͋�!�M0�qP���=�c═�{j�]n��$�z#��oۜ�E��7��~�&r��mA�w��g<�v>g(������]C�=�lBB��h6�8���9��l�������_��#�pZ��a�wW��&<O�S�5ޢe��v���=eP�C����/��Z���u���i-�!�k�y�~���S�u;[�7y���S�X;���r�'�����uF�1�L܋
�b*X�y4�@9߆�������C�F2*��l?X�Ǔؿ|��X�&�<O�Dkb�'ο5�i&ζ�K��=�cq䞥u�*��bT�O���a�J�kc�㵄z�+��T��M�;>���a9��);�����7��?�ቐ_�r}Glμ��	 �R@��hxo��4R��tg��A/]#�(�����o�1wh��<����M��������nHa��q� �/hH˱.,�R8�=�����2�OY�
�{�F3/���2J3�;�ַ�ѪW
��]����>L:�[oN2Z>;���F�	s���������T��4w�-o<�=���'�Y(>��0��ѵ�Q(
E������X:(�����v��'��/&p+�!�JY�ސx�������|��r��8��0��j5�/7(����	��<[�H�p�p<g\�밁+�sƳ9Z[��%c��k��k��;�h������]�>x=�!r�Zn���ֵ�U�(~���^�9�4��_h">[�b�kK�"��g�]	N{��~~����	�+��j�6:3��;�D�ƬB�g�)ևo��{m��_x�������6,)S3�m�8y�5�m��
���Ė����
��
�B�) �M
40���%�w�i�F��ǹ�7�܄R���5V\�L4��B!��~S�{�~��i[�|ݕ<�̲8eܶ=�&
�B��n*��FSC���oby�����6:a�]*����)��g���7Fӓ3��c��)^˘>S�H|����l��dmz	��m���n��/i���{'��~�W(^��"����i#��E�^^����ڼW�Ě�l�lrB�Lq�J��N�
�B�m$�#*�	m�	�w��^ݗ ߃�K0Q(
�b0,��Π|3��OY�B��I8/�����A�l(�9��(��'z�+#z����B%�2O�B�w�8�]�V�-�ׅ����]��w��*D�������:iKbđF�����-�:l����4Y�͢�pD��
�Bц��"x 4����H�Z���=y�'&jw��I9��b�&}
�""�FYB�m1(o�H�K"S�B�P��'���E猖HW���|������^3w�ƙ�,Z�~3�^�Z_'�L+����+T�(��
^����'=p�S���D�Ӂ�^�}�e�w��'���ȍ+�ݤ��o�����u���b�fӂO�A�������&ؠ��,.�����X�}����%
�'�{4w}�:��Qd�g q:�'c~�/ޑ�kC��}�ۿ�g�F1;�#~�O�����-@F�%a����z�V&Ne��}K��h�J�=����i��-�&�G��?cue R��&��ƾ��br!�|���I�;ԃ~
y�zY�n{^��2k�P��W,�wq�`6��1�y��P'|� ����u
my�c1)=�o�`�N�e�n��u�UA,��Y=C��ݔR(籭σ�����g���i_��"��Q�f�����%98�ɯ�h��Bʷ���e���r$��_���סD[��R�͍��Z�����M%��-���%��L�Ӫ;�h���������1|�|�Ǔy�G��;�m��N�D6w��3;�@'.��+안 N�P�yd�d3���*A)@�q�&<�����K9(�:�E��
��1R(�+p*���(��j?;��?���W� F�(���� ��7��Ű�>��#�����b�>Tp�'��>)���mFe?��8�0�8�+�aF��������A��i�a@�KX/��Rg��ؤ^@�uĐ"�&� V/l/s�Di�F��J[��'|�X��u�5���N��Bx�+�����4���`�!F�������,iײ@�Cp���d��ϭ��5
�����ѢP(΃������2v�Ư	.�������b�GB:�7R�*�ŕ�5O9E7k5h-KʯE����<���F���0I�8"g@A��KrF9#)Z7�M��?��}��
&�O������4�e��W���f4�����-�.�y����F��?G8R���UL-@�c��@'uD2��?x*�ۓR+J�|
E+��B�<�i��
A�o�B�2kL6 ̀#@�5ҳ���j
�B�x�j��SQ�����/�$����i-��ο�W�7��@6wh<F�qn�Q �gԀ�����!��XXȇ!�Ja���l�D��&�G��-	�Rۖ�]H�6b!)��~��Mӹgh�B��L4��:�~��	)���h�ҡ�I��N9F픥"=pl:���&~��
��* ��y@�h���3�Nܭ���߼ոU���X��O�������y��=�ς~&<��:����+�\FI/p��-ߞ8�>y�R���^K��-�kV̉a�����<��\޵�찃װp�ڤc�DP(
��87Q;�����F�GGA�zX㽹���w5���4W�}[��L�6��PX;��/�% 1O����F��B/��?"tO'�~xh��G��}b��3�m�z����>K�7X:l�C�ɳ45�*�hl�h�!�b���L���->h��9��v|?x�Z���%����}=��;s2v�U(�&)
E#�I>97mem'��k�,�sd'jr��̼Ϲ{�t���6	W�����.#e\�%y��2�3Gԍ���]��,sf��%I�����ҹ{�����4�o�S2f�*Ơ��%#i<���#GGn����]��z�讹�{$7t�0x?�	�Ž���*8�;��8���H<pP�4��z�ʻ��ѡP(�����pVo,SP�&WY@���?Z��E�SE��B��Ắ��#�l3��x7����23*�Ν���=�q[�{�{�A�!U���0�@�z#D�� LG6��DȪ3��0Sh+J_)��L�m3嶵���1ns�X�&�t�gh?-
����Q2�R�s{�}��p$9L�ʊ��$z��S!<bBWiҐ��-�8�
6V��_�@������0ʣ�J	d���Ӭ-zt*B��~
��N�]JE�t6w{G���`Iׄ�SS�i�3�3��0�'q��������ļ'kf�۱o�O^щ/]	�}H��vj��q�����}k�o�����@���g��>������	�j���&��85�4-�Hw�I�4*�0�fw�y� <��O����rq3��&��:MX����H<p,�(�	Ay�)�N��w�g5T(o@EwG��P\�qMYq�O��u��`l�s%R�뽺�f[�v�
���T�j��[�T3��{�-�i�4��J�D�N>�è�����a�&�K��4�0^�)�PK�#�b+���l���3�rZ�m+�r��5��&S�c��|D�	y�'hS�IB�O�?��W �7����\�О��&��5y��th�@X��v7���@Y��o/hxۘ��XŊO�i�>�E����S(w��/����2�}�=�:�XǛ�U���/�gHyfWE���[���?�2�5�<XB���H�����z�Z�3�������rƜ������v��C�׮����:y6����z�[�|��:cU��e�o>�z����q��a4�8+
9��f�z��5(�i�&�i���C��C�~�u;t�����o��D-��� ��]V�g�^�o��D�g����i�S�˒��G�t��縥�αn��mQ�u�qʹL��EpEp����'��J���U1�.v|��k���#e�ӧg�,���o�懻�%�{����0{x��}dX<)1�C�)�5]���3�B��6��>�U�X[?q��'\kT�Z\{�w�YΈ����' �OX�)=+��v�8�1��Mg��W
a��4��3a�}��B_3hy!��h�=f*�8}pL/�S��!�	��g�/�>�[�c:0����Ѽl �A�Ȇ_/4��	ڍ3"�yA�i9!�aq������i�w��sㄜ�%��`'
���qX2����n!v��gS�!y\>ŧ�}�M�yܪ|$<�thX�x"�X.�?�WI�g����=g��Ӧ㩏�P�"���|x%�m�@p9)�z��C��mL��>Q17��g
���l����5o�3.��b�k>Ԙ`�O'�$!?OAz���ʖk���B�P(ZPf�-
6��pn5?] ^*��BT��¨�()���H��ӗ��`�	�4so��+��u�р��zU��&%��	�/eYlw���! ���,������D��QX�S9!��al�̼p��SRX�Xc�<9�)nA#G�O
�B��	������?�o�&���b9���pxv7r���I�dp��w���)$�{0;X����!H����U`&��x�������W�x����Q�A�7�J�������i/�d�Ɵo���J�s�]�g];��K�뽮�x��}�5��t���gX`�#�U�${$GJ��h��w�����u���
�B�x����b���#����KQǬ{��?B�Anh%'���%Y@��Q)�x�y⭐��a:j���N�^
�,�0�ˋ��t���C!��Wjw),1z�헡ϲz�6ѹ�����&�V{��}mez�UN=���⑔��<�w������M�9�Y�B�Pt�z��b-�z�����`�"@�@��L=N[yc�gt�+L0ٛ�L0t���G^��	�j�'�,�Ef��|ޛ׉|��v:�E��M_�黐\1ٙ�Ez�Q�Yq�i�V��^�ُ�DX���܈� ����sv���
�Y�fN�۪��Q���/��lAɹ�iIׯ��c ��K�|[Ԟ��8�Kn���\x��sF�����R��2��R���2�衴����G�;O{� &��>�G-m͐���>��@�����8&sWM��5���RA��vz>�2�$¹|Ax�`��Z�P(ވMp���,����!�
�Cxm�g���i��
*4Q�w/�rP�>���l�qaQK/LLَ�~�褐��G�01:�F<�`���x9h�p0�`���nyX�v������e
�����czږn����	˕�=fF*6d�X���W@RW.�-s�D�[h~�9�W���.���<��ʳ�N�P(���7�2�u�<��"��Q^1���OI��CB	�chnm������e��Q�g�vB����bۜ��D��y�r�&�UKvg�4,~/�c�_��<M6�d��R�h(�C���{5��?�M9N�K��gH���(���M�6�����-}� �Y>y:�q���aU�X�]�p�o:�+k�����O~�>�6��	���M<o>���U���siFbY�	�׈�����^c���πC({��]�b��'��S���n�
(rJ��k�,�O&r�!���Sr�PR�����kݔ�(��(�{�Je�z�ȕ��I��׺P��
�9���os|�p�sK�!����)���4	g8��R�T�wV߶e�Ǹ��LR�P(~(��5�����2��z�W����3�80˶���ъ:�g�rۖ�8x����٬h�a	9eˡa$/h���:sA+�t��}B:�Ȧ3�������e� �_���U���v�&�.hTaC,*|K$E� Q�P�#Ƀ�i�D�$.����ve/?��cF쇳XC��4�J�P(3 �㌽�lmD������n�٠W��h���!`@:���W��nI�;����Є��\׿g����`��H��i9H�ىF%1Q�c�/�ސ}��#�qW��a����C��A�d��/��\�,��-���ъ}�Ƃ!qc>)a߼�+ DsY\|����/C=ث���G�a0����q쿜aC"�&�������i?���P㿇O�r(Kz&*��X�8G�z���zB�}I<h�M�2� ��}Xx \��o�S�c�y���6����2���J'<|�d�[��AJg_�P����Q����kA�u`	����E��l�1ɷ���I?ċ��9h�����JY"��ZwԵ/
�B�8� �KdN|��'A���o!��Y.�x���`�o�-Up[����O��?Sĳ��?i_eV�^���!��c��i0�ȴC!��l�i��Ѐ@�ٶ���0��eO�8
�[���D�	!R"�t���8W��4
�1����~��ؐ)�:p,i'�ɩ���k�b��\¤�*J�U(����x.����,}dY����I�g���G�Ce���utk?�~�@��!`j�]k�������Y��VG.���ߪ�v��*��T��￳�`c�ԗ���Ԫ���T;��v0�R�����F��=,��?]��2&1n�âza�K�Q����]�i�W�E��|5<�I@�h;���i�YtϢ8aV�����#�r,�%yY�,�je�<"\AK�W�Hu��_���a�^4�_�ٶh�������)��8r`zz�� cʷFw�,�8&��ϗ����
��	蜨�~�����x�0x⦽i^�,�;�sv�:I{\��QO<�g�S��{'�c�Z/�#a�@ ر������Q�AHw��ќ���<K4\+��@mwZ�l�bƗ�u�G?�m-{v�'2�H��	I\�;n�}��@4g;���#��&��ver,�Wx.k�(��um����bq0	�B(
��aHv���Wf�I�y\����Ka@M���>q��O�'��&{?L�[��e�"�&��Rd��?���U�s��-�����Ŭ�����d�@��uF��f�����{����2v�̎z�|r���J9#$>p<lϷ>�y�tL͆/&��vĭ���"�>��L����`�H�H�����.if�U��q�G��i8?Y%w�&*6!�VL����Ov��1���'z��@⛐&��t�zH�5����y�I\�(I���CK�W�H�~��S2)�YnA�x��G��^I����1l�b��)$�u9F�E�0n��PGn�h=��E"�?�/�/��MY��P(��Lڷ�
�3@`������g	e4R���z���^��^�Yx	-�Q�>�g��d�exI�C^,,�FH5�4�t�����������=�I�_@(�C;}�������4=v觰ה�ˆL�U����@K2 �Oh"�څ�I��9� ��I�yȼ����Q�O���*� $>�}���Xl;�uм��@�,�Bq3Y9�]@�.ŵr��,KW"�66ٻ�#q��ef9h5�U�h�@hq_p��c5q�jm� /�6W��2��Ҙ�꜡l������7e;�@�4��i�xN��V,XR��~�t�5�W2�VH���mh���O����Lh���\Gß%4�g�5{L4pI�h&�$���?~s:t�>��(�3�o�z�ë�T��z���P�����y�UWӃ�yK����D�33�;>p��;΀C���g&0�/�D~3~�x�4��A_x���h�G_lT�L`=�t��ky�?��5��#��=��Ka��J��������3�@2Ȣ�1Ap��<��uc��#g�&{|N�<��P��]J����3�֘-�3Da��,Y
�B�(�5�R��2�f��Y��.I����6FM����n�0.K�9��s(��L�W��ϲ|9BJy�B؁g�8By\E`Y|NCW����0l�J;�0~u�T�!QZ�,<<#B�CyDn-Ҁ�A(@`K"c�(|��X05���x�4�H���1ĥ�ӌ�#��85>�
�85�
�]�l+�v���w09�G��� �����
��I�����2n�G]	]f�&�zCʸ�$R?Pqm������b�Y{).~���K{	��٪ֺ�"o�+;g4�=��-�$����|o��Q��ܬ/w�#b�������V�I.��8����e�1(��|���dl��;$�)���!����6�U���{b#��Vn����1-�z�����=�k��c�'e�v���G�F�h"�ђ:?�IlW���I[C��z�t� �ϱH�k��C�Mhp����>�
�|�o�ي&}4�v��Jڐ�ӝ��\e#]X���C���dXqܳ9b��s���h=�,�w2��W<�h���eu�H������E�����Y�އ���Z[��i.zGp�ޗ���M��7���Y���TyD�B����Q!�hA`l��F��y��K<]�Y��
�Bq#�?�Y׀� 	�~3�}(o��T^
LHJ�D�q�ᤘ��!/)�j�IX�r��t�1�,}��R�Z�i�}�*�-��i:�/�I��<;i�Ry�>�^��i�Ѹ�!e$}n�!�����9��p�����H�:�v�p�R�Su:���[^�ܴ�P(u@��d��R �;R���*ݵ��;sqKz �����T��S�fSv��_g�`���Z|@��i(P���9n��7�lzeX���n�ME�ဒ�(�&��{JC^;k��P�ua\���Rf⭁��Ճz�H�r�؇��Ԁ�_�3���xB04ᱵ�����P4�>�H�5ʏ`=���I��&�-|�9?-�+�ƍ�`�p����8փ�Ty�K�4�W��pC/	hӐ���
=�~�{ a�G��-�eY(c��)�tq��˷��n�]� �lσn�Z�ʾ��$�� �B13��M�c�ٿ�I�m��:��QZď,+
�B�H`��+X�]*�P�
��<Q��>q�@���A�M��R��o��Q�*���h���hhL�=VP�0L����eh�L�vk*aF�O�n@���kmw�v*�?���^�x0��w� ��)�:���j�$�A0�ǅ��ɈY~��$�>��B�8p��.
�B�Ѡ�=�z��v�|y��p��O֏�����r���0�yM>��\=z������B��>��kp��˽�p��vޅ;�?�b�1����SC��m��kS�/_�B��������T���IYr�,��t�D��f�P(� ���ۇ3���O/�/��RTO�87^���m�;w�\�f�t��N�%��P(~# ��5e{���r��W^�z�PL��#�}��F[��f�x�Y�c^�)���!	}HÁ>f�,�R:���0�m�z	�m��a����톴���ڝq�!���P���{p��X��F�e��@�F�x����&?5���F�P(
xt���o�G��N���t�L��>ue�䝠t���R&߹���r�=nO���'��+CZꑋ3�-�od�P��+TҾ���u�%�e��0r�(��h9�i��(�Z6�;����vM,�v�B|e}k�#�vfb�Ҵ>;���ߕ�]8[�]4_�o���[����1�4�d�I��8�J�9F�m�pcs����w~���@I
�V$�iknw/vq��P(ǨY9U��
Gh`�����˱�q���S�)d�8�������}@�A�Mz���$D��DoH��L!,���t-���'�o�rΆA�v��- �����F�a;(� ���9
�i(/�ua����DR�Ǥ	��('l}IXb���i>1e���y�l#��xx9Ʒ�^Epm�ݖg�h�&ӑ���B�P܉Kk��yܩs��_��]�z}� ��+Q�z��VqE�
~;�7�_,K��}I��W��Ƈr�f��i?�i�y��%��\�J�tN�+W/)�D[)o�g�������!}�ꕫ�T/�Yn,PP=e��Jc���\��;�J�������И{kts�6.��)=o���޺\]Bn^I���k�ŐN�rZ����<��/���֖"�
|1�)dC�� ��Y�/��g -W����&�BZ�x��3Z^K��,�R���-��Z�-���N�XJ���+��(�5�����@��Y[Hޥ_gyw⎹%i���`Әx�k,��?��~�)#��~���P(o��o��s7�՝$���y\��8{������#Q��OHT���-@P|GCT�¤r0��7�t&�^̳T/�Zh/��R�9֯D{��-a�m����ԁ%��2���� ���=����~�+\<�W �m� $4%q�>�L�k"�#/�a���w�S^]Z�������O����%C�P(&�_�)�c]�D6y�z���#�����Xp��!��d�����?��3���t/�|Z���r�yY�ޠ�O���?Z;x=x{rsc�TV�ͤ�Ku�u��RY-���A�.��Qk�Z^�2����j���|m�"��㿳�Y�{rcM��@��8��)������������wi��g8Hc��q�����Hy����HiZ��Z�Q���=]~K>���w�S����n���o��74��w�`�����������n��O
��&�`ga���F��^�n|u7�v�2��L��-b)�)�e��rk��n�E+��Z:HÒ�0��;hG�8o+��ZX0��r0��q�����q ��7����8�%cy�'
�:�|�������W
h�0���J�8�s<>Q'��d�
�B����D��e���W>o�GA9biՕ���!r��nQP�r$�%�t͈��h�+�s�&�����Ո8�?<�Z��<$��\�$C��A��ܸA�-'W�^������Wx=zߩ�w.�iE;�n����p�����%�uB�<�� k��)��O�h�l�Z�m�Mĵ�-��˧ǚ�T�\��rjek�-����c��폽�9H�<��F{���wɇ���SΥ��(��f��<�B�P�{�6�.r_��uhcVW�3Pf�B����>����Bv_[ ��ƭ�u�����0a�s#��X�YwhT������ �t���l���Ҏ� fG�)��Fo��]�Ӓ��q��9�}�M+�J��!fLB�wF���N�����p�]z��"s��B�PA'�6����>�㵛���P�������e��c$:����r�*���=W~^��>��v��GkY��o1��y��G�������fP�R�Z�r�ZfJe���qr����rZ�k�1/��;��Q�G�\	5���#���ظ�`��,I�6��kqPz:����F}6���?����G��n5�?e҃_��KB,�coC����[~	w�͈-����Q�����sl\��$�6p�B&�ǒR6>����La�ǩ�u˂o� ct�P(��q�q|U�6����
5ܻ'�l��z�(��y���aԾn���N> 
��B��n�)��1<͔'
�yq�>U�Ky�t#������/���^Jw�v+��th !��O�P���ı"�S[�@b9p�����$��; ������H�@ƌH�xY�9�����p��Z�P(?�~E��l���Ȓ�L��{����S衿ft��JqP�Ԣ��R:�*+�������ߥg-����n��G��Bj�\X��Vc�\��U��i�\��8�=��zލZޥ�R�ڻ�a�:!�f�_Rģ�o�0���M���������h�k���Ҟ^8J���p@��i�����!��<a �!){��Sl� ��]��_G�&��B��e�kͻg����qu���=c�x'=�r��O���������;���(�:�f�qa?�
�>5^ϲ����,k}��Ƅ��k9�1G+��EX3p1{��D	����8Q{�3�1泐����Z��n���o$f�AF�D��)��sT����+p�桂�c��$�z��Dq�􌾃�@&��xK��ꊴP��3s��C�V��k
��Ja���baaK�h��т�7�+����� #�a
A!�F�:����}5���E��ۭ���x�[��T9v!4۸ ���ǹB�P(2��x�I�V��!����QS1v=�jڿ���%p�baӴ��T�e|��������J��~��kyN�����7}/}��q8����;^�ܾ��#���P�{)�͹�Im��Ju���g�T6O��g-��˦e���V�\)o^����ϵa�,��S)���(գ�]%�ڃ��y��S<]Π�uޡc��qL�)2�G�?��9�H&�,b�ƭ0hw"sԚ�v\����	w�fhKzH!I
��vu�]}6�}<Y�os���:����B�9���C����H�Poō)�����`$11��B0dȬ�B���r�܁d� �O{PB��zY���4���U��U(
��Ow �ٝ��T�F��0�p���yH�G�,.��P!>}�a�������dh�l�=�P-�7� �hG��I{���K;�-�G	�}ς
u��'�=�ό�ǲ�@�:��1��Iz ��;�z�:��5��b��8#rT�z�Z �%y�x�sV[�P(����7~g���<��2�����Ϛs{���ďD�y~2���ۤ�R)M�=Z�`S����'�j(���8�!N��b=�>;U~C][��W����y=r�j�/�z=��4���z\y�~{��5�]%yֱ<��K����NPK�g��<Zrl�`���SB�[�B��u�N���h�j�,��7�5+,`͝9q�cY^i�RlQ(�P(�wb_[��U9����ɹ& ��������0��<E<>�t�L�J_��u(�����LSC�ĳ��6Ҟ���ڃ�L_WX���h����&A0fc �Qq����
�uB����KUN�"q�̛P��>�;�p�7��r']
�B�;X�u�X5?�Nqu�������ӂ&z�o!�L�Ϣ5�C=>خw�z|�^g�g-Ν����t)xd���&(~:���'�P�L;a觅�=;���N��.
E��?%B4:��
�Y�w�'yሮ�L�^�wJ8���\M:㐴�x2��(���B�P|c׾��N�Oƭ���eF&
�&�	C.��]���h�T�����)��^ՌE⡒cy4�F{.�ض-�3IL��C>�r��qqHg
�ɳ�(��A�g���PwH}�y�<И �)�C����H� �ͧ�@��#Y��_��(
��U(�.����ܺ��6uA�_�c^��.^	��ϭ�S(@��u~��W��i���jd�wN(�[m�哧�Pِ輌5&k�M�GX��_�noM6�Zq᧿[^Ч^u�P܁Y\��Kt[�.���	���O}gÝm��!,���Z��ڂ���٥�\=�����[@=p(
E+ҹ�S���cf긦���k�ѷ���'� �ePan��:�&�� ��ҒH#⠸'	��j,"�`����x����*}gÌ�k�J9V������$O�24T���pLg}HR0ʈ{�HC1�;q[i�4bI9ý�)i�؉�JRKܘ�i�|<|a�vQjjI�+s�P(����X�+	k�����=^������>�~$lE�}�?�V����P���+�D�Sa�b|ɓ�3
��:�����؇tA ǲ����o	^�S�~@�#$�&Ȍ�Jʦ���eѯ]�1g�Ӷ��}������b�p�A$&x���/��1�1/�<g���+IZ<(~|,|R؇e��Z-��X�Ly
��^��<�Ա� ����R�L�����F�]Yb-�g
�B����?̓���P�	|щ~���RU����72�%c�,1��t�&
'��9�0�q�g�<yT��yrս��A�����t����t�Vj[)�,iB��F�>�<9�^�6��>�@M��_���I�)1�q����Q�@b�i'��x�T1��j$�6T�{�d^�[T�a�ݨ�*��*
ż�Κ��"�ӎlߗcTb@��?8��5[W(4`��k�A���g�ҋ�pK�7<ַ8�k�8��Z���B��￴��9�~q��]�	K��ע�ċl)�~1�$I���i�l]�O]�bq�~"�S	��2�l
G꧞rQ���MG?߂'2�0��4���(����p�#d���_�� ?�}��)
�S����ޠ��� ��ij{�}��kә��mH�;50�
:�a����Y��N֤� ��<��ir�O�q#����.�gh:f��+�{w��f4�9ځЎy&�!p$�Z��6H��@�����X-8��3$��y�]K+�er�{G�� %����vV(�w�.�ǧ�7��"�t�1���߉�����[��E~&9n���d�
���2��u|[�ב�4���+O@�����5O��[���Z�Sx�izE>�.~K�w�����y��fI�$��L�!�3Y���j��=[W�y�
��v۾�F�P(�>�?p��0۾�c�p�6ց%�$�0=K�x���C$]v��ʣg^����;������~�ӕ	K���e헴m���z�6"a�J{�m��.AfH�6좱��5`�nÑ�{\�)��q�7>���𩡇�<�C�k7/�3W������S(��n:3��bڈ�χ�mJ�߯*3�ݩXtER(�ɱ����^ �������wT��π�FcߜB�,��4��������^7-J����E��7<#p�Xa�R���txĈ>-�3�0�,�Ht�)ϟ����� +ۼ�:��õ,�����ڎs��<pP�9������C�P(z�|�7����t�9;�Rc���M���<��,�$�c榴��F-�h����&��
���y�0##vH�y�=�@���>�Υ�j+�-���.	#F4^Keioh[Z�K$�'���>�#��������Ӽ4��X^<�j�����ǀ�{o��2��E#�=��!�yN�76Űt
�BQ�w]J�9c��A6y���m����r�����i����G���p�a&	=HV�0�|���4+W!�{I�,�i�`����{��=�"�+�Ws�{������Fzq�
�}I���a^%Esh��aZG�����g�ҝF9��ښN`�T��ܝP��:��$wm��m k����.Ճ�)g���Q2�8�~�׭'�Vc�^#�Oz#�mH��ߺ�)�6.��a�@1�S������0,��Z��;��iDSp��m���'��^}��_$�(<Je��3�[�B��T@N�
�fN������M���A����m�L|���{h�g��ry�21���,�|�!,�2e��*�+Չ�wH� a6����ҭm��Qa��0����=ɋ�L�i��D�+m�ȿ2})��y;��}(Q��1|gL�H^LX��qZ,�ı&m��o��#-d�o�B���]]]_Y�vd����F�ʹ��� d{'A�$ބ��[�
ůC�o~^�C7_a���}\(v���Y{�m���ׯ.���<���w�$À�F�wr^@2���Hk{�����-�s��Zn���A�\�$^�S�⭨Mgd���Cu�a\�[�%��_��C��"���1��.�#����+��E�����?��G�Ju�
rF4Qc�G�@��|c��ĸ�|s�_ɂ�ǓzۼT���š��Ҹ�c��Mr�r�(�&��$�Y8�;o��xΌ0&PC�`A��Ɔ�ȟi�\���r)�n[�B�P�(����Q���4{n r5fxVA9鳠�7��+�s�r�C�R9��#�'4Ps�(���0NS�r@z�Rg�u�:��4��E���@�+ҁ��a�i:0-���n?A��S���oR�!�@�߂O��X8&*��h�P(�f�z8��.
ە�N��y���ʾ�2��3���EF�TNA�+�'��*�����[MoÈ1=� ��&���r'�~���n�Jʣ�P�	R�B~D��?$�'t��C����?e�a������wV��MϡyJ����6;9C
���)O��2x��x����!{H���%�r�ID)����7���~����d�+���H��pql�&x��m̏&�8��/�Oˡ��F��:��L�P(�AXg�s3}���EJ[s�Z�i0� �H���)�'�p% p/R��;)��nIe�8�����,���:�8�-m�E�@C�=%F ��Dab}�Ƣ!Fܚ-Ob{�����Ɓ>�>,����(�{�&�nR\���4��P(� <�D�* �-oк7 �z�V��ŕd�=�z�ງR~@� y�S&,�${�g �s��Y�m
'{H�cpf���^�������B.��ǥ\��㑦�37oH�J<\��8H>�g3���g*�N�sʀ�߹!/쿪�j��H}#�t�$�XɵY)m-����ţI��C��ډ���O���Z<sqs+<��n�������������	���,#p���*���}'qC)�̵�B�P(FB�j��ƀk�ȗ�du��u�}��ǝ�G<����D��,,��FisP#b�i^���^�˕G������No^Ŷ�B�Ia�:���4�Zh7�f�v�@�Å�x1��1i���Iʷ&X��$Qa�xNC�����=�j��ޗ����q�}~n�3~�,2*��x׫P(�I�ٳu��x���^Z&-;��$��Xd'o۴5�t-�<�/����k��d�8l�b��Wޢ�hUl��<��_��X��e�����c&7�{y��=>�ϥ8RYw8�ʔ����~'�]�M�E{@b����q=֒�r��r�3y����'��3��)0B�5
�K�	�]��Q]WMa�� �q��8t��
�C.�-��6U5����=c�͹>�EдW�����H��\X)�Mo@�
}��nc�Z>����^�f�1M<��[��%Bp�yg��c�ǹr-�Zo3-�
�B�:l�����؃G�m�A�y[��B�vW�:N��Iܽo��#��~h�^�[��]�JngP& �&C �+,���1{زp#PE?@�1�%	�4�g'�h��#����ڶ��L;p�J�(}��C9�T/��{Y|`b>G���*�@,���F�8Ć�#]iC����J���\y#���_<B�?ͧ���NM�Y�O1���l�����`$3�G�P�W��C�}�9;;��~�u��eѠ���6�̿M��h^��,hX�����~r0#�3��$�7����R�C,�<��qH��O�Տ��L<��|S�s��o�/=�Y$�'fr���&���y���2�`�>%|'�/n�@��l�F�����#�0���h�e�g�v�qA��)�/��ࣛ*�me�ߨ ��o��F5��it��i��鸋�pz��5ވ��#F3�kc�ϕ���g<��D�>v�`[��B��:f����?q_B�����x�S�`�`ARt1=�PyO��A��ҁ�Y�m�������@C&��n
a�tZD���U,��^ �_Rf-�P�!���þ�K�1�q�{Hu,Ǆ<��j^���������l_R�O/L*;��r����{Ϛ�
�����\�|�ZC��@��g�W�m��M���Z�6$�S���I羁�,tKC30f�Gڑ|G�A;鷧�@Bٸ<'#x�
|�
���gK�fin
��h��D���'k��ֈ�ӒDJ���] @��pL��h�W!�Ǟ/��p�g��'Ю�Zz�7Nr��)ݪP�r^8%XD�w��zWW�LzkwA�3YN�v0�e�	7c��X<k���M b?��ޮT(��֎ U�k�y��4wC�m�Oߣ��mA��Bb{��G�H���ć4/Xh�VGO$�h�4Hy�0!]Rgb�ph#�U�y�Y�Ű�z��9�13�v��мy��~�F��b�$�T�Ā�g�g�7�(H^�=Iî�V����Eq�W�d�:e���X�	 �߽��(R(3�}��͜�g�A�������\|����fr��ޫ%�ŭ�Ԁ;���O�����޷b��P�����(K�nZ�X�~&��0������ʃ��N��Ƃ;���V
N^�b���w��	P尷��D��0�+L��]��,3��#=4���}�7�����mG�j\}���v}�V��Ҿ&���k���̏��P(���>\@�3������ڸ$�A�!����탅�%c��L�g�* n���q_Ȇ�����}i:X�	����Y!,ı�<i ˋ�I�Y�Ԍ�فvN��gR/!L���}fxXK^��0++�I���l e'8����#�|����y�<O�<�q*X͋�a, z�s�j��Gzq��4NE��eY�Y�2�'��EH���K�P���3��(ٮ�c�ȁ�J֟�kON�ɯ%�ai��!�_\
�|%K���<S�,#��8�	�2�4$z|b���hvI���)��"Jx��"�8b�A"H��D3S^��������4�S�p�Z���.t��b$3K�5-�_FɊ;���{x�w��5�/��?��F����� c�!�ߜ!Ę�,i(Cd��4ߡ��
�Bq�ޓ���aM�i�W o��G��u�i��̓F׹��v�k�{�\�w�J�����h �·D��(f��x�,/�Ư�������pȳ1�Ӑ���eۏ�g�]"�Iyf�,�-�]�/�'&(�%�R�g��*{�ut���Eˑ=p0�� �V:&�V��d�7�/���Q�@��v����2`ч�xuJ�k���'��3(�7
�B�e��QR�L�P���KB�pHքD#�`�Q:E�x#����J�s�X��w��p�B���kjr
i�D�q�|r��G���`�9�&����X���C�������ӊ�z0�5r%�q0dYmu�����į��e"��L�o,�w5�� o��l��(N��\����R�ｃ�fe�a�o��)҇u�����He��c�*���:�7Z�ْ�^?/O������Ԗ���V$����S>����4h��lfH�����'u>R(�~�9��:]�V��XB�*J�;��N�.�������o}�OT�-�������]!�����g�W�|B�,!	.��C/#K��gVz �WY$~|`!�)�e���VR�!���l����F&��ڟ�Yl��B5r��HY�H=�ga>��1�]�n`���4�]̃��(�c{ 3b���)}/�
�Q(Ӑ6�.��e�ǫ�?���h��a�H9�����uܼgM���2���1x宫K� rXԃ��c���T?�B�=PY����m��V�vy>���]8�g�ϭѰъ��_�c2;�����Q�"�j��@�J,�{;YCI�H�i*���C���F�8��;6�\nN9�iS(�����;F����7�ܔ���z�4�#�`���V����O��}��x�}���yK\҇�J�C�I@�W��vu�zX��;�����
�;W�OɅO�w���\��	j�aB[')�L
z��9Ơ�F�V[|�k����,�|�r�|p��T�� �OI<�'J�}>��<�P(�!Q�Cq�����
ϘR�ꆥ����ϬxsCR�>����?���C�=(8Ƨa�,�3�a���D� ^�4��HF}/ö��1���aږ�%���3B�kB�0f�$9CT�X��aK)5��-�P���-� a�,_
@2&]��P.����z�K<L+��Q���O8D�����
���Q(���w���¯�hL�u���z,��S����mu�x"*��PRڕnZ��9Լ�>h�P(���o͇�yF��C���?D�.��dz[�����t^��г��~\���K2�=,�4�i˦Ӏ#6T<��N��Ù���C�͝D��LW�~SZ�0%�U|�zo]�L1V1=
;�o/�i#/-���A������IH<��	Q��B�P|J6��L� �V<1u�o�}V��� .��*�+��Y&�1�0�0������N! (���H��a�Ȅ�C�H>Э[+}�>5���tݦ�%y	�Qc��ɧ5��TC��a�[#u��8��,c��ԓr�F�$��|��Irt���&���8(D*��Y��~:f�s^3���ў
�B��xb:l&{X�O.Uh�)�E!5@$e�Z�j�Or�w�+Jy�0"U(���C�%��=D��L�4���rT�z=k��C�k�#]�z����%�ͷ�
4x���D
�L\ɍV]8�]�ȆW�S>������6�a��]�,�T���}-m#���hz�F��_1⠖���������
�B�������RG��q}E*���j����ڝ\�q�y���RGQm|�}=1�
��P���f��B�HX�A2�+Zj�a�*a��^��$}��C�+�g4�O��C�p�4��Jm+ԕgE��6
�tH�P#BO�5���9���fH��"R��9��������\�AM�ʭ��	
�B��WRwz�l�^ȥ�<Lxւ}���z�L��E�H��G����[0�C<Js�Wа]�}�=�9�@��P(ᆅ�aZ�H����3�%:�(��6eX �@r�{�i�����d�~�"/��80K�}q���yps�7
s� �~�s5'L����.�ZIW��Q2,��G�Ң8�>W��J�ZY�g����+��sK���jE�x:�����r�k�z�W�=��Y[��2��b�|�*գ���"�ԓ�A�k��\��@�s��iȾ��)����{��5�,����B�P���@�Z���7��#�d����o_�����Nd�������5�Ni� ߳R�A��o͗�L�Z���vB]k2ɘn}g{!�yJ�[�� ���yU�h�p�OJ���%��w�Z�C���K����<�:�h0fL�h�By�.�\�,��d��0������1Q<} �a�t^Jߛ��ޱW���|�m3=r}H��|Y��r
�l��(Q(
�g�H�wa�+𾿀`t���7��9��<���PY���j�a��nC>@��2�*�{7�.�7aI�q�~<Q^�P(>����7��g��d}��\�@Y��1`�,�3�3O#�)�x�\�^��چ��U̴Ӏ��e�w����@+
:�l��7)��3`����NR4��S�3�����2GBz�s����ڵ��o1�RI}Q�3��BJ�R~�=rF1gP��ʮ-R9�[�#�>�6��A*Ku��v9��TH�2;��؜.�OW�+���;�F
�B�5 jG�
R��l}f���T�xA�̄��Y�I>[�d��/�Y93��*�+ǁB>3�МaMF�	ՠg'y�0)/B�5i�bX�>)��T/!LB.��(���R�,}�@�쐧ɴw#W���)��9U0Xgjh�C2����
���"|���7}�81�`XH$\Z���S��R�UW2J�KS�/n}�B�x8��߃ɠѠ�����l%�	�E�}��K�R��B��W�8��V���<lF�lkj�%y<�[��W���\���\�Z|N.���BO��Ȱڰg���T�P<
��@m�v�ֈ�b�y�9�ǘ#�,���\������=[�:���`B�d���5��tW�ȴ����уڣxI샃��Ռ�8L�D�yv����5�ᙴw�G�����_FI��?KqJy�Ƒ&�3���Zf�x��OF%\�&�~��#�㏛q��w��*z*�?�xcC�<������g������������b
�B�M ���3�g_P�ٹ��H�5����H��3hݧ^��m��L��.Oۂ�܏"x�ɘ\��N<�O�x��j��aR�'� �J���Ha���C^��ʼ����)�Q=a�LC�?�i�|#�$���S{o>1$q��BB��}HL���N���$򃷀�m �ii]��B���`��T��`PM�G��8�${Y�����d8�_��m���o���9�n2T���E�q�g������o�����T���LW�8� �H��.�]����5Xd���Y���Ͽ-�R�gP�ѩ}����Y���~-.{\ul�~$�˟�{�ë{��ƕ.�؀y�M�W�����B�z^�<3ȆJ����0���H��|��W���&}e��b��Jv�4^�参�o?��Ҽ<6ͣk����~�����۩�|�,�����]���?���s�H�"���(]�7��A#xxb����J�&Ϟ�O��6���v;�e�,����k�ۄ����ɬ�Z{��Q[���Zpf�� 6b���+S�7�"3#Ѻb`�a�f6������m .i8�pwp�)7����|^SY��
w�^dp�|.hz|r��ڶ�A����߁�biLf)�=�LC��@S��N>"�4��n��9�O���`�D]�/X�`��_s~Ξ���� 95cKr�ͪ����2����;�u�A�!��v���nȨϻ�m:�Gj���y�;�J�n��s�Ys�!Hp#��y��1TO.8��>D*_I��ʭ �r��\y[�)�X����a�h�p���JDƟ�v��'����}Ѥ���8��֞R"AD��t)�~JV�m���x����4�n�T�:$��ū�o��#d_��	���<w��iP
w)�q����F��v^p��{�`����	�F0���~���o�J�d��x�Y��i�/C�D�|���-=<܎�l4-��l��\�f���\'�ᙝ4�Gp���4����%#������y�N�G��|t��)m�N��+�=٩�yc���������z�j9���ԉ&j|�*^k|�����^���`��~'�:ߺ.��r����2��#z�Nh�D��LVY�b,g�4ځ�O���-��.�C�)���0%[�y�*RSg#t
�~C�2,���7�.�L,0-�-�^)w^љC��X1����ұ>:��d��G�M�\ox��D�?�bk�TH���8�'�_���
��]t7=?hu�kWR~H�,{O0�e�X�}k���֊���ϛ�;��z�l)�'�����W���w���[���q��\�O�_t�	߂�6�$rA5�<��B�T�ޟ�Lma����ux6c��3�c�V�ȄN3(����q
����2���3�G�����:���֓T=�=1@���\��x���~i2n�n�@ٯC�J㱷����dܙ��}����{����A�X�������~�J�	'�:��;e�g*ʇ���pu�b��?h�7�r�n5��*�\o�˳��A8���H4
�'���E�q0�т�MPT�w��hYe�f�z��=�J[���{�V��N��D7p����I�������3����0^m|���-x`�YmA�)J��H�^���*��`~�����+�=i{ ��ˎ�t���5��8d����lZ�7��:7�iʹ�B�#����<>�Mm�����-�ݤadt�;��;*�78���XǄ	��@���`�6ѓ+�<l�2�x�S;۪��
�]�L��Z�L.EC� '�҉�֬�|��*p�X.X��� k|nߟ�o�qnvk�|�Ŝ�O�y	bj{Lx�qm���S:o�x�}~qx<����ru@�E;�����DA��-cІ��̱<��|��W�-!�r�hN�<Ŭ����)�͛�~[q�1��=~_<a��Mf#*03�������;�W��e�я�o@*�G�L����7�u��P���hǕ��!�{c��,{�_�uT��WW�I��a=��l1�?4o����n�Ñ��09� �B]/����>�~��
&=�D�az�y�8��&�]Q��t��U�'�.���p	�G�q��#�|���"���+�ޕ8{
�o� �98�9൹}��s��e�������a,������,��pda᛿���Ʃ��+kw��MM7��c|�I����Ίڰ��7�b�0�@�P(���)�p�G+S�#g%�|<���#;\p_�r�|���A� �JR�`�LƑ0�iu���,وMk�5�˫I�>��re�C^��B��c�����ǐk*L�ߧ<�	��Z�`��M�}���[�<Ù$��|V�']Q(hH���M>�Pn�C�1����}�t\4g|�2]��#�>QV"X
�3 ���6X2�!�Z?&�c֍jϛl��w�먇��.������SE�1��cmQ�'�A&{�c�.��<#Їfl �.��8d���7�P����E���n�ց~�G�
�`|������B���M�� ='w]�h2���|��6��6Q}���,�]P6s~�)q�Qp�_w��ަ`7�m��d��5�xv�Ñ���X�W��0��x���&��ҕ#���v� P�FA�C١�:>#<>򅸠�l]�<��"w�� a�����Z��5�FF��߾�n��PM�e-�K�,X�`���-�T���Y�ے�A�c��0�-�ʔ��7�vq�g������⫭�7�o�~���X``��L����ۏ��۷6O��ivͻ�f�; �)�����:i8�r[�Ζ�~[��(x gڤ�Չ�.����6���Os�	�P�n_QRsҙK��mj����w���{�W���!�4H��%�d��)teؼ�9�pA����+s�b��ɚ ��=���>���έ�v��5���Z�`��~J��79ߎ@\���*+=�o���>L�)����M}�� �h�O/Mp@�oo�[�0�h���{����<,�����|���Ss-AZ��ei�kԶ���O��ni��ȗ�op�J�D��I�ȁ��L!-�M���ct�΅�Ї�X����}`��3�>�O�	�G��,X�YPv6����)[������:�3���g��1��넁@�x,�ze
�WT�{-6_��]��a}���,8f��V����H}E;�6e���3yg�˴��	ok��Bٷ�j-�wi�s	]r����}ݺ�ί%�O�t.�xtz�n�`��3iDeHX�!��V��+80;�q��{��I4�G��Cl�?T/�:�ɔ��B�8�]�K=���.zM���%4e���de�F_d��%@iHǣ�iٴ���������滊	�Ȋ���e騫�@H�v���)����$�Qg�~���:��A^~�a��E<*�)����R&�>�Di<��U����AS�ѱ��Z��݀i���ԧ]~���Y��`���j���,�3#�mQ��S,X�@ �9mvl�~��6̒�;P� (;���a����+��[�$�@�4����F��� ��y8.�I~�i�D��p�Mڰ���&���LZ6�=�@�e�92#<�#�vv�}���#�r�j�ymeqGm%�ӫ�/��^i��f��K���hu�d]S�r!�8�b���g��Y�������)������=L3�*��37�Z��n�$s˺2]���d�����H�x��~��+6}��o�k�+��K6�_2?ve������v�=P���C����TCi�H�/�>�=p�	���_��>47Q��=�NKq.���[ư����0{��>G��\�r9l����H�ܲQ��v �A��L�7�ݵ��e}�i�}�>��Tp� �~�R���;�Gp!�{�=#h*��w�@8,�I6�=��_tT�f��n�HPHE���''�	^!H-Lt��b�ʃC	q@���(Wv�@t-�#�a���N}-�yU{Hh��3��`i'#����e<�ぴ7�h�I�8�{ O4�����)^���QQ�<��q��8�-O��z`}T�7I�I���6������x$e���1��YSr�N�l�5��X��G�����`����������gkl�S�,�ί�{9~��]�d߿�
��\��"�+Dò���ڋ�\��>�g���m��g���$F��JCc$֐��q�0�!�	�B��t��sa�(�*M���Pv9�`p#�l����fpH��l�m����G~�"M!��r��Ɉ�����<�;��L�*��-�Yכ:�Ө~�y84��Y���~���wC���k�맡��ca��J,X��H��5RI���I������ؾ������ߞ�Y�}Q�rl�r-��b}�=�ļ������Nc����i���^L����l�m����{�T��ėr?ko��|�� ��?z(y�'%�Է|_:���� i�8�Gc�����!LS�Y@>��4�S��[f��\�vRk���>M��=�ꚽ�B�ώ�Vʩ���������#L)���.��IgOg0�}����[\צ�Fp�*����tP�Q��pB��a����-S>�?��8�&�>Q��rt����v���v⫟3����ˬ��`�pQ��df���U��ux�vu�:�L�=��G�X���J]{�����`���8O�Y�vH����>%l�����ol��֮���*E�ⷔ����c���5��=
��XƱBpUe!*'RyT��^\�`����^F������YZ�s�o�-��b�N����J�ھ�lSO(w��~&�=8��(C��JX S;;�E{��ȠnAiSA���Y�;�����A
/�)�d�mk���#�2@9��)���Z��잉f�����AbF�-����qx������=�Ӳ����i\����>rٟ�>�Y,X�����u;���j��@2��m7n����� �lHm��;�X,��?����ks��68��\�q�.�Ew��^NA����p&f�*��۽�r����E�a*�0J&��L`~���
�ߪ_�jL��ۉrۿ�0�Y.����D������*�	��D��<��^6��,�J��H=�fk,A)�A�)�Ci;9�u�x/&���0�TEڈ#�o�U�R/��ı�����`(�Ś|&�h���v��b�ö/r��j�Z��{�����(��mc��6O�����E\�G�O�����z�v?̆So�J���'J�:��;gF�v5����Lfْ�G��am�$iT�V�����$���{k�}q�,��Q0�*kw=��w'���G,X�����g-��H����#�0�~��i��'ܦ�P	DS��+���9`�M"R��@�<��yԁj2�l�y�!-�}l>�:^�Nv#_�A9�Ol�nWg�)9��X��p t��}'���9���ƾ����֎��Y|)�I���Ji�,�+�X�v~�D�k.�ߥF�5m���$t* �/C�o��gn6}���&��1��ǺAX�x�����������!�WuDp���~�=4p� �y̳=	c�dh��� ��+�הS�p������wGg�;j�4��uF���;�8��OR>�ic�&�?�7�Ǔ~p��i�Ii�ˮ9BH�g���v��kv=?1�5����=���믽��,�K8ʓŵ�ry��?�y�/�m�.��`3��(���Cpe�ye"#�,M���[���O6���q�g,�݊,��55ZBӳ�3�Hh���ɇ4s�C]�=�i����Y�t6��9�;�M��v�Hv�ű=�~����Cq�{��G,}x�����Ȝ��bZ�ׁ��!��~SO�Y���O3��Rbѵ�3��+Ӷ�jl��.�Xx�־mY�5LH,B8d�I�}$c(��J�,���Kю��3�oأ���g=���ĩx��0�V������gP��,�L�Gyx�޳~O���KM�C"�eu���M���=����,� >�B�L�)~A���r����Y�<(���퍟��� ��;�a����S��s�<	��J���W��7ap}6����mm�|�`8�>\�Qn;�uh_� �͏�*�}݅s���x}=�\��߰��`�������*�v�p�uTT��l#��q��ϯ�?UO$�Ξ=�Ȧ��2*����Cn�SzD��x�����W������W(~D�k��Tv�]g��C�df`z�%t�U�b���-�eٖE��S�b��d���̝]l}+����2������u�;��Fvً	h�֡���H�'u�L�V���,����A ���7���4R�-nL��,;vX�����0]��o��}�@�x�{�Y�k堟��v���=��c�mӑ~hm2O�|����/E�q��&�b}l*�i�\�h|}Qh��<�2b��
q�q��L`o!x�w�;;�p��t��8����4��6ı ?QBّ�(F.�rY>^�Nv��pM��/�m4#�δ�'";١���!�?n��I�ـپ��/�����N�9ց��V`�6�&R�,k�`b~ܱ�a������>�&z�D槕��_Z�~�Uz�P/�n��?�N�֤n����Y�kY��������4��j��_�=��"�J�I�u��'g�����-m?ܬ�e���6=[�u�S���i�V�wo\E6��;J�1��ӛ	�z2��X��J0�4�>��1���ޮ�6$���ҝ@mȢ��p���2t8m&i��k2�G�����Y����s��PNɞ�w��n�O�"�&j#ɓ�[ 	|HC{_,��|���g���5V�����'����}�+U <���|�>��f�U>c�f�����7Qr��+.���D�j�/՗�5\x�~��	}^7��,�]��C,x�u�}��|�U>�-��O��ɱ�N�%�x%��ơ���o�=$ KeOO�R���+��㱽�2o�����e����n�zN��6H�Ϭ8�׽M[���6Csѥŏ��b��8O������H��]�Y���f�l�����!���Ƒ]��C��������F'��clzr���~�CP���m_�Ǚr�f�WƓ���V���m쐗���9���z'��nka�y$�݁?�#v?h�O���{�5�> ?�Wxi�~�=d1�`����a�,���{"�9�ן��
XM�j���7����Q��滿��ZUW5�U[���"٢z�on���N�UR��a��7p|i����&h�r�c�ycEڭ03���	Π�;�/:��S���Q��r�<X��²
���a�
�Pf��J��P>�/��A���@P�3�4���;2���v��i�O�����sX/����fΛ���f9�ٲ���<�Aap���(X�\	e9e��d����J�
߷����V�b�C�qtE��7Wd���J�s��8�=��9��`��?c�Q��Z�L���+k���J��c��r�Aʍ��`��W��$��	�M�Oh2ǩ��4 ��%�ht�1������6��^���r�J��<#Z�|�,G򽌃Tm{䧜��q�l���r���$�B_��yZz�| �3Uߨ��ʦ����v=���C��]��(���'�|,�c��e�S������ٳ_��7/���Y�`�GA�wG��A��7�]^����~b.wq�^W�fife��u5O�wX�◒ĕu2onV�����F��y�������>�WD��ٽ��è�=܁�|(i\:�l��8��G8G�C_���k?�=�����-�q�Wd�S�j�>gNz�����H�s	o���96O�´ڃ�?��U��a�� �9d&_3�a���z��B|����M��?�v��
��ʺ�
�,�Fr
�s`l�$�М�9�_�/�әmt�	�"���;�s�L���E�8��r� �M�@�*���� ]Vħͥ�ca�r6J�p���z�N#�v�hI9:���OT�������`t��hU]ғ�O��*��`�j��M���=���<7���	p:��%q&�����Z�=p��f���~�D���}�I�ɂ�V7�~d�,p2K�bSd����W�j?����t'��$#���������?e����G�� ����qK���"�ݳ�=>��:���lh�ވ�nT�>�<��
g��¥�����p��6Β!3�t�H��"Q�Z�Ȟ$����R���
_\R��Wf�|$�h#�3Hӟ��tWl�#�*^�"�,X��!��w���
���o���������ف]�H���-��P"�1̳:��u<��۷�C����Oח���iۦ6�o�l���!-�~ƿ0��#�2�n�o�P'����8��a��N�R��E{1�O��eh	��Vڇ7�ފ�#��(K��F@�0�z�o�k��؃�n��n��ه��'{�Z=�o~߉�D9���~����sٛD��0G��g�����!����9��d�E䕁bOj]	Zs������>pQ��ޞl��#-�t�ɐ ����BΓa�12��m/ej��g�qy��r��!���ށ��(hw�'h��Jכ�E~�CNVB!�����O]�4Y�B"۹�p��@y$ͫ\�>s�M����h�g}�`q䔅��k���6%R�O�Af+z-q��>_!�yK��LCY�{���^y����+A�ć,����~�����w��d�_* �������TZ2#��BZN>�g����i�b����
��u7�8���n��vP~�m���B��v�"�f�Q%��� 1}�����A�$R M��8ێ�@kk�l,h�
�9rL�[G�+��C]D�~ة^i��'pw�yy�h���F7&���)�)��q�4��.�i�~,�;/9�e�{n5?�J�7��k_��(�Fy ���gp�ش,yrj�t�C�2͘�h'�g���r�c�S�o��k�"�������L�������Ť����k���q� qy8�-�XqK�j,&i�ڃa?	�p��x#`D����mk��c�Q�J��CFx歷w�o��3}���0OK�Tze��������j;_:�a'f�X�~��	
�(d�\��:
R�z"w��6��g������nֈ6V�ǧ�&+�QWE8�8ׅYU��8}�n\N�y4!�H�C>l(��2E�@v���g��������iΕ�p�N6D:zP�x�:Ԋ����d˶2Ԇ�Q�D���8T�GѮ/W�o�{�z¯��%�v�^��;ykH� �O�V���.F%�k�TM��>܀��d�4O�OR�,Xp��]b��V���G�%3�Ò��VG����l̳x|�}��Dp&�l}��rW �2��n��fg�%���T������w֤��0¡]�-������f�>�� Sg�������2~M&W�k[k�y��d����~� [Y'#��Мl�J�z@��g�|�A���сf���c�]������g���{��W�Ɵ��3��+���8rS%�)��i�lh-X�`�]�o��
�c��t֑���u��<��U����*������y?�_�ݓsk�lZFy�����m�Ӯ�L��j�-3�}��}MCJʴ��s�E��y>���j΋�+�'��PN�����N�߾�2j#�q������~"��gE���##�Z%��#�>��'���������:���H��	�	"� ��'F�C3�G2��>���}$��RE�����O�l���?�3鱚����BE	01�L��%�^�D{��Ϸ	=r�_�W�ٓWw,ge���8��|�<A���/k�U�F�`�A-4Q9�rZ�'��a������3�za��r#�T����Вv�PDq{3��z3��x�qu(��'iYr=u*��U_�$��D���v�����殕��b;A@Yn�������F|2���ճ�F u��ג�m`)=��JޛS��,X��o���u���z6��NI��i���������TɤԞ�&���>��ی���x��� ��U�I���f�ˎ��.Q��;p��Qb���\p�	;.��:����t��a��[��9��
$��l~�\�~����y�F�wG�}ۡN�W#�zI3K.lG앒��A��&J'���<��J�.��i7�O�'f]��������>�M�>;5���G��l���j�{u�F�5<�ᒺ`���������-���U�c_�[��gz?�q���/����f�|�|Q��!V{h���P1�����=�o�O�S�t|�b����6^����Gg���mz.���^�[�ŋ�w����S�\�ڹ�3�8���|8���#��7�}�����(�W�����s�����D8��=���z����8���ʏ�!�&�(��YKJ6�|��(�`o��|� ��`��m��Do-���ȿ�d�r�up���Ȫդ�aN>d|?������W�?J W.[��1��}tzT������)4�Bsc��)ѹ�~*�K�ɞ�o��3yb |�������i_�2�;N��':��,
�<��4�5[Z#> ��`*n�|\���r�N��p�N��H��Ϩ����5XTA�T�G��L`yxO�21P橬)h�v���O[���0[7�^頨�9.l��)�}�F�U�g�\_z��)u�o�T-�� ǓD���V�q���2�wl7.X�`�/��)��8�Z8�ѵk����),wY���J��8�qX�]���B1����A>����������ߎ]�#ں�̝]�g���W+�W�C����-9�B>��u��'Ƅ"_�2��rP 	�-��A;`E��[�	P��dK��ʣ���;-���3O���k�K�ǧ�8�Y��9|�����Â>�k=Iݯ��4M4���WZ�>�5�Z?�A���{��<�������E*M����������?�*63���V[����Z��KK~~���l�@%;#<?q��{��3�/�a��|�8�E5F���G|;�Sx�#y�F��?�]��	[���<4�lb�;L�y��G�'f����=��
$3N|��GY�����T�[�^�{������{兟�n���=������96*�]�u�+p�脩M;��k��M�*����\nk�:�� G��x8G.O>���r�N�C��XyG渕=���8䓜���y�^�!hwO>�
���-�~i4AygM�|m�s�1��F����B��+߶�gF����� ����W�w@��oど��	,UY�.���j|�&߂, 8Xt�Ʌ�{o��$1�Eiu�X!�e~� ��C}��C��������D�f�򞟂4���=Ogm�/�m,D�{��r.���H���B>�/r�e�﴿��6J������]�t0�o�h~�j����<�Ϥ�� {���������>Ч���c�[j,X��U�o���ei^+/�%е
]����2� �����y#X��7Ľ�n�:C���W�ޕ��J8t���ي��68�o�	t�{�����7Qo�K>���LA9�Ϛ���Y��]�AV>l���N��]�?�d�Rw�`>�dn�IDp�gSq��析T��Z��w��s:�:L�n��ʃ�G��2��Jɫ����n�}?�U�G{�Ǵ�o����s� �h����������*D�wlj�\���gNb���		>�2���z�V�q��q��p@��^���[��X'�e��ApЀ!.���t����P�Q�F8�c֞�YPF�'r�����9˛D�1 �ds՟E0>큏jL0N���xR�?�� 6��ۏ��S:�uS�o�o�!Kᾓ��U�o��4����^�����w�w4�Rv�.X�`�o�Oۿ�=�,*���<V6���/��m!U�9�0b�s�=��m�ɳ��޶d�Fp.-OT��@�}����4�3���O�y݃�0����E�����?���rtNv����D繃�	���+2_�R��~`�#��R�7�rﵭ�����i��E������_��S���!��ܘ��\��x��N@�����V���* �����j{;!��[���N>��:`�X(��;��4��~K�c�|a/����E�N�;���M�2P?�:����#�'�lsl�H�۽��׶�H���0����gd�h%���:��^���H��rx�`}�|�ʪ��/L��5�v�
�l����"�F�y��w�3jY��L������;�����c�ޅ!q�*���!�v?|��򔫭���8�=�~z��&1���w
��}��H>O���LHPk��M^o�72\mI#��Ʒl����ڢ���Ӈ��x��r��:�A>�����3 �֙(h���kۙvO=��f��غ�zE�dF���q�`�)K��H�9�iiǜ�T!Vױ�]�]���_������ќ��{��H��d�Y�����,ؾ�^�'�+�0����l+�,�L�o�:C���;���G���s�f���&(Q~G歛b��Ǽӛ8:��B!Y�[�EUǒW��f�͵'[�Eg�z��Y�~�jV��8j_��q+�I��r{����H��=;�ݾ�{����?a�:hZ7�mhk&���ؘؐ��^>�u>�u�\(;g������F3M��;��گ�k͓�|�i)O���S�6�v��m�!��د����g[�x��hoJ5�5�h�A�,�?4[�ryP|��~1��kҾ�T�����W_��k�y�ܭ�.��:�{�����d�����W߇���݄�o�d>=܂�Vlp�0T]�x�"ήN�ð�~��"L9�S��S�T�������z�M��"Ȧ�F�Qm����&/zh��
N��{N���QNc���7Esfؓy�uf�[�����٨#������@�o%grdOs|ލ�t � ��}��2j��ܤ�簮������	�ć7r��ك9`�����,W�����y���
{����ޞ�!m�G�i��m�b����Pm�G0�{������P>��}����6_W��.��AUa�/����vq�or�6J��xOq�A���{�LD|gNgy��9���+��� �+�T����G�$�eiM���-�*r���y'I��|�6ؘG�0������Lۦ.����o)��P����~��Lu[�R�a��8!��UU����q��%<�%%E6sc�wh-z�mP#�sZ�6�-������R^��(��T����(9��~=�`���^o�Ǿ>
E2d}< �'l]�2̻nCh:��X���^m�����.;����� 4���DQ�����D�+���Hd����� �L��$��"x�2�y�#�+{ >���D\����Ԧ!��#�P>�^h�[��ό|V>�b�t>�m?�;�t`\
��WŴ�������(�n;���KI�sہ�А�m�D�O���i��CK���>�>�Q�;��޿ը�?0�,X��/s��] ����<H�55�'��a�] ���	Utj���|�7�$�Y�6�c}y��>T:ڬ��O�}r�4����߯���5"�%>��Mi�m��;�V�`�y�vm${@+�w(�N���93ӕ�Aڑ|Q�Р\���/��Br(�dhS֬[(V��F��D�5��Ĳ}��n�����<�ۮ|��Sb9�z�zoQ�^�,��k�+�Q���%���I�{�e�43`��H���/����V��A��U��7��>A�Z�6~"�j!2��1�{��/�CH��Y%�)��|\[`�4�)Ŏ�����Tp.�q��2Bzm�_�W(�����^���}+ru�S�r���,eF@�'WRIW����'��ɡ��� u� }2�!� �H�Ͽ��,X�/�w�a����,��<q��:�>�����>�����Vd��31��㯕�4����p���d\w��L��𱾏}mI$�o�-�@�,.G|F���E�g?�a(�m+�oC�F�U���朠�ʿ�J�c�5��O��>��`��<Z�Vљۍ���Og �
��5�c��Wk��[&��f����(�7֨��}|@k�m�Ɓ,���� �I��`b�����ұ��� �Y�t��`�Gخ�s���=��rF>eO[!/��*.�π��/uf�e�ݱ�f��8�յ��܏>�˨B��pB��vj6���uM�#��t=ؑ����4�q��$ˇ�r��ه�%V�����d�w�޲xve?y��)��T�w���(�	وU'�?�F��p_ٵ�fL�W�Def��l�Y���<��� !,|ʋ?�2#�s�8�y2��wPnJ��*u"}}0�
��c��7]�eWz��²+p���,r��ʟqm7)"e��V�Hl���j�6w�vcI��{��m��u�O�"&�)�=y�}:g����P4�����wMI٭շ���}��.����X���_��mr�4���{�Ҍ��i���ɀ�1����JgB���!��sd�_����Ы�7ն����jf�Z���BA�VY�5�67Ȭ~�W ��<J�g����sC:��׈�v��
2��A��@��l	"b��u1�l/X�`�?�{i{�S٫��˶� �;%�D'�s�7���هJU�W%u6�w憌��|���*4�[$�����W0�D*���l��6�������q�u{8����u��8c��I�mY>�y�� ����߷Q�qv�%�{(g_���P>����J�N�e���-�pj��a����k���5����u��Z��߭l���{Q�୪���q���������t���^���������+TpR4N]��1K�Ϋ��^��q33Wo��[�t��gm�+�@�\�|G���Y�GyGy8p�2�k8�(�#�d�,��hMNP�0d	p9�A�'ߔ�V�z�[�^]Qi����n��W/׵�m�F�:~����9)�\`����5Ys+-J-� �UH��S�*�N0��h��u'��3'&ς�J�����,��~&~����@��c��'�^R��� mfߵ�`���fu���؇k��K��fIlׇY������b��&�oĚW��M�������z���O� �7�Iۼ֣ODQ�"���l��~�[ ��.�O�F!����+�}��4����)�CN���=Q���B����o �m�ݧa	�f�*:F��Wrf�$�R4�ydj�����]k������3��O�+�@q]�B�gsn�~l�l��s�J0��*�ǡȄ; ,X���j\�4�,��/8I>g{���]c��HDtv/���Íg���B]�q���y�hzy��/��2�ѽ3�{�����ߴ~��f��D�����8>��;�/y�����G��u�;t����V�����d��q�����1L�ZE����e��M�X���+��a�<�f�[݋����.���d�6e{?��*��]=�L{�BxCGw����쵼�oUHޱ���;pl�������ğ
� q���|�;N5Z�	jUȗ�F���G'��7��>��=yG�Gel�F|:#%����=)��]I`x��e\����L�������<�\���9�s�!�|�|�S�
pt����ő�i�� ��7f��Jz��W�dŀĠ���9o.$8lF<��t������$%$�M{Oa�:/3�J4��p8B�A��F���խ��{������4�������$���R���}G�U�ۮ^`���"�Z�$�����wj�[��2~��03�F��#��� �����A�·y�8�e���OA#Z�Ɏ|ٗ�����u�������0ό|x�>��5�O�vu7٬�e��[}�k��ʗ�σ2I��σO��'ŖIb?p6 7Z�/įTy��z?HቨT�=���@Ǘnj}�:y��� z���,�D��1O3�1l>��W޼�cv�uq���$���zlq.c������9�����p(�e�u�b�3�{�7�}�<��=o�Um{UM�%��m��i�X��]^˟Ў����� ���|�X��U�8�Ox�ϲ���'�6��D�ѵ�L�B�M���B٬?�Ƭ��i?Lƛ�:�b1�aD��W�E(X�whj}+�Z������#�XO<������>��'���WxͿ.���T���X��E:���`x*m���މ���)�'{�Z�}�8E�2�Cf����w�
�VLd8�H#:�i�{�G���G�g��Q�g���%s�i�TjcX�2(��4����Bfe���28�:�ُ��ԓwA�"%�M�a{P/C��/�=����%U��2��bJI��������L����ɸ�<�ਹPa3�n�o��+����:��A�H� {9Ĩ���w��Y�`�������U;30t���fs��$��~Ggϗ����4����<���p�޽J#�y�l�w@6]� 6���7L'�<t�}�� GG���H��2`~�B?Ŕ��R4���n��A����.���.>&����@���f�I)��Ayl��;\�=`�Lg��~��G�m8ȧ[�~��g������~�~;�:�Z|�z��۟J�on��-�����m�E#�MB|�)o������o����G1J/��X�����5�<����N���T���L���wzg��-�Z�gx+Z�N��y�i���n���fe�d���=?q�ǅ�1������/��0�Of"���&�4~O�Q�������@YU%d�I]��k��:?/=��b���u��|��#y�7�.>���,\iS>�R����9�p.�(��� �XW�;�*$�R� ��Z썓�,����8��>���n�Y&������h�)NKKhN�,m�L��y2@����y�:�sT�|N9�	})��zi�zD�骢��(C�� $���L�-҂YH�O��
���z"�,�ȱ={Jt�@���ť���5�qs���l�|�Q����̴`�����T�K�&�Y���I�B�j��n0��z�ۘ���R�Ϟ��;�3z��~9S��S*�����r��R;�"-d��O%��pXb$��X.��b��8�?�;�+��������ұb�S6��r��m�ψ�����3�ʐf�!s������:�i[SD���?��x��x@)��$����g%p�X��T���'g�A�W��e��OrE��d���3\]��$'��qA�f]ts��,�Y��N�5�E���1,z7E!Im>�|��݉�-�,۫'i�P��~{���ᥳD����~����O�;����6ʉ�5kԹ�m~�ڳ��sd��'�H>i,�]��|�9��XC\'�$���I+HjoDl�9�2M��=&���I��uU>P����F���9䎇��^����'�H�T�9R:����%/e���p�a�~׆Uyn<�Η��Oi���(�Q�³d+�%~���`~*�7����^{�g�D�g�Epx��I}:/�)Q����[c�d-����S�p���M������#���V�4)�j.g�h��g�V���L������� )�A�E���IY���(�5>��Z�U:��;��(�o�D�h-�6.��mw�>6�R!��j�<󒯩˹ �n����S��a�RglC
OhG��P)5�ء�`���1ц���w�����Y���QO�x^�N
�ޑ�ڣ��QKܐU����Y�����#��S�_��ю����d�C���gJ���ғD�D8NC��Ł@I�4x ��pC�� g���`?@��I�zq�����u�=h#���r*��C6}��.����fe�[���G��������;.)kdo�����ؽ3`���GO���'o��H����/Y�<y�A�C�����4��_~ �#����x/�H��,X��p��{�-|����<��z�Y���7��!?�+$�
i'z���Y|����>D>����rm1��M*e���d/��:N�ŉ@�ܩ}��C;q�/�~������^��dO>.a�`���e��8{���K���>�Fv�rd�Rۣ{���r��*����n�hYY�JKrC��5,U�S����#��|txq?	�7pP���:p��\�۠��2!�ڱ�;��N���?��HU�&n�_=�xڄ�+�Ńgݖ�J��W���������_���`����Y駡gd����)���c�^4����t�w��ю���K��q[)~����:'+�t0%:-��*%W��)� וCl����%g��<]�7�M�'�m ���*��v?¡^�X~{�aRn��²�h^�v;�!9rYCɛO��,"m 3���h=#" �q�|���z�k�7��nȌ�p}���;a�FVYˇ2�=6����|�7 Y�u��m;p(:����A�k���x$���0�����#Of�F܂~7x���]�}�A��'
��R�c[;��.OΦ�Ÿ�CE��~p|���zT�Rv���[s�T���������}�^)����-�_�}Z�η����������
�|����O�c��YYF��ɪ�g���J6!�t�3���l}#_d�w�:�K�����GZ���c�Y��	��p�����92�|���Y�N�wmK�rd�B���y�-�%Ֆ�TGy��S��LV��/U����r ��U8?��^��bdޓr�_]Cv&�T[;=�vr��Qn?x�n�-Rj��ꃦ/e� �l��ԯ{��� ���Yw��`V}�!7���!���e�,X�`�8s��ꗶ��>�[`��ͯz��<�5(;�������n=�"A�+���$t��(<x4n��m:k�{���A�3�eGe��������m{0�}A0��d�{�9�.�p�������G7��	_e�>X� ;A9�F#�L��� �I�WQ�gu}I������K��%Sn(�o�b�Y��:dU��������$��[E��>���V�f��z�ok�V�?:��{��/�Q�������գ�_�{F��9�~�Zwy��=�c.�B7�J,��%r�Nn0���..�y���D�v�.'���;�rX�|D�d�2x�~5�($�Q�-gG����Y!�%�#P����v��)��CF�3����*[G>Dy7�D���U�wP�:�.2zcLx�Β��F\��?�uS
�M�.Omsțks3cDkBtR;r�5�N%8 	��+#��c��8�('~�����$��Z�/�+�=m�`���Kx��!M����`�Ɓ~%e:P#�����H�]�j
#(.4}2�z�]�K���r'��;L:�ǂ=xq��y8K��X��x�-H����6l]�Hh)�³���Q>���á�̴�/��-.�a\��������z���d���]��=�ɑ�)�2�{$z6���5�ikbfp�Z��e�|��-��R���϶!�*N�sӴ�Vg���>[Ʈg����d��#u��H��3�V�Bϵov�0^�!���;�]�`����U[����ze����N��TS�J�U�hx��{N{tPffs��=���~π'?;v����O&)m]���SH�|��[<>NUE�������d�pRr�je���c�i�s�,�e�^����oI��}�%�e>��O��Cmb۴�
��2��}����ãx�I��st�lv϶;���1���뗾e�2�� �ƾ�I:����m�����t�CޅJ�$p:�o;%��Q��9���);�JFN�w�`=��G�=�yi��q���fV���샊P�*�y�q�v�yp�3|FFQ>;��^5x����Z�<H��2DtT���S��D-�b���Y}C�$�n���ˢL�X�`��*J��3I����Dg7O�88�"��T�ژ�J��2^�ݙ����+�,n��]؎'��k���I[r�Nʡ�a��ar�R�L�W亓Ƃ����#���!�eF�O��=צ� �U�s��Tk��6���:W����,���8
�Fe��?� �((�f&�v
u�H,b2��E���
�>������`.7\68 �M�f�d�|�����GQ��;���x~�H��r���'ۓ	$�I�P6�?| CK����4?��~i�T�
�ݛ�1�F5XF�f�[�,���~Bg���M;�f��]M�pU���j��m}�}��~C?�'��l���{M��5�~����tv�{������=e�Ӽk?�������Gg����w�$���)g���b�Y��H�|�~cZg���M#;܋IN9���"9��д�e��A;�1�9�U"�|�?��Ѱɒ�R�*�;�x5>���o#�ʔm^��S.���[���%"�����@ght��V�}���J��=��8�sh�·�r0�@�]:�lv�|Vf����`�%ч7��x3,c@@e�K�H�I��9�R��Kћ�_/@*�X5�^�S3ٳ��m!�����z�XIs��<�{�������sdw�K��nRvO>����O��TA�b��-�Y�ߩ~o7�u�+�쐅��*<��3Yװ*>���~�]�^,$U����h��+ކ�с�k��A�}y�k!�ۊ��`F��ވ�����S?���.o=@_=�y�,����#�U�Fk�~^�C�}�|i�gflxtg���'�����n������}S�t�E�
GtAr�7YG��$�W)X�g��?z�eD����3���nmpD�\�)[�Ҋp��'�p#��q�N� ��Xvr��r����'༶%SΓ�Ñ�a>��6i�W���6w� G�|��ʗ��1��'C��ϓ �HR�!2kss4��W�Mp �Z��[[-5�����@��G^�4��{[��OVz9�˱�<�
~���l�lǫ#/_���v��	#z˿�����%��9=����0�tҝB�<c8)G�W�m���p�vГ���y���e���-5�������y.��Ɏ���(d���/����^��4'��B?�&�F�n�v����Bx��D�?�{0�)���\JzLH�Rk�oZ�E�7��~�Wu��1�^p����+T�W��:�w$D0F�D≵M��*��Fu�=x����	�8|s4�l�rt��f��(�������2�u>�qҼ��'�_�SK�����H����)�`G8��9�A�s�\�g�Pv���2XYT~��I&;yO�ly8sd緯M�f����z����-97~��h����xH���K亚�g�s{��!�����ڷ�����|k%OU����LlՉ���!�.i������˂~�3z���k���<�����ɳ�S���A�K�',�M��=��]�w7w���`�>`S���@�L��u�s�R�h�����`e�Ő�fd�ӌm\�`�rf���Јǧ{�,��-.߄���cl$_�6j�@[.�����+�G�)��|��HJ�g���넍�gh�08��Ӟj�@(�'U?���C2���>���:D=@d����i�+\+~zv�w����%�@cT���j$`.���1�*8��G�줻�ɻ�0mc��5��8�k�u�׍�9��
)6Cη��͌A�N]�k2���kX����}�;*?J�3���(�p��և ���47�oh�,(Cg����½� �=i�iRv�E�C�Hvn���v�pt���)��_��?�!m�߿�Y�Ϩ�F@���|��~O������`t�9�� G����\��:��s���9��dƸ_�����F�U�Wi�T�'~2z��y�$�C��D����_y�\��Ɍ`OG�Y��'Ɏ�W��f:R�rqN*�#=�c��ٽ<X��K܀�pM�X�ڶå�����F�ݏ�Ҩ���ѰEg7����@��~�9w!�?�B��P����u��t��{E�j8���@�p�ݯ'��饼fΓUッ9�{�6U���%bz榓H��[�7�C3�N���s�y
��%�s��}03�F��YW�lgiFSw>���W�9�c"�<�b��yN������������&���Fn�O]�5
ogj�[�"- at�md�*p�?_���J�oW:_zhj�<�eT��D1~��rGX��U_�C��.�;Xwzi�W�Ƒ�$d���]�׳�2]��\�62�洟�CC|�����!1�ur��B%������Q�S8���B^���@�r4�q9Ab�sQ�G����n�ΚfIkB/[��x��-�?0{��m3o*��4��0�T�N瘁Q�df�h�W���B�u�7������~\�{bn�z�픥����P����s����E�$���$�o��b���R��,ڃ��g.�&�d犥#[��`�}�UT�(�͗�tg,��v��VD�ؒy�Ƃ�3}�����*�����2��ͮ��/�l�y;�k_����+j�(&���t��{�����:c�{��ݨ��k�N��zP̱!.��3��=���4���sl
Ύ 5��f6�x���F�y<�^��ɡ1�g�,�o[�6���	�f��+��Dʉ}~�a��.��R8�<j�L}k�kEO�X��v���������谚��[+�������SL�}>����«�T���|yO��w���輿v��]�W�y��8�����/�{u`_�v�G �Q��(��3,��g�Q�,
b=XKs�8��aT��h��\K�y=��1�G'�9�s�'�i�A�vudw�y����?8�y}D����Ti�O	��$m�9R�ke���,� 6���:��&ݽ�v}�T+@`&�A��P�(RB��宇:�8�690��@z�*�O��
���>���ٯJ�L乂��ϔ��c|xx�@X9Q��������7X2�� R���HP$��Sg�xdG���S	M#,{�n��p���s��P�\���x m	yip&F������� f+����	ƫ��|7���Vi��GF�e'?�0�s$ӯ����-!�'��n��1��U��]y\��&�<�!���X����!ro�;z����^�( �A���j˱o99�'�.c@�d�=V^��B��</~Q=���{������M;*7K�J�Y�G�붲9�>pZ��7�?�1��>~�ع�?��1~�~��������ai�~B�~�O? �`f�<|���Q�n�g�EY+s�}�]�m�����1��7�_ppV>��j"��|��/�3'�M��D����&�݇�m�M��e�"�|,�Mk�f��T�MFs�I���ڭ��  ��IDAT�q%6�����$�t.� g��]G��0=|���Z�!�o���7p��(7�ց�'}�'X/$w��{kv�N1
�H���A��B-�J�k��`�|G��2D����2�z�Hv:���6;��@v���|P/4�PUgS%�����h�ۆ�.�__�U�Ɵ�=�L-zF��̨�R�嫍��4�ީ;n_W���מ���p޿��� ���b;z�〠5��P˓�_����Ղ~^q>���D�ԓ:���ٛ�c���@Y'�^�tW����(�A��t{��Ɇ��a�k2xӫ���� �)�6�LN�y����}<��i\~�#��u��6T�'�U���)|*&9-bNH���y�SS����#ڐ�� �����5��U���r�K�6^�P;�Bm���+�u=��c��e,8�5o�W��ͫs1����ߵ2�o���ě��~�7�ݳ/�3a�N�c�cv�'�8��.�����8/2��b��gO;�����3ܽ���|�^̄�o�v�s�~������ݎů����Ӿ@h���6!�nF�q#"�亂D=e��F([G�����w�;���R�9�'p��_���@$��O4�1�f��5 V��,�ɤePv��Z�p~|r��3�C��@����vR8Tx���|�N>A>[.��l{�W/%C�oo� �.01�i5<wt�@��#A�#>L19y��е��i� ��`O�������VMA����.�7rо�0z��}��`��	�'���7jۀ�2�+��Vx>:O_�o�}�o'�cm�QP]�����#���)��&06����r�g�iR���|��{pI����������N��GP�Rj8�l�������C�C{5���T��ڕ�Vu��\_�lm�s��<q��+��GW��|�g��ս���xg��gH���Z[�n3����r/�=�!��^�}��,�V[��<|伩�����s�L������1�.F�.�����p �>f�n��}�k����x�XX�Ӕm��{ZB;��}km���4NU�1~g�[:� �d0�O$�p*>�mC��^�|jjy���/�q�v[)h��f0�RB@;��<F7ѓ���g�؏T��&��xXw��#:#��uo �ү։�?\�7t�:��Sh�plr���Q�}׮�ͳ|��}��G[#�)������#`����o���C�U��������6*�Lrb0N�A���N����5HP����.[��C�;*{X$��o+{r�5j�O�vDZD��)ȍa���d�@�dc���1�<���a����k�k����#t|=��s��bh=t�z�7s��(�wմ>�]��S�
����{/t.�9��_9������[#Q�6j��a��Иl�E�����){���L"n�'�������/��Чi2m���U����E��6�̞�rM�]�ϛsW���e2Hj��'����o߷����\e���޵)�W�6t���s+�Ɓ��:�l|�>��JX�b�bֿ���f��V���n���!��Cҟ�U�O��o�Fm�����J6��Sڠi��ர0j��!-��|:_1��S���)p�2�M�x����xC��Z��{<��:�����'���lr��z�7��v��j��:8�ג����o2�j��ˉ���V=������e�굽�.,���_�z}e�F�m�|ilS��]�$�~7����˶���o�ӳ�H'�Xcok��U]Q���y|�}�kW�%�M������[ԕ?�C������ֿ�<���/�:��g W�W}F�I�^��m��k0���^{p��Hq7��Mi�����n½��΍F��ƶ�<>X����:w�E���q��3��B�Fg��l���q��|���g�a�?�ɬ7�3��axE7Z������ڨ�<�6/�/1�fxyz~��5��x�#�h�`AQ�<��Z=�s4O�@�"��7���*Τ��3��}OA��h|�x᩶}߂��x��}m >}���F��<�+l򳎊�����<��w'�m�(@!i��N��A9�2��ӵG����t��M{��7���O�A	h�����6�?JzRƂ
&E�Ņ>������=��Ѭ�K�DZ��n���V�Z���ۗ�-3
������]1o�۶���pN4���!��Ws��Ir��uiۤ�L�S��;z��W�o�=k�>�1.q�l��vL@��������TӁI!���"��=���Nݲ��)�yv�䇠W�'2�#��7#;�Ҕ��Sm4,7���]��k��� x���|��U��P�����n�do��}�n�"Όt��zy�����>I{�M�(���_��{-��<pA
Ruɭ��j����,�<}��z�����{�6}�@)�Z���3���$�!�꧔C�[�
,��Յ���*a�c}��w�=�~�{�/WCPn���=R�����ee�P�N��`ˊ-�tl����p�\����Α����BD���lG��p�㈏�M�9�cib��~FF�/�̶=���(��i=�ћ�G.��}z�Hm�pd>=����s�{(��Cb�@�Q�����]Ա\W�q[��j���>V��N=�
`.�9i��x௵>�P0��zX����J��+N:�e��O�جC����JO���V41���kK�KN�-.9|@O�38��^ov|\�m�lwg�v�g��g����(��1��j��
��5������\����W y���O�J�UHW�#���ȕ�%�:4NoX�:�E��{p�r�H�H���]�I��'3rb�(��:'�1��{Sm��_������j�H�����PT�����>���I��.h�����o�Q��sc�����C���h�ДTH��&ا�P��%��;�-�����\0RG�087){6��$��+Mv��#�WnD��|��B��7�ׄ������,ɼlƐ��I�}����8���$��FR���N����{��Z�4�'ɭL{��s/����u'�x�Hr��s��r_2�vB�ܥS�Eܧ���o��y�[���z��ߗ�u�n֫g�*z���>�+7-��@r��-�{R�p�/j�	gA�S�>i��t���P��w����&w�G���)m��?v��x<g�p�(���<�e [.��*.�����T����uu6�;�ڶ��	N_���~���7���5܃1��?R3��l��n
`�3s?:Xa��CQ��OZ�E8�^>��p�	� p ʓ�ʃdd��*~���3����^�3�\�gT6�X�F4;:�}A
>a-���.�d�C`"]h��*LN�����Ω�-�Ё|����LQ�v?���3a;$�����C4J#~hXf���ʀ��NP9	�2��)XN����)�mԍ���qqv�+v��~��(M�����7n7��>vV�������D��K���=ѲD"$�.lPD��9n#&h)��#�,X��aňJ�M�}	���7���[�n�ƀW������	
��er:vP�=�~�A^˫	��r�C�[�'�~W����2���WŤI.#������qJ��詃b�1����u>�y��=�,����wp�eP~�椤uN�+���>%��	ա��AR������&!�۔t[H�<���\4����*��� o��b-#ر�S|_~�c�w�r����]��)L�Yͨ�H��y��9��-r����&�4��J�`��r�gcF7�f�e�8�ծ��lR��n��|�
��ۿ̃[[{<_���͎ �'�������i{�g�{������l��;�oVv:�a{�pa;��v '���)���q��B��J�~E�G$[6�n�PG�H}���q-��,�nK��J>��֢�jdL�uG>����S�������.����S��/��4��Gv���%��T���� ��ST�((0:x3sx�Cf�(���r�'۹ �+=.�6f��2)^�aAg#c"�:N���bc�py�#�H���=C�u圶��3�R����rV�d�C9�r2�TO;Yi�R�#�41_��0�X�O��V!2��Jsۧ�`s��؊6A��qxe׉R�Hu��>80{��`�P��^s�f��v��#�w�>��N�=}�gn㥬7���cvm}�k��������ld�/X�`��J9���u&c�i#�/�N�6�!)h���؞��C51�ĳ����깞G��=�Ph�x��F����;ц���	m�`�X�"9ij�_��>�WD��A�l�FT�'dT��X3�;;�sp�8�&�?�X��y��O����-{�4�������ܹ�X|,�ٛ��=�l=2���[�mJ$����瑺rp�'��9N����0�w�E�f�yd��|��C�e�%|��4�|0P2v�"}��kAK�OnOY�>����O�Fby���Yȣ�|�|.���=x�Gk˺�x�d1^��-���[���7�«���4G�/���j7t�g�T6���6&��,Z����)���G��
(ǳ�A���[f�,fdW�M[�<�s64O�>�U�O9�3��ʐM9�?"{0�nz=�_���i���>�k���q�tz�vVM�<g����+�(���0���p� �Ƨ�C�%]>>0�����=����j���#ՠV}Z�"�fBˤz������\("�6��b7{��y���Dp�����Ƞ(,�3h4#\j8V�J!%����p��t��7�)�-�H>[�pJC3dϑF���C?"G�[Ƙ��D��}�A}z�>�i�'M�6���\%�eS�I{9�i���W���,Ù���7�������iP6���~�B�3�7Ԥ]�ɫN�P�3���3�f�@L���L��p*':B������~�k��F��c/��(�'y�7���^㲏A��~��`���^͞�I��M��Y7�9�5]р����h<X����薒���Rx��O�v{��Gݺ)�\tT�����Ro�r���6�N'�eL���>��@�=d��k睧s7oh?y�@l,�j81"��D��e_Fn� ;;C��5Ѭ($E��K�lp4(7t��b���>�ݭ� L�)v �P�~J@��e�ie3���j��V�ܐP�"0 MD��O��a��4�-�9����A|�l�3��Xۜ�ù5cp(�0��^���a��/jd+�#�C�$^��-|�=dRʕ����Q}�=���R�<����+u���+�y��Kq��U��F�8;��#K���� �Wf����h/��E'�|q���KL�蜧�I�s:���l�j��f��+ll�������[����S����jP����_g!�I�+��G�PLs(h]���H���̐�Ñ��.�	\�g��q�S�
d��o�p�e�`��#Γ�L9;f�8%!�$���N#�����(�0{y�*�g��8ή��8N1�oc}�{\9rR2�~�/��}��˶�Yq|���9u��T�ٵ�ey���m FO�' �A�+�2�1��#F�'O$-Hҋ�]�!9*f�Φ<@��R��iR
G�H<pJ���G�����zp{���\�*u�^��=>dd�|T/%����=�ɴ����B���c������	"���F_�.߀�2hl������ѡ9�ɮ_��.����>e�;��Z�f�z֑�LުSr�i��(�[tE��@�2XA����:�l6���f|l:K�!�Tx���j�,�����M*YTQg�x�l9O�f-���w���m��%8��z������"_G��y�l$̒!��mě"ho#قKb� ��4m�s�A�(D��n�k~�Ig�n�u��u�L[v��^}�6��(B׶P.�3���h�EN�R׿
��[�<�.'A̬�
��ʗj;+qj���5)��D�6�r�@�tn���A~4���_�:xvM��T���5��vʂ�}�ľM~��ƃ.�<�A�Uo��1�,~g��*��u�ւ|Dq��^;tX�MeHt3�+��nEG�̃�j�xUyYػbK��/�O�@�%�T"��a�net}�Y8p�F:SҌi�'� �{\d�v�q���۹|R_�)��|#\';�䷟�����=n!�ʍd��@�',{>�cxH}�����^�l�&��p��R��>cŐ�T�ץ�
�0����}�����FA� 9c�,�:����sz�}2|�*�le�e�o�]�2o�M2`����y���	ѫ�h2o��C^���a�3iG��|��Ѣ�2
�m�Ws����k.��|(�������G������ +C;$�r�uN4n�N����H�i�b-:�h\�+3��9��_6o;KP�yT�2�l����OfY�!����&�L0n��h�P���X�k��5��br��A*�'���B��!�޹����\m\�"��Ju���T��6��
p�Zg���qK�R����&�~�ayL��A��bi�|��ʺ~[���i��C �'�0��~/�a<��Ɖ|��g4������}�̊�����-?�Y����'�(��O��c1�g�̭.��J�n�PA��W�V���h8��Z�/��A��:{8&�����M9���q �� ���̋������5D��� �2�H|j ��(Yj�U=�5{57gHƕ��
�!z���� W|@�Y'�C�����<{u�����ys���a��z�?�ݣa�5���ݾȈk��y�B���5�w���c�������/z�XI��{`�.�*�6i��+��5�?'͵#,��O����0*G~�����~��G�~j�%���e�qT�ۋ�rd��H�S_��G�ޝ�����i�?����
e��e��]S��n��9�,����8�cfd{r�9�m32�[� �W�MH��_C��*=ڼ�0�l�m���:Kc/3K�� �`��PONw,��{$?�)��<%"�Mç�0�}
��qd��:Y���Q@q"ȉ�l9W��:{4C���8�'�6��N0#�7f���+�X���O�qp����?T�����K�i���uDh�3h��hB���TH�
��������8��qv���w������YB��H5ѤD�]�h[���=I��s{e�37�]f�Vں��q�i� r�S*�in]��[O�e�.X����-oGg���n7�u�㵔7�ҡĞ5��DJ�.���}�I��>��D�ڗ�hZَ6]���-�>���I�=Q�@���>2��[%�.���&��2%HS_�xu\�j�5;x({&Hi4;#ܤ)� kٕ|��<�AU�Ƀ/c���?�iw�������* c���wHL�6:��}�e���H��C��/Ы��v޻7�կ&~�C��.�\�e�������2�������=Ƞ:��qs�#�g�({j}���\I�V�D�`�V p�GKd$��$�f����mx�/�*2��_zh��ů�}����3�揬k�^��F��'��t��/Ȼs;9ج-r�=���������b�)���7��wB�Ao_b����l�}	lF[W�^�i�c,��ϡ���u����DC>N�u��uu���x y�콃���g �1�qZ������pb�F��~Jo�~�?���^��/[��35�'��2�� <��H�j�����g�w��jo�=�So�������Y���eB7�7��>�1���Wh8���'�3=�S������&�7��?��y��r��tpO>G�ԋ�)q���J�����6xm�L��?#������:pQڰm�>B��i�:��HΪڷ0�l5�1��]a��"Oj<tdS�e�6���ONI��ö?�@��(ڄ��ko��6&�IS/��kŬS����~����a(c���T���<�@{dy��=7��AAᔧ��(����}l�z���ʕ��B㹽~��%sk�g�`���T_{�l���:~ŀ�>��][� ��+zt���X��,tvԋ�zh�`f][�����b�`�g���g���Q�A�z��v��(��*6M�5����2PGςۥ�Bly��y������\��7M�véV��ߤ@_�-^u�n�M���~�ȱ�h{~̈��ϣ=�du�$;��C�2�t��yfP;��(�l+g�h�u���_�Y�g[��l+�v���E���\v(��ܵ�*Pٚ������.
��� J����{:ڎA�'!0v��T�5ӕ��t���B�x�l�)������C�LY�ʑ#|�O�����r������������0�߱L\�{�*��r ޓ�o���<���[���+�7lP��p;0�m���$�q*���o��_��ְ���h��f�L��Av�7�2ދǍfn8E
p���R��1?)�=:�b����W����\p���i�Yt�J�Z��錚	<|�y[�Nc�b�#r�4�zBm�A_^�� ���|
��6�
5�|"H_���w���7dC��I)y~��B�l�h#�͉�\;�._���v��������YD��4�)hB� g�Ŵ=��/�ї�ڥcӽ�	�.O�F�oq����eI����|���&����V�P7��Y�s����������X���%�=p������%_/�{[O&���p� i�%*��g��9M��&�NP�Aβ�ga�W3:�Y�0��Az�a���c�=��nQ9�m������8,���T��)�L�L��ZR#	q�PvJF�[���t���~��t���:>$�:kg�g��]�2eģx���K�G��*r3���e�w�CPJh��"0+�>5�U+�@=O0���9�E6$��Mh_be�d&�F��#dV�}��x����[9i�˰�
��5��A��y(�){��n�w��R6i��Q7o�����hf�m�B'"�)��#�����\p��aEV����7�LV���$��I�!�-`v6��/��%6kڹ�-zh�&�3~�YX�	��&�maFD}y��e�`�����q�gv!d��YG����6;��Rh�J�H3�*iT�Hi�!���у�C u˶3~]�j[�yh�!i�\�vg� (�W<�#y�r�f_j�`h��Z񓌡�kqO�߲��4s�pN�W��P��'��mh�0�/�H�Ud&�>�����f��s,+�d��F��A���ؽYoo���P�Áb��43P�M3�6ZeE�%lu��'�;��54�K u�N��gT�w�/���>�<&K*^>Jܱ�����ś�j��ү����a��;!M��K�8�=���'1�Az���B��j���ۏ�vіP|����څ��h[�W�l�DsYl`���Ri�Dg�����f�,О�eK�+Oc>�4��@Ì����N�1��8�����]����F��"Icj�
=0oT��Z����Nm�����9ѥ��q�{�/xx}��!��0�h�y/^!8T�%x��BHt`��>�w��}�(9�p�ą^�b;~G��l%�*l�󦎯��s�V���i�q���ZGTN����mRה�.4y���+�Y����8��� ��ۃ�N���h/��y#xF_d��VנҐ՛�C��m)o� Δ��).���'�lz�T�j��NVbk;�^��d�U�t�a���d|ڱl�abj=v�3R����a���� �J�t�yt�(���PMN>�֗��2�����'���8G�'G�ù��IZ�Ѫk�'�[M�.����1�O;l���<t���Mj���'�x<ƃyUm���:@R�s�a�!�79����d�����=~쵵W~`5�m'�I54���\b7��y�;��E���#���n�}�+y��,-��ꁯ�/���P5E�"���d;�a���/�˝���;~�ی�	�|��쓭Na{�M6�S� ��'���y�v� ��I;qCu�j�j_12�E|�2O�ї��k_��TF�CF�����/�{O/���
���.��_��Byh����4=�I �����n!O��5ܨ�Ɜ�ߍ�@P�{}A�X\K�/�?��	���i^B߬��~P�'�H_ǈAydi���Kpr�	����}.��.)�4��Ly��M�Jy����E�`���0������z�k�$cҾ��<<�L�8y��2�>����:r��w��7�7xE?�ό����nZ��z��C����a�Ѭ��qO��=1"Wz�x)�0��k1FϠ��q9�ż�뙒��b�v]��)�}�<��-����Q��7�C�{���i@�9��hЊI�#}�<���5"��p��P�:�+�M�h[�bV]�7u �x���1�k��(��0:p1R�+֦��]f���L;u���n>��h7p���������Ͻ�q=L��l�)2�P�l�z0��	��0����}��՞�1���X\p��,dz`�	uJ�rŹ����6�����f��7Y}�ޓ*���߼;��s+<���]����<�п���͙.rA_���T�գ3C�N�5BL�r��ev� �\3BݭvT�����֡����h�29>-��-��e�����A�����L������Z�;y��y[;ԓG��		�<�\n��Ƌ��P|�?e�a�#�oI)T����,t����E_b䟌�2Ge��a�� X㱄br[���_��NW �ĵ���9���2$Z`���Y:�w���3#{�yT�.��$��= ��?���D�Ե�@Gmi���,x��oT]��H݆��q��w(�#+�t�IW�bF��� \<���2�Nވ�b�vB�9���}s�{L@�n=�!䩩�e�>G��L��z���ɽ$3�B?���h	�����P�#�l`�0�tn��X��柰�W�/�l8v�C"b4wv�i�Y����W@��>�9HpYV�́�v���3[ ӨI�x֨���Y y�;�򛞷Ed��%*ʨP�/26����Ƒ�����A^��D�IZV/楸���_���bT�WJ_y�>���w,��"�}ft��ĺ|)��W�;���O\��k�n��d��ɤ�[u�g�ς��M�=���~���:gڵ�P��L�ޚ�͎����{}�}{:Lh��}�ﷶ��P#�+�i�QTL6��xбm�mF��<�E�WB��Hw�4UBb�r�\P�_]��{OB�m��}	�F4ݔ��^� �GY��$�Q��G�t�����\����aX���ME�k/�<��G��Ԟp6U��S�B�զ��P���cu����T�X����=l��Jԩt������6kU��w����O��׷>ǵ�.}r��L	���BY��c������u�������}ɘS+��p���i�y�.����^G}��`��ǥl���9��;ȧ���A�N�oVb.�������D���R�Ur�5��j�+'>�PB}-y-�����Q׹iug�������=�ʮ�B\p�{v%�������X�7���[j3�|���a�ٻ��l^��u/�l��7l(�v��8�C<��M��d6�s! ��pA�N�5�iC�e�yڵ9Nh�q;Β\�_	}�7�2څ����>hإ/���Y��F���H鬤���t&�G0_�T��`����|�o�VE&��Tή�g�~��R~0�}� Ǎn�������b��c����\ŽG9�P��3OcI�ʗ.�m����Sr�G����ڮ���-��Sq���*B"`�Ư*�#���墎"�7nf�����5F�,�ѵť��O�Q��rU�8��s~+e*Yy�]�˥{(I�s ��~G%/�p���m�R�7A`�a^F'*����Ӽe7@#�X1F�(��	���"�h�
ogy8��	�쫈*-���m�s����f�Q�F���yܤ2�>�?,����'pg���ɒQ�2+c���)B&+GNlvm$�n�$X��zJ\��O������:��:��}���^n�ܩ��>�wK����6`��!s�n<�e�}���OT��Ny�8�������yʤ8̪kcy�cԏ%0e+p�BYE)���Tp��&�G����Ʊ�6	�^p��!@�7اh��1���d��d)�KW�Rot�����N�������÷��D}��ŵO��~�|{����������s"��-��J�o�8���W�C�P�T�{�ov����Y��L�K���/V6���X����4QS�rHB����au����F�g":��CT'&O���{�#8�����.M��hh#�������ۤ�6��`����y���׏��-i2����f�L�"�Ty�+�!�a��8�NpS��u���ydM�TYsrPٮ�B�D&\C���3�/�~p�O�b�6I�V����`���?`�������������n�@te���0�A�=[�í����C�1J��\� �*��}��G�������r8Cd�mc��h>����G]#���==N��W�3���o���� ���l-���˂t�\P�t�O� u�LG���H�?>���Lw�[��-�+��.��{�6{��o�M�������4>��L_��|ЉͿJYPS���ݥzw�}�mҪ}���s�ϩ�*AZ�lW���M�����
�"Wf6��y�Я��h����f������}��_S��h�^Bs��Qs�J��QU��i}>(����:�GF'���,�����Il�����,t�ނ&s�o�H���9H���yPc���sy~�[��L[�pp�������3�p�Y��D!a��ޣMb��@�;l#�-��D=N���~_�c�����SU~�nО놾}��ۯ#�p�xk��񢦃�ePMӚ"n�"ĖAq����8!O�qW/)�͆�-��2�w��2�{)o3\��;��{҇�G�}�\k����$)6�◵X��VN��������O rF}o@�o�-Dc_��6P�ʦQ�3�l��J��R��r�'����/2>� �1�}������-<�����������r::ڗ�=�ݞ8�jG���\�_�L��S�|)e_�d�bZ�I���v�k�F��	��״��5{���~�+nu�^�U<�@_׺�_p��^	S�"�A���h|7�bz��Y���JڵI�m�~��C!M�w�|�oQ���ͮdˈO��=��e�"�'8�|����<�9-���'=�I�Ox�����t���nt��'+=G�/]���p��m��@c�!����6�ҍ��*|�2�lb�M�FL�3ȫ����������^�}/�-L�}^�N�"-��_vU6���h�Ǎ@���Y�[���0e��)�?��1�#�$I��{z��.������3-�l�����~�V?�Q�ܭ�J��}o��
ݠ�q�_d�}���`jc�����W�y^�5�O06���<�������1�ٸk���+I�"�t/�ޮ�p6o�g���M��7tJ��	�I����&��=8]��4_2Z'�C��^H<&.3R�X͓Bfe?���� z����O�C8��/l����Ifd���bS����l<�>v��*�Nj��$)�����bk_k{s-;<5U��Nȣc/��<��i��O�F�ۡ9?=������%�CW��.1�R�i5�}�f�~Q�7�o��#|\*��/�%����N�nڌ��>]�C���B��Q�b#�l�}?��_X6K0s��B��� 6�7�d��̪TS����bF�vن޾Ac="���r��$}̗���6�س��QM����t����a�Yެ��x�0�^z�y��^v�`�����Z
;=v�~Q�` ^�F���aW9,�w;a]Ƭ͢�n���*#�}������j*XF��o{�DoYX}<4�
�<�]�N��IA	
�Ƣ8	�טd�mɖ��1����;7�&� D�ǄF�BM��r+ק��վ�7ht.Ї�WU�`�$�d�Y��7;�m|�@��f�;O��M�A�����!�S�/�t혉��8N+��G�z���l���,ukb@��g��m��Z�<"i�mH����
2�@��)f_{0���P���%̯��n��z����#�A�7������(�}�1��.J�_�pP�]<���>?c��Wِ\��0ZW�R�ǲfx�0᪯�E��WQ�?�C�����=D�����6{���]�.�������'�#h~RU��σ�������e�{��2j��=�\�y�vh���桍9��<���K��#	<ʛ�3�;-җtvX��<R�~�%=�!��I��I�w���<U��P_�y�&u╘��n=���6��fX^+���	?�(�X���[�񙍵�S������hέ��g� �,i����X�i8G� y0�g�Osγ�]7|����f(�0�!S�ʭ��1"<���M�I���^^F��Ay���o�bǂp�j*dP��'G�����z�&8;��	������Ǳ��'�t���)�%>MV�� �N� �C�ᠴ�K��ZG�������n��9�`j�����J�J#P�֠�\�O�8�S�-��XT �gX�6��W�+#e�m4��c�5���������\p�o�n}P�=��R�G�[�%[S��Y�/^��f�2~m�����3�Y����*�-)[H��^n:����E�շ)�R�ӑ��"�JD��Ъ�K<��l���NU5+�����[�����a���ʘذ��g��Kݒ�v#6@��A^�ގ���1��p���XDA��G�!o�������7p�@Y�0&�ϸ�����ً��n��	r7kT�4�6�d�ZI�y����Su��@��>��V�"m��f{7�C!FG�Hw#���_�3⽡���t�U��ǵ�iiz�*���0![I!�[�0�6>���ĸ����ӗM�s��<3w2[o������u4._��g��(&�eFme�g�P��P[lr��_#:�a�}:_�9{ ���>^GE�Ty�<��x�޼�P�sq�=�Q1�sK�'+\�<N��=H����h�B���?Σ$��~��;y�fy���4ty��Y� �L4R�퍸JQ/��):hg��B�SI�H��ڴ:H�1�<ηh��{� �ռ3�������� G�;��Ä�/���4��j����N��Z�����-0��l�=>�~<�v������=^��c�u��_U�E���Lzj��?S#2;���J�ҳS��\ �JS}/�
h��C�H}��%��n2� de�����Dcο>u�@��I*�A�ki�c�<�q^��i_��Nt�30�|���/�{�ώ��2��)W79Z>n0_7���h2�&�I�@#>�'��2��<ǌԈz3̔3��Fϊ2G���Wo�����z7���C��6=q�A�����Ga�t"ԏ�v�F�gQ�Td���ٚ�� �]v���<Ț�3zP��En�z�Y^�Ol�Jqc��ٸ�&�D�o췾�z� ���O���=*�e3�*���XYSY01ýл��!{�v�G���`yrm�������q��w\\�x�ƞ6���!��.�ӽj����_b=߱� ��y5����:��Ki��y?��D��m�����7C5Gh�s��ڱq�c+4�U�������i�6��Y(H�������>�; ;4m���*�0an�tgg��]���$�\
�f���3�K���_�yd����'�,ϋ|W!��»-H�hl���i�����k^�"����%]˙��GcJ�6���Nl7jt1��|��T������L�3�ێ|��K��Ug���{��o"8��V�&��A��B2��?���у�?寢)��ZTt0��!�_|u�:��f'�M�����۔1��x����e�aٳ��z�N�6#�)��e^����s0���܏��l�U�3P}�� �%�$����\ks->�rtf;��?q<VPV&��qX
C�]u\ѐ�30�G}��v����:���R �9�ņJl�n�b@,�;�oS�(��<�gW�i��>�/LO�˨x6����=�/�!-y�~'�f4�JO_g�:��QH�������}�0�MF�Jɣ|S#�5&��3�ٜʇ�E�ߣc6�軲�ϳ��;�9�ضѡ-�ߧ�C8�!����0��	u�O��Z�0��y�;Q���}>.���/i�mb��2�7�ܳ���;H�ۀ_�������(4��A+��<J�%xy�b���A'��zŧ��b���|Z��EƏY�v�Ny�a^)k���V�$�eK�*P[gU?؍k�/v�v���o���}���ڱ���fA��FC�}{b�r��#e:�k��iF[�����JxͰo%o3N�؏�s��!?��[�~���:Xq��Y��s div�0���f�^��ʑ�g���� o}��/�x���]�7��4�a-��'�K��Ix7��t�X�:��:�{$�͡s��4�?��}Ғ����>�k��2��{3>�:`�Lj�rʂ�zܥ��٣aV/+3�ùkϊ�W��敄�������Tla%~JvoB��V֨�U����&��,S��iѾK�Њ<�&DJ��g�Td���nU�غ�dDA2<I�|� �4?�����
.b/:��CF�	*M.�;k�
'�C(����Rd���(����a�i��2Ĺ�|�`{�k�;��?-�=�򙚝��5Cۿ���;���x��?\�������c�I��Zf>��)���*<��o��[���z���F��h�`�AV�.~F�&ҐU�q�l�E�㤼����a��?;&�p�O����J��h/	og�?���ȏU�v�E~�4��|TKL�ϻ�+ɂb"k���Z�`��<H{�cF�2����}[w�&��Y?����c�x�ؓ�ao��d~�;#s�T
�`����?�8�a��1"�9��9�&���m�eY�\,�	��ea����ŗBfĤ������S(�6�q
EP�tr���Ő�)�P�}����z�~��>�i%�s��> \���{����h ��0ߓ>L�ǀ�Cf����r��V��a#���L�4��2͕w��W���}_�c��"x�@EiG�%9g�v`�{{��M��ɰmά<��*p��9zbPO�~�$���.� uzjA�*�ɰ�J'ʉ~��S�Aλ�SI��r���ˑ�DZ�er`�D�=_�g�eʑ��O��5�zxjc�輏�q"P�n�a��4V%�W��\�tƜ5 h�6�T�p�अ��L]9���8�	�Y��|梇�v7�n>�|�B�%��}����Oa��(~~p�@���W{��e�n�P�[>��]��oXwb�5y�V9�����i�r&�����|�ق���#��8U/ɓ��ݶ�bev����1x�����P�DuW���]�7.��� �p����Ę�*qD���uxB7E�$�#����?����FOd"f��Hyш��	���=f_��g{��������_�=�.���"��}$�o���	o�{Y�Ƌ����v��Y�0�B��ǌ%�q�}+�G�3�G�7jy�F�wbeU��u�����8k�?�Ω��Cp� ǌ1��F7U|8���1��nO	�!Kw@��!��|l���GN0�b=�D�+������Ⳑi��w�����W% 
�(�E��6<	�4$i{4�~v��"�:zv�JtJ_�3��h�r{������x�ͣ�i@;|��7��Xv0��
��AC����&��Ѥ���('��*�"�9�?�$��͜5��u�;˪t��i�����젟޻��i7��:�W�.�`�'�h;n��8��?]��0���0�xOX0���H�k{H���l�g!G�������U
%���˘<1�0ij�� �
q+�ct�Vˏ��;Y�pVpf�맬���
����2��	v9�5����|�<�9�����"}��s���g���o��>G�Y<��>�9���/n��Ǜ<��'6�Cc���	�l����<زI|��&���U��r�a���d'�r�B����8��]��|/|I���y�����P&f,�e �?)����9��NfF����a\]��Ť�}@>�K|�%�(�!�8fye�<*�B{Y_ӽ"���~K���=l�&�e�!oCb�;�O|�א���#�c��҃��9]�b��Z�I��MWݢ|�����lG��V��O������i`+�N�K�8��4r��	��x� 7.C��љ���֋%wH���x2�;�6�R�4Avr|P�a2�`Q�ԃ��� �1O�	c����`ğ��,��e�^G߀�Y�W�x����ƛ)?h��2������6�q�o҇���9̭}z&��z:�ZE�2ۓf�p<����TC���5B���Y�b7 g�⑫a��#�G���O=��6�d�����_͸�� L�qBL��_34W�+�p�&x�f�K{�罰d�.��Ï\p��W���^����oy/��q-"�E��1wH*���t[�0ܚ�7��h)�[��&r]� ��Ũ���&�u͠{���I·���3>>�'j�	��ߍ���Y���W��N?Rۖ}�����0k0#j捌p�����I�s���y�Jr��X>�ʮF�w�J/��<E�Q���m!�؋�rC�Ca�b&��7?[���v�/�5q1[^�����ϙ�1��MK?�Y�^59 Ot��|Dj>����h�?k����<��e�	�u#~٧����i�8�G�m2�ܬ�m�~��x�Mw�|؍�y�/G��'Z��m��׷��$�>������!���E S��$�����<�E=��?�t�{1�Y^9�i��,�%<J����0`.�А��Ч�bF{I�i��r�e�F@���\��V��=qc}�2�n��@(/�	��	k&�?���6v�K����W���3�=��%M�z���)�'9�Z �w�������I�۝ʟ�}L����넂#�����a�Пa_�k�&Z|ctRsiӔK-�c2�������T�������˹<��h@d��r�@����E�j���E�� ���[���p���G�n6͋��=�9����VN�"�v)J����Z�'�u�������B$��J�D�`ks���C�9��C��.E�k�<�w+_T�]ֱ�����H��q8J��_�6'���`��]�I���]d��Ү�1�� ;�Ⱦ�2=�+�����d^����\�;.���}������Ҵ�8�0���&�7��&�W
�������)7(�m���w����MGy5��z�s}r����o��;�!�vj;���@$�i�"��}��)8|���Ľ��Y|��8�Y�ͷ��\�WT�������m�<of��^������c�H	~RR�a�fy�FV����H���^pW����o�Pi�5m��#����h(9����0��	[� y�=P�L)@��h�]w���`��������UB=-�!�R, Vb1߽Q��g�(lf�>a{���D�6{���Z�@��0&��;¤�O�|�Z�K	~���*n8��нÄ�j�������r�O��Y?h�f�|�>	��/�eV�z�^BX��������癭|��M�������r-��2��!��\Vcm������J�:7h���`����t{J[��-�x>��'�d{1�;��ڃ)�JK��w�����z��QO_�WR�|�9�{��e��s@{W�x���q��E��|E��{W)n/;��{8�kȁ���T�`�N�r���f�]�#{��寿<�o>F�Y��^'�A������$�#_�5�H���N�������W��X�t
�R#�`�V��
^EA�i�"����}P��K(|r�7l�K�[Z��*�)L�DA�z2��[n���	4` M�3�s�򰟎R�K����H�T���ؗ~���y]{����4�!O��ˎO@*Y�K#����
�	�������z��4��L�G�b�0�Ӈ���8prj��~���E���xws$]�ǻ��F�`Rx8�D�d�g�l\���A��G�yx������K�N����m���t�C���mcBE)�8����k�����ur��y���pOE���t_褶�wNcH���.�&��Æb����(Wy]żI�q.̑}����,�N���b�J���� +/���_�HY�B|u%��S���G%������AgF��F�CN�SA��둬Y��WDo��h7"��_a�u�4��%@�+��Ļ��J�|iMJ*-��U<ƣ�`9�x�J�?#du�T���ө��S�kvn}�ݺ%�ʀ�=��|.����E��6}��{`]�ہI3VE3�Ye!�y9/��s�t>D��;���9Ѵp�2k�떘�ξ�Og��F$��j�_����ٞ�Y���~K�L�]�V�[� '���dy o��4O*E�K�C\��@��Ӏ���!�/"�m�ı[
���	nǃ�;�;ރ�چC\0��8L��6�VOM����UnS��,�0���=Fs<����g��g o��uz^'+Q3Y��j��F�xVG!Zq�)�Mh�JN����:ŉ�=�ScZ���8���i^�y#��|H��q�˵7�� Z�0��!ɗ�eQ �1�H�$}d
���ݡ�7��`awRǬ�1"�|�[��������*���~�9o-����t 2[�LX�z����IaM���O�|��������GFn����/������ʟYg���d4)�$�tޡ~v��X:٨��������y/z�'�8ʄ���m���q�� V�}�Ä�@D>�JjG�ϲ3u�KT�.y"/�q��P��w��Yf���W���iPf��<���>���uX����� $�.)��y	w���(q���!7tB��1W��fa������wp�Kq�C%��~�^�<G7�O���T�F�xE�F�}�z�ph��X�y���I[N.�`g���
�����j���Ca��t���1���9���#E�X�j7n�~�Fޙ�߽�¸�xf�������}����dz ��`�0`;A�(��I�t�`�;{#�)�3}��}�T�
}��n���2�\=)��y����탔���tD��F����8�p��/�1�|���\	�:9=y�;���q���ۃ9Q�|��z�����?�\�ՙo=}*�E��vLN��`�<��p�>�P��(�-�3��ǀ��Sh�����QYc�.oGTL�#ioQ1��Tu rT�Y�"}��U&y��7���=koЯ��F�CGs�3��~�){�0"��t)�]���K���ʸE��xe�?��`�T�1�zBv��ر�=�j�ù|\5̏ו�H����BrS����T�,����#6�$E�%din<�Q��ɧ�ς���^p��hO����D1%b�g �����w)z]sW��9����&_sᝯ���]�N�E�{H`%����-���|��g�!���ؕ�5*�ď�� Ѩ�ȼ�4d$>����r�>1/�8|�8���Һ��v�^��5~l���70��C��5� �r���teď�<C�˲�F!��q�Cʋ���$9���O˟bvә�gh	9�Q�i-���[��x���U3lK��_��i�P,#q�	~쿦�.��3+�
�����Әӽ�:����)z`��>p��5;xx;�s��������Ł=:Bb�bEM���!r�GC^V^��ZkGʧ��k@��?�o�g�y5,/tf��y;}�����$�F�	�l�C��1ۃ�v��C��{vb����o���w���\zh��놹���8�yn��9�塰I�,oyQpx�D%q"��7ښ�����=���/�zms�S�tj��O.�� K�A��s*��|��v�4�Olt�gJ�D�4LpΌ�H{J��kH^J_��L�i�|}��"�W�p��	���-������)~\S!�$�֭��ON�K����U��E>��&���!������>yo� 9�5��o���`C��`��=g1ۿ�<�C���S�mz������-����MNY��9\p��mQ��7���p3�JY�;���/��.�l �,0R�g���O��_D7	.tm�J�\��$l�F<V��0�k,t�/��{�zxS�Nn'w�e�A�0i:���>��z����X�nV&O�xF�#���s5ma J)vs��\�(�7���;�/��9b�nV;��
����v4���|��(� 9\a~�<��}��g�>�JD��
�)�����˸��Y�W�o��/i�Jq������<S�ٚM07���ĚVу�Iw�7m���F���pp��Ы$H?|�I�}�Ѯצ���0ԗ�*������u¹����)#��� � |���~�b��8��b��?b������͏��g�/���=O �uyh�
9{u�+B�ױD��g3�%�z4�����l��v7h�'i�y�.�%�@|�iC��t�	(�#��H�w��#��l�X��N j�x�����'�Uv�*|����������;˜7�E�Y:�ＲE�>1����b�W���6�L(�;s�O�)=?l8|��	F�*��Yh�C#�ؙ��i�l����}Pf���K��w2}f�������_J|�̀i�2���,�����k����\������.�R��6�by@`�躮�r�0Y�_��`��i{@0uG���0	Z)yo��X<�tr��9v��Vy&����g�L�`����&i6��dԧ�p��s/kWn��x$X����)_�gi~_p�(�"	����!a�u�r����-�(���l7@=NT>�M�s��V���!I��x?n�{��j���5Go�����g�?y���O�����)hKK{3['�eeѪ�V4��Z�Bg�<�|�23��sC|���P���0��q2|F�+|:_)�7��|���7(ط��+V�� ��Q}9�B�K�!ϭ�DV�ʐ,^�
X�kF�����9�"��%r/�I���N�K��:��y�֌���#j�07��A+~��U�͇��g�PV�S��\�ZMd3K(�p�@�k|��RP�Y�5�v�����^?�n|zT�s+�������-�M��r��J�"�];���o
��X�۲��0��wqa��8�������ڵf�}��i^�/�ϓzCڅ��XP�k'�ļA_;�Q�ڊ@��=Hx�F�°Z;f5�x���	<tVJ*�����L������.���ƅ^m���FA�C���ic�7�K�p�*���*˙URlпKIΧ�Ѻ<���"y��O���gB���$PI�c!Ԗ<��Lh�#�$�)B)�y�t�(�L��q�,/���c����3�~گ����%ݧ��1��%�iF;��SkÔ�;����G��>i&��k+G����n�\Q�n0����o�ٵ�{O��A,��t�㚰[G��V�	@�t�+����{}�(�_�3wI
�h������׃���.��`[�1��2=���)⧀&I!��~�W�׃j�@�����/�zߧ��	n
����&���O��ƟO<��=�P�g����XQ�aK��Do��{����"��	�I�����
���)�7R1��,�K�7C�i`��D����س��g��p	���z �s���dc���@���{Ѩ5X9�������1m��ȩ�#��_��@�	 �]�x�b�('�Zۏ�uW�.���p�P�Wj3߉�'D��]p���e����ҹ	��<"w��涣�_ˍl���Ph��gT]����'�c�|2 ��`]�V��$���:��ooF��A�4��,�h���Kh��ђ���J%�;C[�Ĵ./�:��W7o��$��0�Y��\�"������{܃�6��~���������O�����8Ԧ:��f8~�����8Ve��~�&������kALOkM�MV�]^�DWN�5Pq�\q9w�Aۜ| 	�'�~�4S���{�<�i%y��,o��C��髶��B�C?'mwr}@K��7Zk|��� ����ڦ�P�h�C��=G��J[?���3�u�?g�.�M
xrk�G9�m#�)�l�*��0��V�bt`���l㳔��8vP$i��OA�i�D�����ۇ�JL���`U�����Gwi_d���"��~bc�׳O#���3�~ܦ:c�C?�R�߱{����q6F�#͉���y�(Ay�E6py҆��*�|Ѝ<EJ빍`h�]���c�w���c}rL�(��Ŝ{�
CW�Z��Hd���L��60�n�d�R򻅘��J�] W`�_��E��A�W@���K�����շQ}��8�)���۸$�[p�Wcjq�*{���7�$�.�wa/��>IvH�L([8�q�����~y�Q{�rZ�V.���?z�l[�vH��!)�ɜ���N�N�M������l� ۋ�$�юyb�C=�ԓW�e���a�<�;HJ��gb���k̳֟�����2�2��[pW)� o7?�.8���~��R����V�����L0?�������P��š��!�� ,:d�;hn����|vƳ���j��|{��gA���.mh%�M��|�������y��^�'1�'D �<�N9.l��D���v&�w��f�Z�CƿN�hMPbа�W7��#8+��Vm�^C�&t�+n��3��_X���,rI�|e���A�2�;����6�&8Jz�u��P�I���Q�9K�ǣɭ�����v����*�u��|�ʼRW��R�-t_p�� ��nAo�_�ç��sv�K���H�Ǩs�ݤ[����	Q*�ߪӝ�Y�7�ϥ:'�񉮧�&�������2;�!7j��"g*�D(�hWi	2ύ��Ykd�y��a=�шgx�3��Z��C��V���'+D�N'��#�u*�c�O$7:��d�I�O0~%N?q�����Se��>�zR�4��#�G;�D��J���=�r2y���d�<]�m�d��`s��En��ŹM�Ydu���6����J���!]p>�������'�r\p��	{1���)�Uv� ������ud#�c[�.y�U_�`�튙�Ѱ�G�X�tA?~��U���`6#���S.�i}����V�,�g��9�!��'䅼. ;�/�h�_��{>�ڀ���6�{,��p�_x�׵�D���|��mk�?B�,��@\&�#q�!d�ɘ�s{Ml�����11�'�����u��8�x5�Hy��`�bdu��������[���E[���ƱD�q�:���)q�����5�>Y c�.*�
[�R˭[	�m��v�򈟣�A��*�R����� �e��� /�o�W�<���%�g���\�a���HH��b<e%�vP�9�j�#���uG'�'�$��������Y��:v�A&�PVgy��c�W��G:�w	8�`��:^��<�^kg{eJk��> �f��1z�����=Nk�eJ��x�Q&wgx~�~ �p�|�c79mz e�B��r���-�"�{c1y���	H�̢zj�;�Dz���}:5;ME���ΆC$���[��#��vk��,�/��|;��3\����������p������R����/_#C;ӜYY���.�;)��-��!���7{�򎖂�'6�bM�ʍ��a�~�*Px%�L3��4��m�[�+Md>�%q�]�9tM��k#De�&��,���>�jr)[��}���#�C��V9�����k�����A�����jC�s�����v�YxS�L�[�#�$p��CA��Q@�E�6��n��'�3(��H���.�7 5���҆@vX�ɿ&'�a�������`O�_1��K��|/�����<�|ip���#[�̀{5����:9�G㩳��+3p2���u�������	R�����q9`zwy���'y�~K�yY�ҼP�������������e|���W(b?�Mo	IN���r0�++~�~b0i��I�7�����X��U>�p
�����ܷ�)8}Gc
'ُL�w12��+S����r$0�_��_7�@G܂o+�1hٍ�K�}�$1|�"�PC��� '��ӂ�rm��#��q�� ���J��I��Ҟ�ӵ��<mb:.oV/Ї�J��l��2��*pP��G���֍:t�FJ�P	�v��>C���{�Z�ி�1���2�[ųlp�\�����/&<\�T���AE�b7�Ƭ�~����z��#�Q�
�����L�F��mp�����N���WH49��.޶$3#��C��o{f4�ᛑ�~�~x��>ꣾ?���2��ڵ��?��1i��x�zk�d�F�@�3a�J���?ڶh/;���b�=�w�f6���œ������Y��zh��0;;���w2��c�����
�&�5���޵����!*:�r��`�O)�eЭ����-γ0�p� �|6h�I�Hg\��wو�~�r5N���B���<؂��d��%����o�m�7�B;�~4����.�ཐ��,�#���R���3߳�4�v��ڔ���������t�qS�61w�?eϯ��q�Fmcٝq�,h0f����O!/�½���*}%�ǃv.���-��w{+YZB�p�%�]m���Ŕ����=�3��ړg��c=��S�R~e�:J-�i8"��'B_�Sl�W��w٣Q�d��x��:������0�7� �pl�i�V6��`c9�p��8�����0
��7i�����w�� �,)�?YX�-i�(GD�Dx��|H#���S,��j���8��������v'��2��qb�.O�g�H�:�]�\����	�uLJ߯n����Z�5��a���Q���N���Z_�M9EY����.�B�5����ʏ6ivm-nĽK��r�n�!;�v.#����m�Zk�Y2k�� s\fuv'	>-�
G�_p�����Jr��F�YRxI�z�� =l��A��O���u�� 5�3`�7�1�:���ƛ�L���4�s$T�%�C�"I��f�q�Z���X�G���6�#,F�q8��?��۽��o�ü�X�Q�F;�%�������;�|��n�	^�o�Q���S+8�5�-G���>S�z�6��B	r����O��X�.0��cY�B��~n�Ín?���� >y�0�~5�2�C���|���.����Dy�����l�}iu4x�od���O�3���i{�T��f4�UJRm��~F�Ӹ%Ĵi��}��ń>�G�:����E���e����>�K�SO�n;������l,I����9���zgRw ]|2߉����H6~�P��=��݇b{���������8�
�=�'&��yٵc���E�	��'E�#O���3������v���n�3��ˮa֮�J��&��K;<��Ң��֣$�Kw"�+��R�NT�1��+����F�8""Lٟ���=�C�^�7����4t�_�N>	ʳ�ei���bh{l�{�cGX3B��JwX
����2�^q0S�&?�M^�Uv#�O:H��o�f�m��iSۢ��̡����=
(Н!}�\pf���0�_���ξ�n�����o7$=��?���;�^ݢ��{����f[�Bc�ty�(C4E��B��\!���$-�i?2o	�))���B�Glܢv-b�~s-`��@s���Om�C��He��%yhG��s���xa<��`��+$�P���Fɤ�֯���å4�F\�˪meTv��e���� H��#CI�d2?'��!�^�Bpˆ4}��}98g���A��г��A�2/��'4�\�߃����ٛ����6���H�2�V���ATo����v0�S��A�~�d�09o���,��N��<�.M�#|��Ys���mE,�sm'�B6�+I=�ub���]����'�K�f<����6�J�	��%�&���d?�Ù�?zR�H�4w�mO�6D6��F@��@���/��$ۃa�]R�[�F�ʈ��3��'p��F_���"��}��zg��N���Ҕ����pQV�>Uȓ�7 O��ҚY8���Q�cڀ�-�
4Ww�0)����0Mp�(�',F��-Y�'÷v�2�+4�hOx�mrt���d��X>#̦Sƿ�N���';}��?j��)4����pm����(��`���*`Y��{�91}�
�����C�[���w3�{��n��3��Qy�6�������e������z9>��Q�����.����<w�'��t��Udv��s�5˙me�����9�������-�q�yj ҂"f�}����Z��ÿ}jt�����UX00�.f���1�-��o�1�$Dm��k��l�XlMM��h�gM�����C��U>�:LC��:�{����2�G.��R(�)��f%~l�����ЏL�,����ԛrK;�Q
m���t"n5
�fr�h�v�im_�t�gCI�}e80!�����-�2-��j;2�m�q��Y�~&�N�r���a����g�cy~ߤ7^��V��e�9�n�h6n8�����!�B�%�g{�5�m��.&��l��4�ݍ����'�'�����[:���i�Ǩ^��\;����~�o�G	�f�ç����k��QC�w7:_>��h�m�E��U�G�
&琞Z�\?�Ն]����=���sD�@ߠ?��� zV�}�g/����.�>I-���s���0����`��O=�0�S����w?HVU�<
�P�ݓY���9af�93^�1�U��X�p��֕��ة����n`��;]�\�W�$�Dd�b\�ћ(ṆASߎ*rEw���h1�)����y�CC��ޘ�4i<)�w�e�B����1pX�S�X�vA���� ��Sph���grD��r���up<"�P����2��Z����3o��fmQ��w*d�Yz��-��6X��0!��b��esD�i���8=>��)uˆ�&`�L�l=�%�������t1�.�������9z�8ZY�`��vY AP����!đm�H='-K`���D7���sN���C�f��'��:b��m�j�n�x��}AѺ�c��#�E�O�	l��X�S� ���s1�F�S�U�VAH��L���`Ƨ.a���0I��%�V�G���R6"����p������zj�4ry=��]�L|$Y���L��X!�jd/���,���9���N��#�)��E�g$���,�Tͦ�����j�^z|`��QqEu6���<�a$���llu�>=Y�\�
w7_�_2_"^��X��.��(�V嗀�AJ�=+��uz���6�2�\�YqQ���Tx����{��5D���[2_#}���->7�� �N��vG���l��Y���;�!�D�qh�����v7q`�xX�O��t���FU�N�G0a�7݋	�"}+�-��=��gѼ^�9����U�Ce����+N��{
ڌ���k�%�9�j)l=nT�P�����/ ���3��g�gb9���;y�L��&r,�-B����"�.��h��8��������N���}@���~���It�N&0�T�m��PT���#'܏u(0m5�
�y�Y�HK����-�A=����h�"}h9��<8�o�/�\��5�� 
3�kg��@�� i�5�-&�ڨ��F���bwp#�ƏڑIo���	�mc��'�f.��^�����S�d�I�����2Ђ��$+����璕1�d��KP\E�Y��J��A��N��n��.������8ULo�$�E)���� �%����@y�DY��������vl_�S䪏���Й��Ef	2�)�֊��y�h�çڸ]+���!ь<��%��a��#/�'�"�3�c	b�F�р������!N��������p���_aHr��U��IE���nK׶�iߚ���V�>ۃ��=@��o�K�/83_3��K���XB�|/��ˀ	��ҧh����.��	Q��ЮL�j2�g�I��X�g������L7�#!�|�؋]=�˷t��M��:�n�p��?�Y��s��y�����,�О�s4�<��8�}D���xK��z�L\��u,fF����Wۓ�ƚ�����9^|�B�ف_珈�֦�Q�ud����>����{�=��x�Í]�u�>�ƍ���9dp� �:�rj���
`�6�x��k����p��1�7����B��@��v3?!����5!HB,�
�m�"Ň�8�+�, ����y��1/t��0��e�O�5���Ef��:���z8(�o������Y^Ks�w�?D��1j���N���:|;��V��3�Q�8i�C���0?\74���y��5��y���@��{^����~��UX�����'�t�|"</C�F��P�=W�<cIo:��'�F5���xW�����@ߨ�(�o��<���%=8�ĕ��[�vwĿ�"�I�%#���Z$��5���y�BG	?���l��Q濽Ĵ�6;�Fu��ҿ���߰�Ç��n���1�'S<2���BL׃H�����q���
+�/<D� ��,���p�M@}*7L�xj���,~y���� 2��}X�nY(`O�\p��X�ģ��n�~/�A��X/�v>�%Dw�����P�1liݍ�ŗ�L�t��b�c�}~�{7�ѡ���HRfG�5��ćP�ɞ�l/fo�&�o)�~P���7���\�0�w�BUD���<�׏��%�,7k��7�n�O�麠��}����<�?��V��5횬��|��J�{�������>I�	^�X�mb�z�}0�*z��ߠ��X��)��rA��x�`D	`c₼1�c;1�g=V�JB��2�Wg�d����󠝈k)O`�^F{֯H��������W�ST�Q	�q'���0���usY�%;�
*�Ƚ���FM�y3�����4�!5>��t�5C�
�v(���C��.����9����n^�v�G4ZlPF��]���	l���
�wB�^�j4m�l�
���R���,p��V���j״V�Ő�/i+�fX��ʅߍ�ڏX,N�Ȣ�1s1��E�#W!��fr�}����oIP�"qaX�$<��Q�?^�3�c��y��b�Q�-�վ��2��;[�WH|����c-��p���8�?E������B�L���:�3�����<y8@��i+����z��/H��6�@K��9�;��rɼ.M~_p��V���y��|�X���e!�)X��#�= {F�b��a��"���Oy��E���il3۳��fg�T��z`���t�h�G	N��xү�6�Q��@�0/kG���6�~Pqc�����!�պ'gk'|9�O� /��� ��U��@_���޲|��{�N����4z��z��k�3�l��Ȼ�n���B�Ǘz0Cާ�������o�?�$~�A�����0�S�~�!��Y�t�0����4�����-k%������4�`;�z�)��2ڳ<�N�W)}ި�������j�?���'���J0��x����º�˓]�rZ_������j�;�։�j�W���޵������_����gX6�댆�[�/���g�;��*=���]E(�A���N��I�o��JD�\��}{��r�
��r��������x薝w��w��q��}k����;,��=t��}G������7�E���O����� ��S���]n��#~�'��3�aD����4w�*i��^m���Bgиn��:�d<	0 ��i����ڃ�f��0�+e�S.s\Yۮ�@�
J�z��)u�.�i�o�@��!\����i@�����C�c�
]V����)��ƌ8�3��:\�Q�����G������*�k���o����4�S6��n�H���^�3�4�sa]㪣2���-J�^q���ex��.��(��ͺ�>����z�n� �8З~_��W��JA��zA�7�A��Vm��7b����E�6���1��LQ�
]��c��G��w�,���繸?C��^��,/kg�v��2hoԯ�0Y�o��/�+=�x�z�΀�w�+gH��{��N��%<���#B���(m6e⏠{&D5�/V�%3�${x�g�A��)���XٞK�����
�A�iώ�0?f��i�?=�Pp,����G&E|�}u���bn�d̼l��	��*�<&�*�!��y�?��z�����P��
c'/�Py���E-�v�㘗����e'<²h��W�^�8��ya���A\_�g+�OI�a���i{@����d�+}�i��������lػ�c�ka"��x���uSUg�o��nȺ��.x��J�h%�����/KR�'��S�i)���:eMemO�f�K�X<��SO������@���3vo� ?~�O	�Z�e<�b���,S&�[b����&��؈��(E�b�W1k3���!s��.^�|f��>S�tTr���J`^16_�?4fO���X�͛�Q�2w��!߃�e�ȥ]W���oυ�ȇ����v��l��Vp���;��#��S�� ��'$l���n����0\p�o��mT�h/d��eQ�G�L�(�����xˠ,��l��A��%�՞9��{t@4KwuKhh��gӗ���
���}j�qA?�v�^^�yq�h�$o��� |\��|=���A��^LF_Fgt�B�p��u}�OoȲ����m"2��+&��<�o{��;zW��zF��x��z{872�;{�,� ��X��7p؜'�d~��n�5�Y� ���Z������O:�B�+4t��{F��C���< �J��^�F��z	o3py��́���X��o�u\͢C��8)��h�#�?�� ����h4��$W�Tn�PN��A{��z���+���\�On�ק�ީ���B�u�ӾW��C���LJ?��N���ÔWh�:{ݞa����Aa��$�#I'Fb�߀O��	)�����k��aI����溶��Sm�#k_��̝��P���vS����_��������~dF��y��0�M쉑vZa ���V�1�>��G��_���=t���:�ƻ��>z�t��8����M?�-G�Ĝ��`E9?��W��Q,���g�w���H�'p$��������"莆���9/$���� �gh�|����^̈�zw���};H��W�;�0� �2S7>��4���+=]BL��$�)����Y)��>�W�W���x~�@�<�
��_���-'AVR����ɒxM��գ��O�ŘU�(��ef4�\i���r+b�A�"�<<��N(B;3T�@^�qhD@];4ɛ��h�⓼2����e48�|4h^��e&iY8��B��I���ME��C�C�O����V����R28�t��|�U�
��ꎌ��
���Ikgq^�ȸ��X���?
�0�\p���]������^߶�e�-�$hx�A?���HΞ�ػ���l9[/�'�u�^�=�*3?f��9c����f�^젮s�����2t[󖾍���� ���h�dtG�C�>yP`t�X4F�=�3b��^#�1p�eN1 EH�Գ��g�׆F}&M�U�ė�Wë~R�C���<	�F��m�?1���aUW�6���\�e�N.�yv��OS�\p������߄�QA����<�6�씗5�OB���S�0�rw���B�Іr't)�MI�tO �݋ѽ�0�$������Y0�#6�s�<}�/�푆lodH��Bڱ}�C�4�	��ғ�*�����E��R���D�6ڎ�E\і:����wG���W�x��`� N��q��O�K���^= #��4XPڗ����#p�x�}�Ly�˔q|j�][,̣�W�<��W�
L��qPd��*�ڠ�C"�ռ��4�W	�����%���{ʓt�)-���څS��Dŕ�̾�&x�y:��(��Q����م�+�Fr�h�����$5������u���U���땒ŏ���0�kёC������@q~�\�4�L�>�2n�߲�N���w>�)_�=+�Ѡ9P���Q����j����M���o�.&��!�c�jCf��}�j�K�օ� Ģ��>��]��?ϩ�͏��h��ft��Q��}@�~h%�>��Q������6��f��	��|�Ւ�86L�S�wP̼"�r��P��O�zq�#�8����ǖ��j�<�9�5����.��+z�5�����r�*�y^-�b]�<� _�����$���y9��ꥸ�`�E7ƅ�g{��SyΉ ���l�%͋
eƼ�}��1�=ɓ��+1�y�S�9����	�\^�GI�"�K�mRok�ݬ�l��;[K�~q~v��8���$]��n|E@��\��=�«��R[ml��ae�}���D��yG��������;���_�v�e�[�Q�c
؏O�rx$2ޏ��[I{vQ�����"�`�4��$�}4�SŔ�(�Ǎ�N9A��@_�s��6�3�83��$2�J�c���4�<�>�����U2ZY�t�ŖmH<�+���\;���2ؘ��&���x'��H�E���_�=p���Qf���=�6d}���zG�ǡ�*W$uj����rlO%3�I�c�S^'��\p�i�� avZo_�O�ܥ�y�4[ta��5zj�n��7j����|���r�������������c2�;j%;�������DV|�w�����M���T�31�k^y�J8f�[��ܾav��{�H���ص��?�i��AoSX�L�|�U�5�i�eu(I'H�A�0x^�Q�}/m�I-K������	��\��Hmd�1�8m(�d��x#�SܬT't�T�/��;�+���>�//7܈��n�[E���=w�h��g4�ҡJ���n��i��'�s�/r��fَG��M���R��}��f�ޗS��H�i�F�������8���%x��u�7N�����9Y�jtg�#���~K�g1���}�%y���l�"�t�Gy�~)?0m��B���p�L�����>��Lh�x5��|:���r�t�Fx�2A<%�\Y������!O��q[�7H ���dEF�rԷ��O_�^��eӃ/�����<�R´R�C"��c8p�"d8��Ï��@��㉦O��z'��Q�"+��vV��"�Q�pl���`3Z@	�!�
���y�4�mq��{4p�w�v4f�ʘ����sBѼ^GC��r8�_����^���r t`��
4���h�,���3	���8��g.cήӸi�F��%�l���~~��͌�y.E�q2��qλ�$���.�A��{�Z�!)�F*��45a]o��r�ɧ�?|kܥ�4}�#�mr>��/T�K�Lr<K�����k'��mu>lC��aG���� =b�|;(	��X^�?�/ņo��/F��������>�vt�W����u���9{���>3�I�qzz����z�އ5,>ۏm~n�*������������Y,ł�d��|ZX��Q��f4Sݶ�uO���O�~#������;������x�M rVݭ77�=�\p�������z?.�r��O��j���}7p�[«���դ[�jtHvH��fM�_0����b2\ۇثI;���g1���yiBߤ=7�#�%��x\�f�%�P_,����5J�g�۬^��9���KIDE|�p�6���C[�F@�G���U\ۭި��{���3}νB�!��N�\^��A<U���L;��q#oS�[��t���r�d
����щ<4 J�D$4D\<���`�1�QV&y��S���%y��b�툾\�;�C��hhpP�kH��AA��	� ��Y�4Z�����jٻ����y�D������\����\�`V5�fX�g������{r\/���>z��\�H����2�	� E�98���ƔpV�%l��n{$=hy������~��I}D��K��������jsaO)t}�<8F�9�{��=��Qn��"�ȕ��&�#+p�C�s�4�M�4��݉P���Ҽ���j����<�n�6�}f�G>/�C�~Ɣ��� O?���os�'h�"�\�&��s�/�|_* _�� ����\p�Yp����%KJ!��+N�S㨕L�$g�o�O���m��~�_P��+{1ݞ�y.ǋA;�@;��s{*e@{٧}��wkχ�E{3Ґ9@��Q�s_����Y�y�n`�!�.��$�=�;*�k�^������φs8�8~��xK&�'���,��^��q��,��~[�����~f��|vr����9ꩲF\1��v�4 }�	Dw
6�2�Ї��
�!%�3�_T�3��a^=��h���S���6��$W�Y��s;`Bֆx�k� V�	�6km36���M!3��eܳ���d�3:��?G�,Qy_9��R:��@e�k�$�h�{�\0��&�n~���'��'�$` v��xVGV��Y0q���<���2-�����e�}T^��N8����ݗ)jO���B
Kڰ_V�q�4{�}yܛW��>��.�_��+�Ԯ�/o5q�������O�b��;�������̧(��) s����l̑K%|G��F�q_zs�NrDJ����q�:�A���!5��NGm�p?��ʜ�m+2�ه\����;���"SE��x�=�V�|���Mz�.�o�+��δ�;�y#�>���x���].��C���%hII�[���.U�cZ�/QJq6b�{��Ҟ�yIۇ�[��HM�f����x��Ѿ�� ���_�e����홙�=.��d��b?�ğ(��B�����;p���=N��.��@\������ލ��y�������\��iI̽⊬w��( %m�F�Kv���SԤ Q�w�QQ`S�+9�i��)�.�hV��z����P~/���Se���00�R@��4���fV6�P�㻷��_gҚn�Qgk]0Pt��a�H�j����m,\��h*Y�������޳�ɱܻ�������O��l¬4Ґ칠�F��'kr�y�"�$P��T���E���k���u��M�w��>/���~�^?a�x�ou+��wQ������?ޞҨ{�l��Eg����� F���v�_����y���o�l)�u��'�������zf���2���P�^Ŕ&=XDX^�՗��fwz�o��Nш�?X��O�#�,���<�5��������pd��E_wMJ���j����@T�8=n�iv|	U�g~�qL��,��m.8z$��
�+YV�d�nL[-w����۷G��^B@�	 
�@tJD��M�q��c���0��:���@\�kk�պ3�\p�G`t��t�3n��^����σ���w��O�G�ۢE����	����� b���2 � ͳ����y11/��q?��e���A/�ѓy[~0�f�+�	�������H�#�,;;Hb�f��}�����bs4R���V�=�0��簃w�G�tEV2Ng��+`��u��u\�~��sgQ�=���� �v�ׇh�� ����j�W?��O�]�Mo������<9Ks{�dij��vdW��ǉiX�b��ż}�Чp�v�l��,��3�&Hz��z�T��PFh�oC��_��}l�d�MT��l-0S0>k��Q���,$�����fJ[�Ø@w'o�ص�ke?�0�s��-xC7��7����\p���L׸C��D�� ��A�r\�8B�p ��4�F��>>|�w�*��@�`�(}��2���(�c�����i�Z���J�9w������h�'�y��8�g���3?`��Ϭ�F��Z�rG�O!R'�#7$��i�{�1�1�YqW�!�ϣ�[p�=����'�b���{~�+b�u�G�,Ûzw^&iG6��|�ܱ݇�l#|���>���.�����w��]p�;l��y���>��˜�����|F���F`nI��ų�n��uQ����u����?)f���	��<�q����ѷK{��4�~ˌ�دnD~�1�ߢ6=��J�hH��@̋'�a��+q���[���Ztg����Gbb1�{����9E����xp��ߠs����7��[n�o��:��8TZ�&��� ��4���w�G-�̐A�N��P;�{P�C@!��s��p�k�Y^b�,�	�1[ab0��&S��� `D�X�"oG����ڈ3(����ÿ��4h�I��6&+K�U0
����7�4�O��F�o8h�GӃwQ��ozb{���Q��c~�-f����$�|�\�_��ֈTϓ�/���!�Zy�Q���{�^ĸ[CK��vf������՚��T���'c���R��~>~Gש$߳��L�v�C����	C�uY܉����4�"�I�n��x-AO	�� �{⬸�:_$^C9３�[W��`s�7ܗ;�.���.�\�ѭ�-lo�<�?��#����@��d���L�am�쇊�~FB�����A�wO`�^�W��7lg֯@Ñ���>���H�}�?�}�mh����;{0dIV�b0�8O�u����?��(4�m�R���ǈ�s�g7p\���N<\N�B�W8U��~����,��b��h�dH�Ț��e�e!M���Jpb�.`G!p��u��"���0ùC{�ڑ��X>֝�=���*��3ފѱ�w��EA�$�l�_��Y�v:=�Ȉ���Zˆ�ȫTFpo��ՏO&�~�n�S��3�'�:7r���Fz�D�|8��kS"��.���_�d����Ւ�r�?g\��uf�۱f�1���[#7`5�l���/M`d*�ļf�'�Kt&%�&6Q�o���lk)�S��
j׋�<T���P��=
�ܗC��[�Tln���x%5��l5E���#?#���qN��܀Y�5������yiq�6����6/Z�խ;0,��I�tE)�]2��~�S����4z� �'��.��������>@�&�
�[�~b�q�7B�i`d�v{0\:�Ƿ3�{��ﻸ� ����E�Kv����C�-��2��޾If�}KGW���C|O ҧ��aV������,�f�A3������:�e�Gƌ�o�Hu��x�U�	���d���������n�U>�������D�_����9>�uA�BtF�G-�`@�4�!��.�xY�C\��Fy����)���!���i�f�&�K�W�2%�p�@{ ���sɼ.�SI���W#Z������|r��0�b֒���v��Io��izTT4^~�������?��w�o�)����g��R<�.�����F����0!��oK�������}� �m���c��VP*�+�фډ�0����7}����V�s�{�@�$� 	q%�I��DѶ�JI�R�*ǥ��R�$U��/�7R����C�8qʮȕ8�K�$Y�hH� 	� GpAx��9{w���Z�z�}�{Ϲo/��s��i���k��a��lf}j[��2�g�(e�A�&qePva�BIJ)�,�b����u�I���/{�E�2��g��K�@�C���5�kT& ���$_�A8�ԇ�}�q��,�ҧ| N�!	F�ש�p�IRr2���lC�u�g�R��&�uu"#�����N� ;�����1�L3ʹ{:P�Z�$\�ú�z��g��0o��t}��}�X@\��v2�&����ѽ����ߣ>��h�P��x�b9B����*��W�0�l�0��������Ԃ��v���d�d�[����C,}J��d�#N�(��|Ec��Q��<k�Y���L��������Q��ƺ0U�q(����C���X��:�����@�&��,s=vAӞk��$�P��=�yrQI[ȣKk�j>����0��Q�r4M#^���O?�'���W���n�j��Q9,�a�s5X*F�D��'�>�+0�[�y�",�ˍ�M/�nWan3���%I���ߴza9��P�#ѡe0�c��0,�FS�f ��7�F�d>�Q���o�zR��\���Cp�J<h^�w�m�3��N��'p�dR��̏N�!_�&�� �:��2���������L3�t�(Lq|��y�sD-�f>����i� ĉHa=�m�X�kpp��jNa0jX۳�HVn�����u�GT���_��I"nB�m�7��R͑�[�8I��ʚ�8��2��p4��l��pr����I��Tó'����r�|��OZ���a����s���a���XS�A($�TA���g���X���i�I��4��SV����c$4�57EFf���B"Je0����<bQ�94�e�>f(�����<�g��U���'��c�r���n��F�XN/4,Vs��v�-�立���NwzN�کsT-�n�,���\�G�9]�9�L3]*�	���y>���!R�#�xo�:������r�Ik,;z9=�.��-��p��A�������
�C�����"�D�>��ԺC����׶��0��-IUn�e�J(�=�#�Ac|��07�ð��H����ô�¦���(�%Y�(�b �s�;��d���I'���Q>0�\�Ԗ��)���)�lz�u!W�S�0��01y�sQ�YE_��{�[,��Ƶ��|Z��K����"���.�����<\@4���z�4Ő���kjy��;ΆD�	��
�� �}��PX?;�=!�=�5�M��@M[�f���HX<�]\?s�����C�}ZgC9���G�Q� ��@ �e6��<sҋ|�`@r��r^ZL���<)=���fz>���|5)�0y�_~��\f�i��fڄ6YEJL&r�.a�M��kv;w
`@�s"n�� @wIS�!�g�O�`4���(Ny ���B��_�1�6`#'�&|X9R���C��
_���4�<�O��8���J��	���H��:/���NE�a�aj�S��5�T�E�#�Zt�$��!*�Y�Cgv`ȋ���b|δ)�Pߗ���q$K �%L�Ți��n6��J�ǀ��T�!�>�D�玕�����<��$xÇ���5�16��!|��ތo�[�0g���p�*o>M޷�Y�KX}�8�I����6td9@8T�
�z��+�qL�=r�z���Lq"���J��1��+_�]��~������P�#$"����́�K!�� <�,pj�9z��zԜ7j�����G�~(I�_,,)��D|&J�r�����0�Gm�V�^�̚��4�'���V|<qu񳬳۪^� �@hx�բ��t��>�� ������]0fEd�F�+��������}��]��8�:/bcF�n��R8���f�i��f:?�u���c�?C3iӎ���w
]�Cc�MOĝ�C;`��Ic�QU \�|<F:~}��pn;�*|�`�ZF�[+��%~W<YM�n|�CFь���g���p���(V��~S{J˗Z>*�W� �VbB�@�V�[��]-�&녲�˄1(J�r��4hr�ql��E1J��=����Bx�?�>O�Iʎ�%�>g�i��nV�N��q��eg��:�I�b�&'�=�?�di��S�}�%��Ψ落e(�A[��K�w�������O��z��m$KR:)+CK,tR'P�8ehy�r֩�#��DIfu��#>VY(t�����6s�p���c�S�E�����|��yt��+C��$RU,�GS���혣��?�3({8����S,�?�J��w^�J��@XNG�t�yca��~���a:�J;pX�'�/F�P� A�\-�b���P�G�a�O��y��J�7\�;�K��*AA�����7D?���=s�?������y�Yc�_����y�nwY��j��������zyf�i��f�-����۵��؄;׬��IxjkK	�×EvF��X�9�|��EJ�8����S5��$g2��h*i�ǎ�k�E!�(��p�)�8:����|�â�C����3Pl��<�{���C���8��7īj|+o��Xߋx����� ;O _��s���B�֫0�]
���t4�]��t�d���Ԣ�x9��iS�>�w�F�6#�o��$�+�4�L3�tT�-�m�a.w�_^���^	�H�l��B��ZW�X�z槸"|�E�O.�?��A{�QP���LK�
86%]bF�3�^�v��v���j�0�#U�9X��f'm��M�Ű���D8��L61����kUsȫ���L,O��V�R� ��B' ��,�����7#m|�
�1��1;��}��ࠊ��^�I;�+��"�k��˓g1�:�5ZP�U��v0��Ɇ���f]����Xa"�ZE�M�"�W4��EP���)l�Ah���K%5���a��d���+���+��l�	B/���uC��x`�"�*���#^�Žxq�II+��0�h!U6�#ּ!�9����σ�����¿W�u�67)��Z�X��۲���;]�0�Ի������m�� ��nh�L3�4�E^m@f�)�$�����ȓ3�� %l�����6Y�nK�s>���hs<b�� �rt�g=�]��S����5��S;��V>��`�G�kX9�E��]���-$�A@;A�R�N2Y���:�8p�5�Z�Ԟ��Ĭ�WO���XE:��_��B��c?K������S���5�}e�,(ڤ��`�(�D��;�?2��~X'�2q5��V�,�©��H������BSO֝�1�dE��1��.3�4�L3����i(�}�q��,�Ѯ�����=gGU,�w�O%����$�!
��Wt��3��4�O�`��,�~��@&�Me(̰��	�t�0,'�$ȟ�r�.፰*A:$��X�
T�x���F�&�Q��g���J����&�ħT�p�~%�(��)J�L��6��N`��{=*6���3����P����3Z괱G~Y�c�ە����%��t�^?���>�������(��%��/�i���:��{�8�9'��Ee�~��L���0y�<�b˪�rګ�$J��`��@�T:�H{]�j̒ۉ�]L�n(����T�~.�/�	�}8T�`�@�q�����c@{z"pPZUW�@��q2o~&��������_M�����#�^�Ny� w;vrY�����w�:��,G�֠v�z��pL�\V.@��@��L3�t���� �;T�8eS����Q���ߛ`�WYN��+����q�~4ʄ��S8Ź
�O�8�e��3ǓN|����Z�����޸��3'��B�x�N����I��ޒ�V	s�-��P�����g��X����<u��'���_\���2g�����Q�ħ�d�c�K�0�Du2�w0�`��ɀ��m��Y�B�=�,;��k���T�l��\�����Yз�"AQ#ϯ�ѯZ3�4�L7���m���[��M�]��ͯb=6������Z�̃lS����k!�N}<Qh.J�BY�n֏H�4@����:/����+�ܬ��e��b�1�y*�F��<Ⱦ�m��A;�Th8L���i�rjafUx��0fr';׈�
^�S� ����w �,ɾ"�5t��x:q�Yt��6t���rt'p�4��>�������vp"XtV����ɍ>�d9i�4�V��e�Ĝ���re�YX<c(.�)Atg1�&رTj�cM�b%���ڽ�¨�����u�nQ/���9�y(X(�[ϊ0��\�Rŷ<�'����c`^�Oa%@hR^�C4�VK؇��H�G^R}96F*�N�"nyi�B_juFTF��u�!�S�w�l���)B��7h�.I�z.�Xv6nx._�\�i��f:�(���Y0�yF��1F��M*�OI��õio@MmW�@�[£T�GQ��΀�����&^�1Q0چ�˖1n�8�����c]Hg0��O�Z��#��	y��{�)���|��ۮ����O��\Q�һ��4F��3��҈J9�:ҭ��cX#�{�yr�R"l�؎R�����L�װ8���d�C���RR�W����<��9j0���L3�4�L�F�<�c���i���r����n����9�?����>E����י��A䰺-ƨ�V`�ނ�s(�;
[�3°�z�R��l��QT�J��c��6,�x��G(�J�2�?-y����bW��Q�Jg?Uq�\����r�VtS��q�i3xä�����TGv<�.hȻkm���z�W,��G�3���<c[�mZP�ɚ�4�̼�	�N��R�]⡜�C�3�x�Z]*��P~�w�Q�uQϡ����E9j�&ڬ�. �JX�`B����0 �"�3�89T�v�aiLqj�b4�Y�x���>�����JM�c��?�#u���ݕ�e��Q�D��VF*���.Ϧ���O����L3�4��UI�7��/��Ǵ��F��s��|�m�>O�R����ف"��ZWyPV:���_NPp�0|ķ.b�����E	�jG\@���S�j�5_4��XR���y�	�kiD�)x���6��,m�7�q)?T����<�+Y2��A�<�"��,i����-���x5d�c�k2����q� ��ɶ�f�cZnf�i����oJ��kT�uZ4�����G�<
�b�-;\_�R2-˰�+�_Ѕ��Y���SiP�U�B��a�XU����[��FF��U���6CL�l1��ĺ�@X�%��7ٶ���0`;�7G�1�br�R������x]60wq0��r��I�΍a����� ��r������X�o7+�fN�7x�FٝK#��#Y���Ia��e��m�U_��v��,��!�V/8fQd�~F�,��T8e��|�59ANX,`D0f�`��J~ �H��L���������$�Zֱmۓ����
�D����3�ڡ���|��O��za�=GR�38�s�����?����棭�&z���a���0���S7(�U�3z������n �L3�4�a�I��]�!�q�F ���ljtm*2
�<l�]6�>�b�=9y�?��!���bVd�}^���)Y�:=0,�Z؛�@��05����w2�f�o�Xv�-��:g��/�����ɞ�I}��ׄL��t�)����e[Һ��O�'����E�\��կ�ʁB��S�]�G�8�G��O�8c����OL[�>�S��MCc�
c"���yӧ*�����b���ʻ�������<�9
�#�g��S�N'����X��d���)�7�U��o3�4�L3�����w^��MG:�P:��vYN�<�J����� �숝~oR?�|\׍d:+s�GU-Գ���C��c��e��-�C|�,��a�L�u�t�%x��Ȩs%̊��mY���Xm;ă�W�QC�[�0�����Ԃ�`>Y�mr͓,��,Db}9���q�Y(�s�-�oY��+��>��!����F1�8]�z+��g�l/Φ���Xہ�z�����Z�)�l��ц�;��-\����=nr�6���i
���z�cݵ�a t�^t�31n�3Vn�},���/>PF�Y��O��VU,7^Ғ�*�ǅK #,�Wh�/�m�� gٶ*�|'ɤ��5ðZXNjC�K�A+�đ�\�]^��}ޢ\gVQ�]7/#��V�f	����k��1?�]�^<�9	AG�LtO��7�>�#0���a��޺�z����2'L�3�4�LGAi-j�6x�9R�G������勸�����!�wK�P/'.�����x*A�tG푰�1�&���N��$�G�4�8,��[.V�W�@�a~;w� �Y:q��Y�e=�ׅ���)=D����<7%�$�#��ϻ��e�g'owq�Z���:[=_��0�ɂ��Zvm�.�3�L�I\q�{�:�MNة���VG�=�C�3}��S��(�Ǜq)������ ��	�6����9-~�����4��AWtp�H̟��I�	9H� ._�<'�f�tZvs��enN�&�~j���a��u4����]��ޫ:ȍ>C���1��+�Р\�O%��e��i��f�M]g�t��+��|�A�+m�N��݄�&����ֱ��iiפ�>�%gNѳ�����exFE�6��(@0��1�D��a,� |+ ���,%`�@� ��a�֭�O֡l,%hmo�9�0YG�y�I�I6����	�EW�
9O?Na��$_Nt��xP��eoɲY����"bg&�'��Zd��d�E�B��������G���8˙ ��8e˹6��8�\��S>c��Tgt�07���Q~��M�f�J�}�Q�����'����j��lv�.eCy�\��pѩ
�^|l]�A��?$ݶ���:�?��!�O�
��].Ƌ5�ð21��;y3`��VT E%P�Gǖ*�\Q?E�+7,"��A,��f���s#��x��E�$X�\X�O�uZ��K�e��4���:d��ۋ
��Dx7�JH�s�kנ}͍b� Ɗۙ6k%�jj��߀�N��i��f��4&Ԟ7��2D
��Y��
Iȕ�ʒ�����H��q24<����K���,�S����֤�t$^���B'���x\)�tn�'n�eC^�M��K Z-uצt��{~}IW�����n��O���~p�:=ߕv�
�Dg�X�މ�KIMC'n��9���E%�2":�)�c�bR�+����z�z`h~*����Pi+±.�j�ɋ����E��g�Jq�M8W��S~�p,z�E8׉dX���!"�]w���"��ks���}��S縍9���%�Ij�����i��f��i]]Yv���@��
7���>�𚴣�e;2��B1m�M������Tl(�+tެҶQ����I��ܩ��5��?�|FcLF,�R�0��+2o=#i,@C��%��TY�1 a0�[��}X�b�(��-�7_d���
A7�x �z��t���z�r�5�#剀1#���a���������w������9-'�v��D�؁#�t��f9ׁ�# Rʆ}�:;;��ӡ�����̺Yyb�th)(���S��W�p:�R�,H ���x�� c�y�2�8Wv�0I��ʈ=j�:b&��4妚4K��j������ �9�����"�ڋ6$�l� >S_�1V�i�	e�y_�� ��)џ�R�Mʣ���� ��Q�3�4�L3*���ސ��Ԏ'x=�ԁ���7�χLB�]�n*�sY*����i�U^���(X���N��nB�� �ʪ�����.��쾜^�~��;���n��_{���;�5'�����꙯ҟ�����/~���~�^8Y���k��3���$�Ι�d�_��d	��L���#v�|�J��t�J]�U��I��/q��U��o3�i� {�n1��9.�Nh3G��!r��"��;�C���y-e��S)|���ۆ�n�w�`������{��69�f�i��f�i��9c_�5��u�xD�����? �?xx&�&ʘP�Y�a�(�S�2/��@X��ao4bo�:L�.�e�[,�ts([���MZ4��8�]�H�y��p*���O2�H�����'3ƿ>3�FH�e��v��+��Ƨ8Ubz�1���m�u���紁��P�l�8����è��8K�y�h�I��u��#���7��j��z	���3VL%%U�ǥ0ɗ�t%P��=/	�3�4,��˪�������x��Ma�nP���k8�x�kn�wf塗Kf����@\{k<h�fK � �ǈ�	�ϙ	��V`�o�Մǅa���@�ř��1Rܛ��}uwF�Ӿ���L3�4ӱ�g��LK�ˊcZ��$��·�6w�ڥ�iW
?P:��N���N�	�z��ͣ��%;ȏ�}�{#NN'&,�X>j���3Gw�����]���E��}5]؍��U��O��w?��{�M������{�����}��g��Wo%w�-t���κkm��7�7V8�S�.�i\82څ���nc��u���p��%��ou������ ���4>c9�{:R6*�9>Ȧ�'�!,ѐ�krl/����X��� L�K�a,�:�����\��f3mCiܦ����/�L�|�$3�4�L3]�U _�碓m��i�Ӷjy�F�M�XՕ�C��k��Q>��e_�PF�r��
�Y��ͅc�˲��6���/�,²ݰ��y�[�Ѵ �5��B�A��d^�ޢ�P�G5�d[�9do����2Bz�9r�g.N�/.c���OE��Ŀ$�����=�#��Nc�g�6�[C�&]���܄q��t%[��u�S��6w� :�
�N�i"��^�iRR/��͕.��2'���;߃�9'�?�y��� ��qr��,/"�Qf��zS�C�N^,��4e��a�є��Z�|"���=�~J�:�m�db2\s5f�>����"P! ��A8���PjO2!.�q%O��?Ju�vbO�ͩ���-��
\�?>�@Mt�Je^n�W��^w�q�&٥<�+���D��h`ڛi��f�dtxkXZs+Q��a�c$c/Fc�����1��Us$�����ʊn��k�����]M�i�5���>��3fV�Oµ��Y��̐�jyq��Pk��F%Kw�F{��՗��?}ϻ���ߥ�nY-�V�\%zOg��z_]�y�;�����������~����Oҿ��������������bՠW��OWŭ�Y,WE���n�sG��\�°��j�a���Z�0�7	����΋�}Z�&i�,g,q�т9�o_(M��+%�b���/�&�G)�K��,��T��1j)��1�ޒ��Ϝ��!���}JS��hp�Ƥ������}6�L3�t	ȘȻ)�a]���gq��<��}-];����;څ�H����ܣ*;�d�3�%�,"�M
y�,����	%o�>��4��$2�i�|����l�V�a�P�b8�R���s�����rty5,{�rBj[v� ۈh+�>�rx�}����'~y����H�$[�S���v���W�v��1pl��m���t[���؁#��q��8��ilpv�z�=�jR��A��8r��k<]�y��.��3���z@��J��TnZʔIq����$<q��<��gf=�	��)O�G���L�:��s�w�O�m	��|(�9.�B}NK�9����a��K��N0+���C���s�>��ع",9a$e28�0P�iC�X1�$�C7�%�4��
�W \����[P؅{�1�Gܢ��9����L3�4ӱ��1JG�G�����-.��p�&!���\�b��\�	'�՛�$P�2����*V�������t��)7^�7������G�k'D�v�-Be;�9{�4���-��v���;��>L��?�/?�m���>O���|�����n�B��	�EK�k�U��T�uJ��h���Ex�5W�MkiN�fN�f�l`۽Yn4Ter ���t���#��dU�!P�@	��X��D�w������	�(I��T>����qD�3�Qrv����h���=4�L3�t���I�'��c��;mc/2�)��-Y��}�A�r}���I��y�T6���A>�,E;I�9�NE���ھ�m1	ց-F�W0n9�S"�3�?�<��-ȕ��d큁�ޢm1�m�Òܙ�E�u�-5�ٲ�������HqȔys2̩�W�Gx�G ��������W٧�?ˤ�#��P�����#���# �g['ܬC�^��Ii���8�@�p�.m�;ّ���:�wT鎟���$�������f�q6���u��2���5�!�H9%�Sf&)�I���3�����0�����a��yz��b��I�"�sT���z������'��	�b=�%�� ,��!��	 �|�䔺�@7z
f�]�����l�cY���b1�a'hӸb�`s�r�svbk��]����l[���6
�4�L3ʹea? �m�'�-�9�;���ꗓй>;�f��� >)�F����ʻ��&%CH�����ؒ��"qs��f���_��w���t]_�]rAe�� ���/����
����U��u���>�z��o,��=G��c��>�}�G?�_\��n����-�;�c�W���9iN�|����O[I�v�qT�05�� O�ݣxb�z���M^*+d��b`Xv�N1��YƗ�B&�ߚ���T4y�B"f�e�T�z��Ma���0<@5�D$��iG��Y	�O�ݜ�_�6�L3�ts��`��Ǖ8�&"���ݙ�������$V�ԩ�擁g	�§ȫP�[��e*�%j�� �`:o��� ���D�1�|i���Y��l$��P���-&�E�J&��z�2�ԃ�O�,b%;
��cF��2/b}��Ê��rm��C�+:G��	����%V��@Z؋��9��W�����s!VRMX8�J�nlr��u�τ��T�����7�Z�e�� ��*)犼�`�d���\��ZP0^NKS��>2��+ac�K>$/�=��������"�'e?�:��d��
C��,p����E맊�m�Δ��7_�b.?���L �Hl �<o)�;�J�ѐ�Pq��/X��q�Me|h�s�8o�6���J����4�L3�t���$�.���<;����'I�
u��u8�������B�H=���G�OIYFcf`R�Il��p��FT"k��>NK��PZ8!({��O��~�]�r���ϕp�F��;mxxok�2C�����ƒ��~�ᕯ���ƫ��>�!�ҷ�M�~�Y���_�ǿ����t���N�5�V�-�VXl�Jݬ>����>����;v���9Rn���]�����u9;˕	��?1���E�1<�e�s`��0�Vm,��$;y�v�r.�:�9;u�8�!Ʈ���Ɩ�y^t�ؙi��f��棤�eL��7�I^�D�u�C����M�V�oM5y�M,KZ(�M#�� �1A��&qAW�AW�e{F֍gT��O���o�~O��fo��E)g���̟߹�>�j6��F�'�v��!�9��0̄�^��*H�F�?,�����,���BI�O��R�#�/�<�m@�7{mbO>�>�0��5��n�P�;�T�2��+T(�Չc]bG��S7�TY��b(-��sgCgYp�je4o|�0\!A�+Uؓ+.Ѹc��i�+�UN�xQ�ð\�'\:t�b�;3�jFU7`\a��y��w'�D��N�)���
K5N�8Pp�,x1��N���1f����¨ �*$�q��:MY�v��K|���4d��?H����^�֡0_�r��#�,d���g�i��f&s*�hM\���}��:xu�������cݡ�i������}$��/��ව�l���06�fǅ�x��L�r��%�w�ҁ<�l�<�9i��K�~F�]d�����oI42��ɴ����e��G�_���>��}�>����ǟx����O�G/�Qs��G�W���mh��ȢY��U\,&8���d(��hq��Kn\&Sê��{Vv�vD�ⳓ8z��~�99>�:hR�u'����?y���¹"�dY�1�c0�qrxJ�dɴ��Ͷ���s�3�nu##�Ɇ�mT���YJ�i��fZ��s+����탊U�����qtROu1��о%�fo���s�46(�mPY�e���O�}Oڭ-Ey%o�p�i餦�'�����<R�Q�m�(km���9W��!J[�+ygy�S��bS0�c>aP��'Yc���mQ�ɫ頍RyzX�1�S�p�֐��Q͈"����H�s�=FB�� �r@��F\Y#6fFE]��dL6��Ј7��w����}>6�B%}��r���.�(�Wn�ֹ3I�q6IPw�7,b�?��ǻ�v��U�.��IYZ������FÙNQ�l���y�x�֭��x��v:Ae2��N���m�����t[P�R����H��{'�Km��F^���cbn��䅿L` M���Bb���`�c�I�Ҕ`r�>��8rŲ���1�rM�s��Zz��sD��L3�t��"ֳ�2%&/1Ag ^��|��3iX����o�[��g��
�M��K�w�3��,�k�MЂR��p�s�o�l��#p�v.�)͈�f�ګ�%#�2~�2�K`&F�m������Ψ9m����6}������o�y�����������_\�h�!lxX���i��z`��A�������g�F��ѿ�?�)z�{?�WE�-]�v�N\K-;�v״t't�W�]F:Z����>b%r���^��(#��0�-�����x���1���ݻ��e�<�o�#�K�c���#e�X\��K�������8)5W	�0�V�+&:o���S�uu�ͧ ����W��8���չ�Թ��vՍM�܎I�7�L3�t�k���{�6紞c�����A��yYf&���>�Q�*��ʓ�Ki�2m�n[몕Wuu86�
���Av���1�渢���sD�X+���[�i�{����f�Knb�Z._�^?�"�sH���3;Q�,���<�*�����`H���আJXj9�9y/d���Gޣ��֐�B1x�ќr�d�-G�߱ľ5�"O�O�?������W��y�H;�J����h�A�q�ڃ!r֌�
��0�/�%��Z�
6t N�}����LK��y�VX���<�r�J�M��v#̹�~Ym*���	�a��̓�����eB��;c ��A�sƙȬܡ��wP���S.7Y%��8��BP��z�F�a��r�:@*�� V���O�6Yr	'pd~/9�F�F9��5�vM���g�i��f*h�%�n'2��Z��/�#��%W�L�� �jZ���J�f?��%��e��1��3�仏ӆ�����/���o��\�#�m§oX磶��}��^A�
�{����dU�;x����C�������w�K�����>O_����ū׈n�-��ewL��Խ�L�z�߸iXxj�f�_�J�Dgm�1��w��G�C$�2�Ӱ����%��ܞܦp�#5ʤ<��R���I�����I�[V*ast��f�d���r��L��hnN����f��f�i�KL��'��c[����c�1�3@h�fۡ�@:�N#�w�����!��Y�1l\��4��φ���?7�<���ax�f��-�'B@�*6�ɶ�k���"=f���<EK�\�^@��F}Ǽ�Ma�Q6�ܦ^���G�D�r<�fб��I��h�]h�'���K�ep3����f����1�,�;ΆDX���`��,<'�xLY*�&�d ���[#�j�M�����2]��(Zaж'���,[�zO.F�$WI��Ұ��%���{�/��*�[-� ����<�BX�#M� �R8��܍&P1�NH
�K���8�:��6�?t��E붒���O ts0:E�4�L3�t\�uq�9b\~I�N����)�ŕ(h�F�Kcw_£F��S�f�"A��1�H;8'N;�R�dҹ8,�SI�½D�g��������{%э3�����W%9(��· ���,�;���+K�W�z�^��ѻ^������sߢ��/�G��,=����O�/i�9g����R�ھ?N����f�Q���ǈ.�����;����(�|qK
��۲�w�����ɜ�B��F�C�_J�	7���XH��O�ҫVR~�WrB_�y�-�l=���r4��S�y�~�j�fwJ�_�8���3�4�L3M��0����hv^�����`6�V�i#�,&mq��"� `aC��%��6�ֵ��c�R0ƺ��9��:�0l@��b�b�a�q9,	 ����a}VR�+l1��b�Y���c�٩����:��V|Rxi��̬�G�l��6��\f�j���y`郙_n:is?�l��8`�Z�c��q,�g��8�}������I"�^Eā<*�<*Ő��d�n�܄0�}���<[7��]޼���	ĶEǂ�(d����Wjɟ����0<.�&<;eۡ�U�w�A�<&O�P��T{�7�n�v��:�3ev��ŅݕCo�vd*�jb�L3�4�L����3�tF��������Oq� +��9�����6&.�`@(���Z��3�^���X� �+}�ߢ����c����ߡ�x9��m�hù۝��e�� ���ج��Y`\,K��b��R�g��,=�{��t�^N�x�#�G/�@�?�U�7�=N�|���OF?[�H�ۯRs���e�Ҭ��X	���V��>�I�N$hb#���s��Ģ�TcjP������$!����X�I[����r��;�?�q�1��(����0��R�˴����X
sȧp�Ͽ��hw��+b���W��_(9Ҥp��F��f�i��t^����]l��J�^��g!ش�Z�[�*�N)L.���:;~>���
dC;g<3m4�l
�5æ�w��8n�S~��	��e���۶��p^h8'��S���l	}]ږli5%�@:�����aN}�r�AnL[�ay�Hl��N2e{"�c^m�!ch�ġ�qf�i�+T����ϣ��gՇ�++4�R���M^l˻s�L� R�m�M�}���:��|��$*�jKI�Nd�\����Z�܆a�?��ɥ�0yl^��ZD^(t1�0�s�KߡY�0�%�1XȬ�VOq`P�5;�
�..�I�6SyvzYN�(F�����J�l}�EzG�Ay�GB/Y��n�x�	��\�\1�ڢ�CZ�ې#��B�pY���<�%x��f�i7t�`=���h��7:�0E�W�L�`A�La)4��(�2f�!<4�[��l�1��t3�HH��q�Yn�k��5�(��s�P��)��2|_�+t�{�O��}�������҇���t͝�D�Α�,xtעx |d#������|�������pH�W��Y���fA���6��o���[��?{����/��>�8���H_��t��mݑ��*7gt�4�%[Z4'�]���Ξ����x�G�OL�+��PjA�ѧ���ԪQ��t��i.�8�B����q���X���/y��0���T�T��4.S�R���St.F�YW"�q�.�;�\�,=�L3�4S�p!_G׻5��əw�x��'1���iL�5��kt�sv�2x�֔�#ٙɌ῾�
�P7��{i�J�aH�H�O��0�xj���<�~���g�=�{�-�j���Vf�b� [1�B���4�����j�ʋ�%�U]��xeJ�R�Y>�DrLO���:p�[�����f�q�؁C�0���$y?mTS8�0%/�!A�>^Vm�tQ�d�B1P���Iy뜬�����
����o�O�0Ra��ӫ^������5 �S��$�ڏ-G2]*_.����D^ccw$œ"�G�B����y�itl�+w��P/'2�Kl �g|$w��\�4!�t�M����4Ύ^!�H�������2�\��)9�CT0
�A���4�L3�t�T_+ұ�.���+��rS�q�dct�݋2c�@S����vB����Pqda��t96����5�
�|B�ݩ�?!�ˬ�'+,�R۶t㶫�W/>O��?������_7}�W�Nw]�%�{0Nr��F����ۧe`k��>�5��۵;�#Ցz���գ�n}��+���������_>�U�ė��O~���O~F�Xy}qJ��N��d˳U�pE��*��E\T�u����g ,��.e˩��v("g�tv�p{n`��dY$G���ɰ�3��e�,��w#a�,&��e�s\<]�l�m�O��cQ	�4�L3 ����tm��AG�;�v���)�[G^e+7]�Q�����s��=�\�y�s>x��?#���"I��oڜ��;�pta�����k��3+OKp#a����(�x1e�l�a�E�M�i�-&�)�Y��dU�4�w$�si5{� [�c:�\��B���߇�vX�%�P�F��!o�(�d�U�ݭ�F�{��f�W�vk̦���`�)��=�?�v.��������������w?7�2�Q�Z�����X�� �����ML=�@������2��7Z4���O酉K��sdp�!%�&t�)K�?|vVȊ�\'�bP>� �����w�I����.�ħ�/.�� �7D� �d;0_^�wJB+�,$柮�۶o^�-J oGS�#ޭ�Ӽ"�j9uxܶ|�8���f�i���b��y��څ#I].R��q1�� �!��H�b4d���^��r%c�puI�H:��ޡ�;a��vB/�4����6}������O|�~�mo�w����}���j|8��Oӟѥ��(�-��,+�r@�v��ҝ��{d��Z��Ŋ���}=����?~ϻ�[?�!}��/�'�<}��ߤg��~qz���)���劷ev��|�"��k�C.\�5ˠ>�����$�V���'�_�MXMe�4�=���cd3�� �ᘰ�@�Y��I&�)]�Ydr<	G�?�������t���43�4�LGB ���2~)�]M[.�;?�qXޥ�=��Zȱ��B�v���KFF+U�i�>2��b�U���i`n�dV^��ۨno���UcjJ� �x,l1���bH�v(ѩs���!s�:����a9$}z�O9����7����u��~5�1���:�De�9�a�/�x#/��iݭ6-��2���X��U&�~�0��ZS�U)�xV�Mk�)��K�	��آ�����j�D������|��N�#���x�|i�|Սg^�#�o�����Ι-����]�Z�nL�p�8#�N:I|A9��מ߇��l}*N�@T����${:�� 	܆{`I�<&0�ip��f�i�ɴI�<�#��T4z�.� ?ڼ~r���W���j��q��W����=HΧK=1`����ʰΩ�]�_=X�e��]7r�S�W_���_�;]Co��^��;�A���x�n����g�{5CF�����	%7�<i�]��Iq��=�Xw=p���>��nz�C������O�3�ԗ�L����O|��܏��?�B��+���xq튧Ūދ��EWjんGlT���|��5R�����H��C�썲�@�gG���&YR+�uDaz��/�L`_��[��^��b�V��,���Mq7��ob(9�[�d1����Kvt-p�4�Z3�4ӡ�3��ҕZ>��H��Fŵ���N}_S�P�ڈ a��Ҍ'��u3C�׵��xc��C^j��j�_�ϱ�<�=�Iyq�C�(`�TTy`�Gkb������mUM8�i�`�T��<[u��T�"���PNj������7��â-�P�/v�Pie~�H���t��н�ƺ֤������uC�G���fe�A��+���G�	9!$�������9n��~h�0��K@���0��<՞�	aS���y� �*wW^��Y��ɥO��d�Yɧ�U�'4H�9��g��Kx �	�b��8��Y���FJ�޴!�p��0+_{�k
��U�޺��ؽ2�8�������p�'j��dO��6�<W�9��g�i��fڄ�
�f�Jc�u�!�k�o	������mi]S�;$;�G'9����.ۜ��
 YB(�|)��J�\G�j���B���޹�ߟ���_,;G�������w\��;o��g�荟�c�(�O����Ɨ�E����Co}3=�����k�hѝ�֮J>�x:Gw���T�;]p� ����ar`F�!Rwh[��K�>�������v����N���O豯<K��/?K�~�����KW��z;�X��ޱdIg��}u;��0,���p���tm��[ׅVNƙG���p*����O]���_�g�Է�����ީ��O��1�NA�/�D<�^��^N<�;�bAQ�&��x5g����nz��v22�y�!~d+�fd���5�L3%];�:��zr�[�V
��m>���v�@�<����m�2�N+��e�yN��b楚rJ���&cв��J�*П�M��O�Mŧ'u{�����M�CM=�!�[t��Z�#8�t+�}F�g@�V^�M��B�k�#�#�����f;BA��x���dZ�v���	�Fۼ����v���qW������xQ�'�\	#�e$��
wI�E�A���*�lKQ9O4���$JY�f��8�d��ug��x�q�u껉6�:�O��|2���N��MC k(��lܱ�Z�Y݋��>}�
�,�����}��!��J�s��В3x�?�	`E�ܿ��C�����8��4�|�j�q���A���C�1���}W��PR`��a0��5�~x�%Ⱥ��Ea:�L3��tR�8���z���؇܌�w��إ�)���2�?o�����.q� �4�w��ZS�>�`J]T��F}��35�J=N�*�x���*,��W��0��X@��w���	�,/N�9i�gg�>��_�g�ݣ�>���_�w��z���#���~鶗��+W�����k���;����>���e�R`��{߈Б'=�D�}���_������w�OO|�+��?�E��׿A����М��.�9[թ�Eӹn��.V��&H;������;�¸���_�	*)]Z2u�M¾Y�I��:�r��{@}�,9�`����Je�S: _��yx� �	n�k�:8|�t?��S�����!*zO��^��O(�&#�9�%���&��L3�t蔖}m�����@�r�6���㹨��Pfǽ缘A߅��5;���ޠ��	F�o��I��q�p��,n	g2L�&�JUР��Ԩ�.S�gZSBX5����xpF�Z�Ny�?�q���|���%��(\o�`0,v0�E��Y���&�-2cuo�;�;��'a|o�ˈ���u�G��'��+�bb͝gSD���&ӱ���:l��a:o���P��FfʟE�it!��úX�F6[��,�v
��/�(�O~x)�z����d�EP�A~ńѽO��qLR&P�,CM�)�ʮs�Z�=��S^lg|�t���/��iP`�kݰ��r�!�hۃ4�V��,<BQ1H$ʱj_��� ��'pȱ�O`p,�g�O��এ��?��̃�푁Ue7O�GK�T�����~��Nq�B�]�K(
\a��f�i�ç]N�N�;���~�t'��Q�=�ܠ-�b���[C��>]�n5o�J-�ۆ�aڈhs�J�6c�&�i��u�h��R�=�]6-5������*�w~�}���}�^��O���\��z�����m��^M��v-Viݲ�;8�8ZR�����9B�B������S�t�AT69]ߞ~A[�	=|�k���_C�}璘��G��'��?��c���~��_����)ъ��ICMw��"#M�z���4:7d95�а2�L��������s'[@��C~)8	}����G����)�o������k�რ��^�1��@��"+��BN�i��f��⨀n�����xJm��E��O=8�ԒHYW��+TX>�ZW^��s�
������\n�%�i�\�bW�¬[Z��!�O��{�P��6+�-��V�I�-������"�C=w��� 	ST��sEa�!���	9�Tٱ�/�:T�'>Ɯ�wA�	�E�Ykw��:���EMV4Ti3,{�tw��J:�Ю���V9!�ڈ���$tFRO�l�@���ód�]��A�c�Y@��$]�@����5W�\��Q��xgE���%[��A�&�����ި�j1�������x��JH�v� 8�[�D]�gvQ�[4���yY����fj���`l�d���eǙK��q��f�i�åp�@���x&E�C�mF��ὁB�E�'}��T�/�5�M� ��,)�}�3����c��.A.���������Ks���q����t��̙��=����O�^~�����}o~#���W��/��׻�PK7z��s�=i��n#��3��t��͸����i"�>����^�o���_�g����'�@�z���g���5'���)-Ot�Js�Vuj-�E�g�,��0��g��E�Y�ic[��	���2����x�J��Z�*� p �����܋�B�	Qٱ��tE&Q�m>yP���1V�VX�?@�e �tK3�4�L3ݼԝ��L��{�&�Mƺ'{킑��J$�ġ�^L�0a��S¦�`��_i��+Sl0c��m�15��g;My�b�m�����+,8�`eo���Z!w�VV�����T�l�	ɝ��@6�<Y�s8g/̵�k��w����|"=��l4���ܑʄ�9p�)\i<{���tx��SF�4�g�:��s�g%�W������Pu����7��ȭ��#��@���� �;��:�J�� �o��.'��R4���u(7R\�X1��v�aN�h�EY�������
G�W�+��	�it��}C�&�NJI)�o�| g�YH{��y(9�9��Cx��,�S>;;�4�L3ݼtl:y��4R�̴=I����\y��}�e��h��^�����D����,f���'qP�j�]���N-`��.^��m{�����GmC����3�����|���.z�~�~��o�_}��t���ɢ��$��Xr,�?��h@���y�Ee_�H��|p�5g��+^^Mo~�k�o��}��o=G����/��4=����O�KZ\[Psz�kdZ��bI�h|_�._wA4�D����0�lR�E���a�_A�Z�r�#$ey#��<����dO	9���U.)� �9H��-O��i��w�ѡ�[ZQ����f��!v><&9F��� �5��7�L�9u��~~H��X�Q6��o�:��G��5T���ѹZ�iiڗ� ja�� ��>v��]%�����I�M���W���7�ɧ���ޙM�a��%6$$��X��Q�	��,���&���M�Xw�xP��rJy�8�����]��cs�IvyU�1���뾫�}�8Ġ�����!J/��1F{�;~�}$�:G�%\+;��G��˳�cs�]��ο!���N��%2��y#�O(�r���b��֧���f0$�cŵڈ6|��6�k����e�����Ni�ٱ͡h^�=�)�N1����N�٥ګZOL�e''�Ә?�h���t�vN�y�iaLA��� ���Rs܆��6���ǌ��M���4�L7el�;�Q ;$!�w`��5�C#��ɓuBMI�vk��'�L��p�v2QFژ���z�1;.P1f�e��˒�	�\�����#�;'t�������mޣ�UYWW��N��r���)=q�E��/<M��Oћ>��7ѻy���W�=�\��fA���P4�<�Nt�2��)�e�w�g6V�����G��nw^����Ƈ�=oy3���>O�~�)���=��oѷ_x�n,W���[��*ߓ΁ey#`�Ω�s�]���(	��x}b& !�+P}೘R]H֏j2?�?^���N���œ�|D��T��5��#�Wa	�<v1r�>�YF��\F����B^"p������|��J�bǨ�M᭤�o5�i��vI�T*کӝ�/2�j�ܒ��v6A����p��퀴q��1���ʰ�~���lȁ$��U��B�	��0���h @[���cg}>I��b��o��0eY�`��߲%J$�p��Ř-��$}��aY��I,�Yb4�*>��n=C�w�oo(בyUh�kL'"DVl�wݛ���mޗ�\��l
m3���p]�́�x`���w3�΅|ҹ�,�/�>�6���>2XT�F��R��]�����}�8���`�q�A�o&M�z�T `B�&�8�6��tq��s�k'�����8�ҍ��AW�S7��w�$&����E]'�r���N�*|�H�1:f���!��e�;�q$]��/��#�3����퉏����g�3a�����,���f�i��&<U�I`0P��+�����ӛ �:�h۫$w����5H�)2���B���0�S܁zGцw��cOZp����&�w��#��8�.΢h�]�Ԭ�r�
�����ON���O�������[��_{�A��[�H�y����{��쌨]��0�#=|zA}�!
'u�f���9>�\�w��AbK�kV�"H%�뿠��^�����ч������>��/�?�E�x����*��]�[O�����Z�<�������m-I>�\>�#��:���RtB�+v�Vk��r�e�ɘ�uYq�R+��o�q��,�Pͳ����+��%{�d����#�����w�
���Ե�Uh��f�i� ^Pw�؃hw2��Nz,�ߙ�CRu��5i}D] �ίOـx�����vU΄������]�e�!]��x�����6���ՄI���M���6f�����Vn<�+��-�Hg�b��h"���݄냧�����9)�BQ�$kYd?���M9�0�:0$��/@�^wж����>Z'����մ��1nb^ہ�/����c����m���/��B�O#vzDd��*�OTΤN~V�S�2Z�R��� �5y��Ö���),�]H�^���q~o唺[���LwkVH�8�A|-LP1fЃ2�_>�J(;9!
,�������E.Up����ϳC��}-�5\n��cI.��
�e�w�����O:� ������$b�&�(�{S*���^�^�i��f�,$��[w��O�t�i�/l�$t� Q�F��ȍ��c��%6+;<�#|T����r�eA�?�#\���d��jCgW����O���+O?E���'��;^F��A��=B�<� �}�mt���a�e��u�s$|9r�I!���1֧��`a�>�x-V�|�(�h�\��w��~�������wD�)���<F�����WV\]�J�ӦO��-�m�}��Z�S9z�Oѭ���*����Fo3s��gRV��V-@F�� ���)B�S֔�̄�ȃF�<B����Y��O���B�-��֜��`��e��f��Ih���.ͼ���8t������fc}����d7���N������ع&1�~���e�Ę��-�U�F�<���1d �p�H,�o��\��Dw�pТ�&�X�+����b�b���^
�F1K$��]M�;Sʃ��sm�A[%�#�-���U�47���&{TsQ�6�A}�7p�p��A��jGM�z�Ɂ˅GG�z!,�4φz}�sy��mj�,$��5�Ȟ�eXT��3(�1{�鰮��hKf_	��S'��gJ��ë0~k=�MG�3��̛Ǹ=yф���3,�x�ZG�v)=��r��԰�A���YQ&Z?��@�\��=xz��˰�	*�̑������S!v�)�X��4��>����]�]l�@9�L3M#K0�Gc�]+���;��L�����!�`�Q�wcWG�^���7�\�� Rl�}�k8T�y���"����Aݗ.�ET����������녺bNW�b����	=��3z��'��z�����w��Az�#��7��^��k�ѕ�WW��u'hEot�� Z�6�߷9n���S9V��-z^;e��W��=�{�����}�=��o|���cO�'��u��Ϯӏ���K�)�����w$i��W4�$[t��Ӊ���,��A,��������S�r��|��\���q"�D8hO�|��_��L;�n̴�K_s#�4�L�J�\�]@�]�j��}Qy��~�M>�,��{�.p;�N�������^4}�2t�N;�j8�r�%(��$�L���;�4xʆ4~0V�$�/ �Oud����rNS���O��T�O��g�i��Pݶ�K��\��t���� P�����yRJ�3\.��w�a��~D%�EP��<��XxQ7���/��e�7�\����wע�9���W�ȶ�F�C�!�2�.��v�X��o���q
�S���B��UU֤M_�Z|q��A,�1�M�(�#��Ͽ-в�4Wyf-�N}�_��/.�b�4F>?�^s�?�Q,%�1�K�����\�*�S҆߸\j��)wA�Vjs"���< �8Y{T@棛��G#�Q��)3�t�Pb%�弡�i�+�=�Rߙm������lG���/c��<���%�.�	���2r���	a�2�%��4�L�HO����\ě�AY 2�̫��Gd��3a^\5�(+2֧�!����X�v  ��IDAT���b��B`����Lg)������b}�'>BTl�T��\~�J���0o}��; ��>m���s�AmT�y�\��O��U��ԟ�qr�B{��`�����>����|�t��	��/?L��η�;z�~�m�v���e��s�X-�,��·���&��j��|�sIW֊=���;�}o~;��-o�������/?C��g�?������ۮ��U;��(v�;t�����(��$��^a��2��x��su����X�q��4>�S°8�T�M;�B�PD)!��r?����~�{G��-g�-�p����L3�d�%�+�Ӽ7��^�+�wυ�y%쯼i(}-Ħ,�d�!m��/�����.lcܖE�M}�eMؗvL���8�;3�l0N��塌��<��ɫ��
.�]R쏽��'�ZcͶS�h ��Y���g��O[�����ͬh�)�C�#e��@�1̙!��<����>>��_���O��Yzt�<Gx�}?��.�..�f-�rx�^eg�q�������u���,~^F�w �N��As4N*�N}�[�\P�m�U�j�
�o^8�A�hsF��cM,U�b*,HN�E2:jp��0Tl��o��Bo���\�6M�)f:J��l(�����y�-�����q��C�
�r��?�W \���K|?)�����:݋���>�Au�A��FwW�[��)xb�տ���n��nLwF�ư���p:�ݚ�K�=v���3J��8A�l�k\�b5qrs8��cė;;��y9��f�i�a¹���x�Ҝ��껅����ή�Ө�3;���*!��;��{�E!��
�9Fs=����#k�}����d�j
�n��2�k妔Au%�����-���ī�)M�,��R�� bz!(, ��;�=X��0;�.O��Yb��#��z���Pc'��J�S�~�'1��q���)�W��*��n���x���'���ﾓ~��oz��k�{Nnt̞��9��/z''9���]{����`�8��R���/���ú�Q��Vz�����M�����>������>���Џ�]��%��,��lI�$��-�]8�X�雲�8臀/ɠ:�r��8t<ȿ���r&�;��WQ��|ʛ�>�;����_�~�����k��S�o9�B�i=���RG�u�0(��8�=g���Ik�~o+�[ynBzU���ug,����7�X#X��s
]'�4��O��ׅW�ۗ�������6�F���׈���&����e�P�+��ӊ�?��GM:T�;B�l`w"L {�y� 2��Л�a�[��E�/����Q䗯� �VŨ���:jn}�I�A��S��X�i��� �s(?+���/Yg�3�0i���x�F	��o]��]4��_S��r9z�CЩ��fV��^�}������6P���8i���8?��.�sޕa#thv�@y5	#"�.�	�+��(Y��!˞�Vz�߶�&�{N������.a6D^�4�c������&�����]Pf�8��}+�=��I6?���䌪���ŉ�C`�ڞ���b4��N	K�Q^4��p�۪F�ȦÆ�Z�����A=^3��Ք5�3ӈ;�D0�"���m^�E�-%��[+.�gy<��7�,������vDlP�h��m��V�~4��`�p*\��gv2��3�4�L[R�E�)s��� H�$�R��D:ϿCR����[e<3�P#
��q ��(�_"7���q��%𓦀�I� �"��G?��՚�[�v�N��+�dm�;Ltq��[���~@������ԣ����Io{����G^Oo{�C�����1���k��Z�E��a��2�,u����r�X�ΎC�e��V9\k���W�?�a���������Oҧ~�z�]�+��o�M_����}�l��Ri�^�)�_���$i]���Lce�)��il>8��BД"�dKKUC;�q�:ֱ���s��.�r>8��~O�ZV��ȉo���pN�?�1�1B�\tE1�>�f���i��(�>�wL �u�R?.�h�!W�'�z�t|�Ry�1bSeu�q��3�m���YfTU�b��7�P����6�F��Q)�g�|��"�hAg�a�Il��s2B��8xU�wX���i��N�!N��N)�g����8_�S�8}�e�w�r�����`��f9o�S�m�iWxe�+T���(DoǦS\t�O�0���˵n'x�-���/=�Ŝ��~#�9Z��F�$b*�ji�	 ��ҫ����I}$��$/����GBx�����I�Bsa1��@DYsYo�wX�tU��G�?������O�fW��8��K0�V�\�h�;��/y�^���0݂ō�
T�F��4�$r��3�4�L�G��s��E��=��n�L�`F3��*�-<|l.��������+m��xVh��sH;Iɔ*�+�O~Ӱ
���\��1u8'�t��p:G���ZtgbxjV�:猳+���܂>w�E��矢?~�iz��k�[oy�>����ￏ���JӐ;k(��m{�݄"�~����H���6rQ�rħr�ݭ�$8���s�=[��O���������������?z�������VZīTN�K��r+4��=R_�F^)�.<�5�`G���`�])_�������\K)Y�<6ϓ�!�N��ڷ�&��7d��f�i?t�3O9��ku�W�_���9��A���ŭC�.nB�M ��B�5�rY����G<�N2� ⟑a������9Ŝ�k��N�#��2õ��UQ�V�m�+�k�t�zrY�eo�� �d�)��M�r�/������<8;.o��N� ��#Q~�_�uO�Y�9��SG:[~<��ph������wS��8,ҤHGAIyz$�w(>7=|G&�����{ԊS�_�ǷIcu��j{	�m\.nyە�_)mh�6r/Ta��E��D>�9#Am�5Is������8(u;� �@"�O�՜3�A����\��E{'�3�H夬�B5�S���Z�YP�G���jh
|���Tl|H#�T'N�0f5%��v�L3�4��tHG�oDj�ܬ.Y)��V����v�P�O�劯�@u� �J2��%�ǻ�"�AO�VI+IF�9���H-���B|����x��XV˿��^P�n���vD-�H'}~'����5z�7�č��K��|�iz��k��_��>����{��9^u�;9�ڳ��es�_{��v�ʥx�ҷQ��l\.��X�/Y������"���H��qW�������޺���_���]��S����q~�}r���R�Re|y?-yW�T���c�{TrR�Jt9�VV:L�ys[b�x�r�$�|:Iyd���3�s�g�i���]�Ƈ��6'\/r�HB�z˭���s��/��eaS�2Β�P4�� -i�����������t�@�A�Z�zNPɨsg]���`�&�вUa��6$��2�ΏMz�/E��bqien��*�:�fo�cGl�}v
K�,G�rO�kmv�*&ͥܨ�F!h��򈒫7\�����~�|hz��c��F�&1Gz�%̡��r�L�������%��=��;Og�4\���x=��!"����3�˚�y�n߿CӶ�x񺑒�EDP=�Y�P�Jg����e^\ ���5z#Ҡ�(~��9�{������u��8ƙ�&Q�ݛ���
k����[.�A�0�d*��/s�z?�VP��^
��c�9O��)@	e����=�;ָ��6a΍%��������1�(Wm/]ya�L3�4��<���Щ�O䪈I}P\ǧP�[���æ�k�Z�]j�_sX݇�?�o�w�#|�NF,�x�p\��Ӹ��RB��2u@��#�9�<e�۝v��q��O�p,��xm�:_��9N,|�f��dA/�~?�n����>��|���/�������7��>��[間�����[�����e�����<�I �*��X��ĝ�ď�.�N�/��~�#�����gh��O�	��;���k�}�GǸ�)N� a a��s"4Nϙ��0B����:$�살t�r�P|�Eڞx.Hk�Q&�O�%����J��f��i~����hs�@�Og>-R9�e7�ݘ���Q(�g]� 1�u���xsX��ep�����M�T%�Ǒ�ʸ̤��9�݈-ƒ����s��Alax��жge�#Mz�km�*��jh�)�s���SlU-!�v�βD��`�蜀B�`�̗e6}�'��k�	��<S)y�Bkߒ0�k�̅�*3mE9p�qOqP��`�q�<�bP��o�"�IoI����p���V
ΐn��R�}Į�Պϡi&�I�L\Ϋ0hbY�`��F �OW�D�=�;+��@�y���Mz��M	#�,k x����N ��������5�E�a2�|�WΣhT1�޷f��:lq�G�Pj/c^�1��qx�<:ie�܅z)Ez2U�54��/<KS�C�	�#�}��'0���t�6$V�y.~�Yd`�u>��]�>ι���淙f��N����{��f�a�I�;���k������7�^R�]��7���B�%PUv"'�e}<�T��3��q�}��@�B��g%��;�X PB�۽�q���;�@�U��(b���1_/S�ƏE�̀Ǣ���^�׺�~��FcD�e���e?u�l�Ѝ[n�Ͼ��ǟ�:�oO>K���.z���_{�+�W^�*z�]��;�ܲJ{}��ǣ�s�e�ߝ�霎���s<鸊���eH�Z�s�������G��p�E�W���1*��Z,g|Ͽs�p������]4�ȒY2s0�f��$�y�Z�9/��5����t���k�ݤa\�w,U�O0�L3�tl4����]����}�k���P�L�U�P��� C}|�_ue������
��E#uY[�#���3�3�ʳ5�B�S6(�*x��\�e�4���Oϟ�1�C2���N}�4��;��j��-����)x0�2�ldw�%X^����;!�O_��Mf�,�)��>l?��*� )�1m�U���>���༪'��y�PI5=à�2�jv[|vN}ڔ��m����f_�ǝX�W���b'pE A$�}�Dq(QҌfdk�x�猷��A�~��w�����s�#�aF3s��Wp �� �{ow՗�\"2"2�[�����~ܮ���%r�Eddd{�ʾ�*٬e�q����W1Q���u��N���qh�����ݿi� �@�0Pˊn�ކ5�ߵKpT��8�3���˦Bpe�̥TkE)q\�_��}Ks-��y�5�{��ĝ������9����Ъ<��J`!G�7;� ���y��dI[mʍ����?i|���E�YZ��@���oz��8x&�&�d,�P>Ԟ6��_�	RM4�p:{��,������$�]��d��)
�JM�C��ʕ0�5�Lr��^�ͭ5Ek��c���q��\G&�n9n�~sc͊񪬳��ROE(���m:8�
��^.ۖc"4mK�IK�����f�\x�Wo�7�}����Y�������;_�/�N�V�JY�z#?�$�7�h�
��Ew��F>���]������Ń9����6���;����&��Ε�u���X���bc �ƈ>��	����x�-)r��]ל9�!x�d{� ������lMtn�KF?�\u���ѧ�u@�e��qki��~��
��S��m�KvZ&N�kLh�5Dmapf�gm��&���[������������r"=�8�F�C'�=��ΠT#��?�F�P�!������o�|�lj��EU�P��t£�=��%/V����7�6��O�a�Dg��3�H8��mNGl�Zi�ŔV��������L8���>�M�M�j�a�eVy/���y�kI�Z�pQ��k�UÒ�܂�N)��|c�_[FmϧNC����R���~Wؙ�8$N	~�LK֞Ų��X����g�eɊ]��]�YV�t�| `�<��N�u��Z�[���aM��L�VP8���T�5,9�$�9�Jj[?k�"�ָ�p��yp9���������D�J}��Sm��~�Jp$�=u��s\�J^�ea����hCU6�B;�I|=;�n��0�T�^��ѵ9���6P��=k���!�fT�t˫�'I�|]H���H��t�17�q�x� ��j,;���Zx��=[�t�v��_�~�����7^���>���<d�x�L@L�.�I(q/VsA�s3�s�f��Xu���V� 9Q6�qU��G��Lj�<H���^�vA� ��ߋ�o��:��sz�F�:v��-�чDX/]�m�j��JM�К���26�D�髶6K����B���2�]Q8>�$|g��D['�� ;(�#H�G�@o��{r���x� zⳅ��
_�s���n��G�yL!���twa�FGEmaU9lJ�Ց�i�R)w��t)��[f��rM5����A�������7��[�� o�2�ZNYZ���^�¾'H���3Q�J]��3� �[aR��W��^7�7������^ݣM���(���~K<Ȭ�2��H	7�{�R�R6�r @f@���t����@���9��"�K�����L�-|v/�p<�]��.t(A�Rf]5gT,��-�7 �Ҫ�I($����ȂTWć���%zЀ"7���/q�#q\D�{#�1���5���8u��]�A�?�s��1��-��AX�cD��o��O4��G�ûxkH@|�Һ��1�}���}���������h�e���O&"2;��#��*O��j� 9�- ��C:mg�Q�N<��T�EC���Ӵ�{�3�h&gU���lP�F�磣�x]]��ސ�%1[��<laf���7_؇�|���>�I����a�8���^��$v'�y6�'	�6�{��Pg.7s���_f�z�	
mn\1������1�Q͖�L��T_$�`]�_B.��DP�@^�0�8�9���1�v�3�J�֏�!�����e������O{&�h�����;�� ���wۛ�2$�^���;3�GӨUO1���h�v=��W���5U�|)w zT�A�TG��Ox2���S��̶N�O��	�Ԫfh�,,����ߓ���wp�?M�]W\��Ϙ�R�ͦ����������R�O׉O��Ro���@|NB&� V���?t�\�A�u�\�U�T
;Aǫ�Q��m�B' pb<w�m������1�А���甮ڈ&#��4���I+�����po�J{@Y�Q@d�:��h �Sd�Ad�La�3�1���Ңm���P��\���X R����b�֬��C1�0P}��C�����\�mO��7�U>��A�F']��c���R\`�ny�'�ծ�+U��M���9����vwo��?q��U�Y���X �Q�+�Eo))QC�8��"T��?X�49KM��`����`�A�LO��N&:����y�|,n����
�-U������!v����6y�g�mOm��Cù��zc6�a$�(�P/=�%�$������`^���yW�3%��gT:�_T�r�"���'w�.u'S��o_c*����OXe�n)GS����aQf�@Nq⸊�m����բL��\��hP�^�kV��\�/~�����/|���=�]���*��!̖�����N*�a�E#/�]��z��fz�M0���h5�/@cX����P594���N�69V=���I2Ċ�4�%5R��m���r��<JOP��&�Z��h�q�2���!=M��������7#�n�L/ƻ��<7�=��*�Dau|5��h\��R��ݵ&��0=a�#\I�h��&r�u~5�wI'nճ�\ ��p��gH&n�xX�܏iazK�0=Gz�Q\Zn2C6��Ze�$�	�ċD.#�:i�m�3�(N ���B������ �[k��؛l�K���T$
QP`�����g���5G�g��W��|�'��m��<]c�
�ä�<.AS �5��uO�8I�3�H�F�a(0�'X@eɢ�\�̂��F�1y$�]hA�k�''}�B����F_����j�;�1��ؑ�%��R��ʟ�4��M�0v6�*=��;�p:�k�Zܰ�(�R�J�E���RW,d� �%I�U5�p;[*�W���<oٚ`�����ҢMYTۮe����K`�K��?�`B}�4b�d���TJ��I�� �%�pԁ4��Ηܗk�S�� �+_�-K���D~F���ż���e��R��>x^�����9��]�qN���m�c4�Y�h�nEI�b����I��wM4�n�V�&�89��񱓉k�P���v�=��J����:@Qu��L$)�F�gʲ϶����qnC�����FL����l%	eN:�i4n�l�G��a%D�g393~��_�߽�n������D����m*���^9�Y{��Z��?_���S�n���.텅������.|[4�׃Dsl�����8�a�k ��.�3o����o����7�m�X�A�6[&���Ը8T@��-r"���	�G�ir{�JGH�ٔ��d0�ڬ����o{W�
=������ 5�����5�hX��k���a��ҹeFK}���&�h�ݢ1�~�p��֎�Vv�����K�� 	��&Zgr#��D1�AWjO~�������9E�r��F])߃�U����acc��S��b�Ll��`s\��C���i��Գ��Y��L8$.�ﳲQ������ϸ���U˚���X��o�L&KX�qS�tc�;BC�(�4��0$v��`�I��k�C�x�)T� �P�`��tl����G�ϓe`}i�a,��R����z��̒V$T=ͩ#u��ݥ�+^+���Ja5^/u-��I�K��i�B�_� �7�@���g���[�DKqmL�p�:,�e��j�aϊqUu3j��=��R�X}�~3&�bX\�e��<��x"�?���5�;�����[J ��Z�U��O�?.甒� ����e�M��\$�Б��+>���0N�)������G��r����:�D珺��q�d�76H\9�
�1����刼'�I2�gv4(��l�@��=�'�V5���mJCl��0&�i�$��R��H̢,e�K�N�&<�G�Ӻx-y_���ӂY�R8\�u�>z����	_���~/��7��ͼ�F�.�HsgTa[��!�<A�n��	a�ðg!x��ή��K�.���<�4��kG�^6�N˺�\٘_��C��Y�b(&/q91���r�ݱ���X��AM\f�z2^�(9UG�Ǎ��_�PE��P0o�L4�D���ډ鲠����l���A(���t�p쉕�&�FC����V�ŵ����OV�--��s��؃���`H��Ӱ����,����N���c�m�7�ߗ��
O�-�q�{1z`a��N4d��T>���od��}�2胷����,���O��O��Ra��a�8�t3���_cI]�g��]TJ�j�$��r�2�0��W[��5҃{����CNCm��dƓF�z���X�-��pe2|�(AA�P�*�Tp�xQ&�u����W*4��� ���Y���fU H(���*�t���a;�O-v@%B `@e��0,Ua��������BTڊ�2l.��!&+N��]���R�3���i���0� Z֮9
�ƀ��w��z��m<��7�(��;��y�j�LU�pl���P�q��&�h7��	��"�[�{ad�+R�yv��@%��͌��!�����|��kc�3[N��]9�=��cG�/*��μ9gHa�1=��Z��N��F%���ӄk/Z���a��..Zx���G�೟��o�z�50[����5�:3s��0��?�\����ߠJ2�w,u0܈�<{m0�03����Vi����/����_���>p�u�����aO)��>�uU�ޚ��kr)Ҋ7�rU)�erq��2�n�����L汥θ��f��֪z*�s}PTc��J���G
o��ͿB�^9'�d��&�u:��
͕��P)��oB(�0�����ǵbw��ȏ��2"�����������F�����rLF�<c!�8V>�q���Ͳރ�HY���k{*��k�X�;�-�V�v�=�T��ԣj)Y������qz"�5�,�3��d@�i�������.�w���K-��`�*�~#��v�=j���X#�]��\�8���x0�mT����U��t����	��;�³�`S8�I�3w+�/|4���^_+��J)�'�,��2��-]�2p`�%��A8� �Nqܵ<��ڋ�Q�^k��w�����y�1�;A/���w�p����h�扊K�0�wt��K�V,w���O"RQ��-Z�&�ړ�S�G�-���6Ӻ��H�� ��:o[K�a��qC�;Ȏ>l!S\Z����8���_W{oQ���$3�ِ0M�Kt^��I�k��Xz�8aK@=�ۘm��`����ڊIsEA_����FwT�'Ъ�)3F���u&���a`i����rp�;����,zڭ��a���2r{�P�}�k�cnĊ�c-X��Ie��<m�xm�fX�����+-��4�n��Z��G?��sw���x�|�5��:OG �K�vc�U��MHW�����\��95��`�1##Ke	�݅�~��kୣK�����߆�<��p-�g�{߰f7,Ý��e�T5�V��T��`P2
Nx(FY�y&�6#�*_[x��8H�O�Iy�$�����]+����ϢX��<�~��WW�0(����a�t�IyN��e���a&�h��8�a��m��܈i�w�]!1�l2��8��5��h�6R�9j���9��i�4h7k�iGh'6\���G��q/2-�)��Y�/���,�2�E��b�-�N�eٿ0�1:R��8Ҳ�p%��"��'�~�QU��śf�o�&ɇ",�M����$qv��{�hcHb�!1��ib�īR^B�:�:���Y��#��ݍC���i��9�9�r�)����W�8��t3�1��#�.�r�q3���\�Z8o�68q���Vh$���K�Ϣ�.��� i���KK,ʈ>��������15X�$�K�uB),�|}���bf�,����)QG-p��|�g8�z��S������:�c�;�c��h)]�%�w-�G�ӹ έ�[m𴑒���m.�,
}}�p���N9������5�l�@̄×�d�\��	�A�ɛ���q���o@P�-H��۴���0�5ͮk�Re��&{���J�tȳ�ֈ�&�<U��s@C��&H�Y���� I0�}G
���K$o�M�oL�d�J��mр��g ����ڱ�1������,.���?o�f� ��W�����п-��&�ԗ	6�$�e2O��o�~��8���WjI�1t|����a��&\'8B���{�)��BK�����.�>x�u��;>_�ȇ���ux����>��0���F`�z%��7iڀ8Fx��Ր����a��ح���Vcc	G�'�y����/�z�Mx����}�7�Ӝm����W��6�������\ꉊ�,���x�
�p���<�2S
��~�p9��Rc��vvr�an��ے���O\K<���ַHwdd�G�XM����I2ШS[B�}��Y��EI���y	�C!��<ⷉ&�h�T>�����
>�q�p�m��h�EIg4t-"d��$$4�����{�,�_�Fn��,p/b�o�椩�qa���]RF7��OW�9�l��l���=�#�#�&�i-�C8@)���\���{��k	����v����pV�UqJ�|c����9f��z���a�?�)�OH]&�8�������Y��ɵ3���CP��|jS}�by�I������1���>�9�.A�%��9_�x`fSc8�5�j�7�o���立�x�@��:
�����h-N� ����ky�_Ʉ������8�}/�S�E� ��5�����T
%��Ж�5X%]�q�3�da%�+�����])g]*�~'@�� X���p��x�0DF����B[��\�˼��w��Jc���<p�V����<��zj�3�A ֗cD�T&\t���X(�����9l̳]�]]t��c�x�Hf�3�v���ސ9�	��k�Ic���ct�\o�T���d^�.M"�dGҒ���O'\tPn�Qb7��4��r�4����6~���ֵ���8Z0�U��b���|���|?|�w�g�� �z�;`�XX�ˣU�h�k�aH0	߶��n��q�hg^5���h�kRV�������/��x�A��?�����9_B� ���3#��D���X�L�Lʺt��p2�=���˫!�����}D�YIt��PN�uR�lA���A3X���XC%�G�]���,��M4�nS��:���O��O����|*
�p=�I�3�6Eː���.�Ƀ��4Q��Cyzc%)�O�c&�k��"N�fI��wH8[uYħ~S���䚡��d"��,%_ڃ)��nm�K,��jE�X&��뵥�[xg �6qeS\Ēg2�7F��t��
��A�`�^v�L��(Kq��:P��o����A"�sR��8�M|#;�,�N������w�T��H{���������p�;a�3��4e���d�� cW �S��wC��ȓ�Ė�M���*��(-�e�P_·�3^�}ql�sJ��B9�w��*=��3C9���R�H�)���ps'\��qy(3Dc
�t��:�ٕt*�3p&@Fa��e¬��ڔ0��<�0�����N�<�1
4�DM4Ѧ	� �y]}4NIZ���	�zrp�B�e�E�B$�-�Q,��2 �A���zK�|y���_�z�]����@k�`�,����{�5�۟�~�K_�O��=p�n	��r�.�s�§�hp^68��^X�������K�+��Y�����ƇoW�M�\��Wl.��˗��g���<�s����.�ϡ�v���^{!�ˀ/c�x�\�L�֦��o$����4[<K�����{�I�T�!<�t���]�3�y��g:-�%����yN���Q�@�NM8�DMt�ԡ�:9�SZ��N�,.�5,�NQ�.<pЫ��W�)rs=J�$���H�i�|����6%sC686"}�Xڏ)$ ����!�S�{?�p�hYx.걽�΄;K�#�)e��<��Ɠ�,]�@jqF��g�6K>'QҸӰ�I긗�>M5e��[�~�:u�ܑ��4�r�"\~b'S�^�X�;FW���GM
qB�=F����+TԾ���<��e���K�W8�sw������D��IU(�1��I7f�>L!!]��~�z�ǆG���''Ҳ�J�5�������NW��� �GX��\fa82@`e�w�0h.��h����U�Y8��|�%���cʑ�8ΘR{��$��!_'ɺ��o
gO+Yc��9��Q=Q�:���DM4Q�p��Tk�K��^7�����K�5�l���4�N���%��
��@MGr���"��{��%�ò�H Z<b?��ē�/K]�{���!^sC�꾘a<��wݽ�ݢ�߆k$��A+��h-�usw]�֧����]�?����w��-ay��Sy3���\��=]�{�ȣA���a��kf�k�K�]�⬾7{>�f6��.�=���{~
��x���U��l.\{��o������8�z��il�PO�B5�d jR�}��	�(���6�iYs�Vex�t/�euz�2�w����>��)
�z2)�7;�O(Ʉ��`�@S�q哭Zk �9�+"�A5}�6Hk���:�D�ƌ���V~5��7���R��8y]��j{"I�jq[�S�%�v|p��nˠ����1���AFQ:R:���bRxu � �����,������`�ɕ�`��B}��j��%
r��d�R�����W%Y�$�w��!��܃I��ʥ�YB��{01��@j�5�<./�R'�JW�n�x��CN�h�_��[��pO#=p M�N�4��w.��r��S�ē�Ɲ~[17k[8tEX����M:�]E�A*:d���n!�m�R�=q��G�/7 ���[i�~���/wd|Q��u��'f�T��������#����$��:��x�ʅ|H���@�n���^}֖\S����O]�"�Ӊ�ku��.��0��,%�ڨ'|��4Y���Y~Z�6^�����`�za�Kʷ�ĕ�b�6z?|�n
�ٯxL������z���t*�E$�S�z{��b��q��5S�K!�3����x:4�شq��&�h���đ'[��?q������v�E@F}�^{��S�|�j8f��=v6o6��zRnl�ձ��{X�ϑ/#©��a�rLQ�UJ�mࡂ��5�]M��a���3�rf�pf
�R�
�AA u]���xe
���.*J|ܺ��fWp���m7�������>���]pˍ7�����*��(������a�t;Z�$���J��iC�~6k��$

�����n����˗��^������??{�x���8��u:
�F]J�`� 8��I)�d���m�[�IH�a�f�u�z����T[Iim(�(GW��<�f����i����)��Qi>����.�vJ�N��76H#�3\���׆Ks���WH���?�a�o�F�*�K��5��"����h����q�G�1�Q�8�7�<����(����)�Q��nӃ0��?�$�� < 
��	?�ƚZ����I� � "M��N��T��� _+�5)�@>�L>a���I���܃����&��~X^� %�m;q����-�U
k*�9V|�z�9��x���Q5��@�j7Ĥ������7j/�� �����)eY*.��[�h訕���k�pF�����4�s�LT��d�ǬǛ���U�,�3�|�Fp�X�wBY��NW҉���iv�m�P��M ڈ���.�9$����T��3��� g�~�Z\�{��`U��iM��'��Y������z�ԅe@>cl��{�P!��������u�/�Kt(۲�%�WpR����qB����"}�}ۂ�"~V���-o�Ⓧ���,-��i�Q'	����A�_�]��k��F��~��9�����4���M�e���h��&����ζ%E����g��Ȱ:�]���Jݩ&���Ic����k�f*��>��RR�KPű���Pm��.h�98}��S�!^��7���W��b��7X
F.[o�q�b	�_{��g>��������p��}0�Ucp�2Z��Þ������� LA�EA��5�g�``���x#����|ţY�x��Wỏ=���}/��,0ۻ fo���kV)�ʁmᔏ��$^��`x�Y�$b*�52�l�I����Q���<jRW2@KLj~	���/`��.Ee0II�J�GID��'�)��T�e]C7e�Xg�qd{�t��v\��RГΐ0M4�nӐ�gW��&l�5q�e\��\�p͜?��Mg��*�7��FLږ��L�yi���`V��u����6�� k�U�)en�[ڃ�F�i$]�H8��4�.�)��r�9�u��{�J~�bR�M�9�0�o��g�w\���]��E�Q�h��i�Q<cb�����;w�"�=Qsc��o�q�;��P�O�r�I��9�Saxg �.�D�Jh�ϸ�j0u ~@
��
��晓�(Z��<�, �Ӧ��;���$����~G*s,�Ż��ZL���A�H�VZ(�8t��� ��b1�zB�.@E��0E��3տ!i�j�-EAHO��	���aHms㯡ͯA��	#�+��a����#�΅p! ,r�aJW)��\V���@cR�i�,>�vNe΀.	k�ߕ`X�7�{i1J�+aڛ[��Aa��~����~0��
��a���7"@�ᤴ��eH6�Rx(��;�&�h���E�Q��t�	i�B'!�(��F���2�0L(������#��s�|YZ�f�iH�(FD-Y�HT��h�j#����d��r8�d���1��c�N�_:��!�|��÷�_���w�~�mp�5��ܹ�X\9r�{/7 G���-c9�G�Q,~��_���m_8mjBH2|q�M���*�|�}��}�9����o=�8�쩗��/˃=����g�q�M@Zw�J��a�xq^��c�RD"�G:�;V)��ްfB���dq0��[�KE)yM
�z�GK�L��޴���L��2�q�~�%�8�
�6�8}p=��w��"�w�f�jz��&�u�s�5چއ�����Ҿ����u�A�6���5;at�ў�%�J�5ހδ���m�S��(�8�I�o�鯓��G��r�(L��}T�OqN��6iX�{0��n�z}����*��@��ej#��{B,�g}�P�H�Ԫ���hۂՇ0�0<��1���;�i&߰�4�pNJ]��hQ��;G�t!ˋ^8x��8V�#a�T:�@"C�\�����x\���,���[w[�%���_�(|%��`:KT���?ϯ4��"�҈��T��a�, ����8�Ҏ�Y�'v�Z}f�8�N�Zx�N�E��:m|�6g��.VYSmԼ����kz����>y:W�ĕ�yC�A�p � �+EF��bL\�I����3ύO)C657�r��((xey횇�P������,�l�`m�F�4�����rUo!1��7,?k�9��A�hv�B٥��h�uD��&���Qm
;?�;�Y:ӏ�mwt�
���I`���1�叱�me�t����6p����r4�,Z�mM�E!H%��D,k��F�DInj�o�=��N/��;Z�v����n�ۃ���^��>y������7��ܴ�S�a��g�|�;����#�M�mP��Y,+
A0�W�4Mr���˗��_��=�(���g�O?Ͼ~	���Fsp��=�Ug���lc�w�w�����%��f:5�(_��x�.Y��T`͂�Y*}���.u]4�Ƭ�b�[����ch��ׇk>���N��M�Z�Q����w=��q�POS��7J=��4�{8�����k�5�DM4�z:(~=E��F7O����yh,C�	.Nb_��!�m�T��F䡖��w��O7P�X)��R�i&��蓙���{d���J��o��,��g��
�����W��.Ul�݀=�.��\����԰p5���?�/6�JB�u��/(1�h
��$�x`�|M��ڞ�_p����J�	�$ir�II{��̬���gvmgWI���3��_��O�;NI���6�ݞ�5i+���F������J>��`}S��Pb\�.�/�=[d�
_�"Y�Z���a�]��@�2K�mm#o��LՇңb��ӊ�!@�$d��xY+saҧ4����͝-���q�>ͅ[ ��P"��C�Ph���c���'!ptQi��I��F�;��Zz�uO$(���i7�<p`K8�|k�U)���TtּIx�8�b�9"1��
�h���Cǐ� �+qz�Ge���S�݉k��/���5�")�y���x�ʢmQX�w�W��T���mU�<�0~-LD@�8u1��5���@;딵b���P�C6`#�F�-f��a��[0�XBsh�A���¬]���y|������9���o���{ �G ����
�ux�*�Ҡ�@Ąm��x5�cƲ��0c\��yi����yw��Rf{0�x{��^}�y�1��< ?}�Ex�=�K�0�.\s�r:�����fLf�&eՎ�JF��B"HXO�b*?�����3m�XT�&aXʻ���Pr�w*���$f���yP=�� d= �v�؁i�g�d�:nȡV4I�N'͙$���G`�Q�H�c��'wjk��{;��Xi�>C�:�w��J��WӉ&:?t���f�:�s.���:�� p�#�5,ঀ�~뿘x��X/�\���u�I�ݔ.�K�{WN�C��2�@�f�Ơ�fN�h��ܰ��,��j��ڲw�2X��M�WWI��r�*��6[�eQ����j)�n)^-��$at �p]JG�f�� ��ZNgV��q�|$�FŧL�8�N��+ %����C�aouX��m�)���7N���>�i��}���pl�̑s��@�2*G�p>��i����Y�m�%i��
�����>�u-9�pRO�x\�=k�d(%�H0]��3�n�u '0P(�w�ł˕����b�`�U�� }�����vENzy�j��?�&�)����?jE�V�����q��S�c�������������E?C:��� �(0sE���0�T	C%���Z�L8�-&��({F ��~���b��X�X|	@�Ǽ0�*�����h��N��L����٤��b@�87���F��+��,��*�5�\]hw�%�X�94��9<�*b�5�O��H14�o�-+�?ml�����-s��}�iU3�"��=awÐ�E0�°��4x%
^�´Q�B'�D_������\�/���,��3���s���?_����[n�k.9�]��� �G��ڥO�]L��E}��p�8*�8?^�`�1kf�7,�|��./[x����'O<}�O��=����h/ ,`������`ng1͐O��hуG��� ��ٸLo�;`F�]�����D�%)���m�X�Ry�l�d�7]�P³��_���G.�r�=u�2=�������z^�D#۲�P�6�fD�_Z�e�|���k��:v����a���7�֢�6a{���˪pzԵv�n����!����&�h��P�Mq)ǋ��/=�0\q����,�5�B���mY7_7B��yY����r � �ʔ���F\�8	,Q�-%�%���O Z��Tu	��Ƣ_ě-7'�&y@#m�Ǫ�g�����E?�؃I�K��(��0�#릾��%>���	��L�(<�񺰆Q�^�\°��4؄B�pqB�l?N�н���`0L�#`�E��g�a�wK��.�����>�Τ�8��Պ'9՗茭��Sg��8�\��'�	"�@J���r$�8��j�U�DpH��jAuTj�܌�f��x��Uq�����o�ⲒT6��,1�r���`
���-O�Z?�l�@�o(��i���(�b�������7d�� ��X�M�P�L�~a+�y���EB�$��������`:>jl`�,M�����=�|uS������<�� % ������97�iqS� S���G�
|~*)�5@�s�z}~��M4����ꌑFI�zW�e�.�(n���q�&��I��cE$k�h����G��;D}�h�P���CNjڢ2*��b~���^��"�(�I΀åޭdҥ�����¥Ko���3��;o�|�'���|�]��Ź��n~�{ō��o���<��4�o�3�� o$Qnk���D���CBY���}�|��.�/�~�s��pϓO�O^x���U����*쁗�f���=�٬����܈��� ������P���. e�4��՞���@^���\�{�W�D�9�Q����~�� ��(�'%�U�!���x|Wh���NZ�=y,�?s}�]2:*�y�-���(۪��lT��V����.�̉&���)��g��Y��1b�6�\�I#x��<[����fjӐ����W㫹 l�K��^���^w!�i��S��T�;$��t��i��^Z�'�x��l���r/���zl9^��^ђBz��� ���T��R����g����-h~/cZ�\6��m�2:��H̀�`09u(�*��YƜe-R.W?�c����;F�ח���'�g���n5�\��L�N�X1�X��4��������5�7�?�8��IY�Ǥ4R�1>�Z���QG��1q��)0���B��V.`��x��)�tEKȒ�F�T��е�4���VV+��V�J����:/z�y��&���Q�0�R�s��D]�#p���Φx&�˳f���;`�ªZ�*f��tT��,Ↄ���`��3D/�=��$�y2m@��N"��M�l�)��Znn�O�P�8祧:(Ί������L4�D�I�1��{*�IK�0t98w�<�&���9{��������:kdѶ�@\�Pm��&	�^���4�-�Do�?g�aQ����h+�t�������=7����K�����z�p��kB�+�dWB�ή¥��L�th��������QX�*e��if��]�bѸ�ú��./���[o��z��ޟ��ϿϿ}�\����̺�>��m���7�����SwLNjD'nܡg�[��%��E�b[�����"�B��J��P9Q��쥒�ᢕ՜�6΃��Q��E8\XC�G����U��I�aU���d�Z��zT�B��פ�q�$��]����ޟ��7�Dg�N{c>�'yV�����#o�<c���	����Xlp�ٞ��U6� ��LO:�����$�P�S8�}�>��, ������M�3BVA�p�����|�Ǫ�l?�������Z��O$���4t�`X-��d��R�4�|Xb��t^-��c��/x}���8���	c&�y����xHaO���t��F$V���[׀u#�&��Y0��.��7������/>G"�D7&O����,�P��������|O���o�d��7�TТ5R��p��t��rCk��$7����2������^��TN�����e��J�&+�X��)Y_�)��M(�4�(�E�>��[���!׍���^$�kR�Jň�L�i)�!��i����V��X����8_��'���=!v�/,H@صnv��)�L;�%�5K3�c�d 8&:�T�7!��=ߌs_��Ru�� �>Gs/�V_�bjLM
�����HX^�s8k���ݺ;�@_�U�Z!�)�2Pl���Q~�ЖDX�`�< �����ֲ�G�����>�w¿�ڗ᫟�$�|�E��{JV�=-��ШJ�&8G�(H�#�J~Tй�6�6MHǧ��N9�z>s���^y�m��S��������s�.��`�g0;8�=�K���W���ޡG��?�͆$�`-z����ʍ�`$\��x��d�Jf�r�4�,i�rZ���^��j�Í���W�s�9yX@�	�\(t�Jk����C)ζ�4�j��D#f�rd����Ξ�h_Yò�)��%�v�������~[xl��&Z�vmN
^���S�g�4���H�A��f���S%�>'Z���S�Z5�=m�ނ\�:ƈ���܃!U��Ԧ�z�o����z�;�m����!w*�.�ʍ2/�
�{���]ɖC7��ߵP]��gn]!���$,�O��Ȗ����ߥr�v��m6S�g#�E����iI~J��%@�n~̨O�(�?��i�Lt�������Cl��N�����gC��p"��hȀ�d!޶OY�{��ť�m�L�$���-���'��E3���H��)��-*�*���\��{-y뵸X8%e��^��e&*�P���5��9,_ڢD@o��)DCl!�5��Uk~�=��Hj���D��iQ��و'�!�.ې�����N�	��d�k�IY���s�څ�GX�NM�p7p�'��O
�ϒ���M�͒��/ �T��9զƆ����zF��z9D>d�
�wv��Nʹ ����(�[�����[�ޝ(�1��O
��g��$Y��rǶ�}i��&�:�|6��:�=��w��	�#;����Y#a�I�9�7lB7m�:W��2�e��X�= ��Smۈ������y����f�ļ�T�'�a�M���KJU/:M�7;���/c1�1dR��+r

��a1��V�'q0�m� �s�B?��vd�+Gp����}���/�����w���C����aȠE���L��"�$y�!,�E~�8��M N��ƶ�����s��^x��G��<�(���s��ކ7W|�V���"7=e�ʶ�@3g�ѶF��5T����_�ɕ�k��+�[�i�A�l|C!��L���M�Uv����k6W&�{ò��Uʳ�^��!���5u�Q��'_�J��g��pܹ!���ޢ+n$6:W�0�?E:k֓���� G��=~؆MޯH.�nVXSPn�H�L(����}�C��wa������Tz}�&�h��#��77����zQ7Y
#�%�U%�,�3xU��C�Dp��ƐB)@��F�¤N�h7i(����)�����P��tS+�NJ,��Q����:���'�jC2��g�x�D�@*S�d�hd�6����xf̎�|�!�����N	�:M<_���B�_C�,��&�LX`�)�atx��ܥ��楜K�y.��-��di3���2���Q�=�á;ԩ� ����=�R>�ֺ���8%�)����a�T3�mO�L��a33�]�����+���,�E:[�i*YY��y$��M#�b�Ɣ�o�lT��N�X�u#;���+.�&�bh��R����.n��KkQ/�O�9���o�t��;�٩q�w�0���<A�4qb�?0�%TR��v�b�K���}�]J#-F}-�'�R�A���62&)���7t2|!gP�WQ�b.�7H�p\����p��?�<�����k��wumV�tNӈCuE�,�{O��4D���@r��{�(Xp>���l�6$�s�]��$hq���g���&�h��6@�[c�o�����O�5ފO+���C*Mz"Z�Z�W�j2z�8STS`$8o4M����N�!;��I�%�bjL��p�p�M
[��Lbum�ļ��z�>�bT����L��gf+�F��o}�.��_�m��m����3���u$ �6Z���F��F=~�ʱF֑i#$Ŕ�2�ac2�@H�<^Yx��g�?����gϿo���up�+�h��RT���+c̿�`��*�u�v{���$L��`#��Y6-��E��mg��y +��r�'>�B�?$��da ��|&
[Ёh�{��N�8d�&.���65�����y�b�(�i��=����-��,#�<�S���RORM4�NҮr�߸F��&,�z�6l���D��	��y�<�X�k"���	F���]���̱�וՏ��,ۦZD9!��S�<�G-��PUf!}g���DBk"<�`!�a.�>���]no�ظm�!f>�&��ud�*����b�{�F<j�%H���K�V���[��S	!�َ�1�e��D�9/��Q{0<n��y��6���G!�nȕ��Θ񍐇��m��,�t=�����"����}�m�dD4��澍�n F��mT�梬��� �[�7~/��70�Fp�$Ud�(�~��.^M$N���#����m�h���!V���)�*���_M!�͌(@xo��>��J��iaqx��;پ���
̏����xv���&-C=��o�����lq��RN/u�.��
E��H��Nb.-��fo�o�^���p���o���?Ǿ"k��)��FY�en�ӑ���wZ@�+� �o�R2pi�����e�4ᤛ7�����|9S��GZ6�G���DMt5�x�HcQ"[h�0����0s:I]�9^�N�tѶ0�P��O��ߵ!�0 z����������(\A��r�d\l�rt	GW�`����������n9� pti���_Ҷ4.�t�$��[�(��p��yy�M�2��4���Ǹ���6���_������C�̢��� {�z�9̽����Y�_{`\�M�60sX�$e�W�2e!W����f�mY�HP0(���ⲋ�[�@֖"�F�H���@9ɤ@�}�m�{~-y���3c��V�R�"/�e�a� ����#�ӣ�|m��_v�1ĒB�r��9��	�DM4��C���&-�~�D��6�4���ѓ׈�,����߀[�B\���WfW��] �ث�Cc��=>�3��,������ڈ�2ܚ��`b$����xͣs�.��-a�z����J���k웕4А!����7u�C���g���ʕ̆�c�� Y}��݃���]�*��9�VKvI[��ﵒ�=��Vu�C�$/v���H �l����(��ȱl���rW�7qφ9O�E�~1�6�H�B��2�0�g��w����LZ��;hŊ�S���zT�j2|�(�Ry�Az��c[�( ��,��tnr2�֙�]v������y޽|��fp���jtZx��ex���b�{p G��8�FJę�E㍰����a���-R�r��h�3��5�cBv\����ҵl��'o<�������Q�P(Q|��K���p��R�J�e�_:M��P9�\�)՚��z�H�,9�E���!��	�|EJ�s�7f�@�U��f���N��(x�n��i#���.&�h��N��ǝ㑢�76��Z�n�ܵp+��uk�S��I,�1
�c�t��7��4�M}��E�t����7��B�i��໬�����
>�g�y���W��U������Z�Y�����mA�:����4��^��r��j�G��*�٬I����N������X�Q/�����_�7�~��S����+���>̯Y�u.	�����LӬ��뎚��@�y�:m�	�_���.�Ǵ��51���:*�y�sZI&����W�yŷR.v�>C��Ĭ@���A(�Y���
�'e�=pp�+��p>�1���u�4}���Z�
Gy0�oQ1�Y�'�h����:�R�8���kD�v��z�xh	���'��q��e�����[rO�J�x�#a`��)v%�C�-�U�C��
@*�A�~���(������U��%�V�ޱ7�k�`�X��.��C��=h������@�7֘�C�ޔ)r�[�aZ`y68N�[)9��lІ�E��ǈC�)�)5ra&q�����FY�%I�<O/��#��,�c[�ec|��1����x��1d��0�3��փ�9�齜]ԅx�#��8���]����PAJJ�_1��UJz#V�Pʈ).���lr3��JI>ykWE�[Sk��
@��=N���"����e	��D��.�2*��#���������_����n�ۿ ���K��#������G��V���xp�*���U��z��88����8���� S��:���Z�P��
�R�����U�ݿ�o���%4@ ��\	��H���Ft���އ#��(�W�C�:LÿQ��Ɨ"	3�5���i����6��R��X�	�d &.z���l�RKm~�^��Y��G�@b�$��.U��g��0�"b+QZ������R���þ�&��ꢒ� ���������]�������"���&�^�w>��`-b��0D2���}2bsDJ�AYXR�8�㋯Q:�z�F�����g^�K�H�u-�tcJiH7~mR����涁��z����p�l%�,��X4� ��X���ZT����M2"��cQ�g|�ʶ��|~�q��{��<�<��pi�v�N�^);wqZO]��WLC�o�w�*xOy
������F^�?e���F	���COLi���T�>�2X��
��6	'�pi�lg�F�K1ۜ�[�<X�X�)���x���lZ��_Ί1����j��^FY�{���F&���Sz�7�;��Ұ�"����+re�<�HXM4�D�J]�����a먇a�Y�y��V|��P�M�¿��IKF�#
�ɋigcm=QB�?�����%t�F9{5��>�}]|�rp�84N�&l ��:j=6i���raGW.�����>�Y�g_�n{��+��O=�|��G�?��>����å٪/_8��U�C��b���*��
N&i��]�05�EN�i�A\��<"~�oT��ZU���7u��Od�z�yz��°�����[!u�'#�
��`Rw�R*;�J0v�?�T����)9i��l����4���(~j�V��\G:��m	������.KZ�h��<I�����.Q�Ŭ�'��j��j+ޡ�C�j��畾%��r#+�)�3L���f�+�tP	rF���ؽX6p�p	w�����{�ُ| ��x pb�������~��_��?�|��o~����g�W����+0�2c�|���{���@i�+;�ƨ�R��6X�Rq%��K6=��qUŶЏ_�Rץl�y��T���N��sP#��S��,ۤ:
�\�3��y|�����S�?,1MHN�Ӊ4�F�1�S�@��f��١���R���r�>7��yҐI�l����-j��H�_�l���e-�'��o?q�9`��&�y*mz�6zC��u�1\C�,r��3��m�^tb����2Ga��di�j)�z�5�p��m�j��)�'ymJ�L��Q6$�(tqV����؍�U'^�:{�����[n���}�"��()%+Qb�h4x}	^���ך6~#b�.���[�⫯�=�=
���<o�p���̍�C���oaiRk���P��LFv!87	���Z2�e�	����KVe�P+Y��2Z��~S�\���W]p,��s�c��H'�Þ�a?�ѷ>lC�ѥ;�8���� z�ө0�2���P m��h&&�h��N�J_�y�=�Ç���pۈ���^����s�7���hɛ\�*�Uf�w@��Nsp�q��>�!+�i�F�w�  C�?u�O>�� �m{1+���p�!��?z7����
���wþ�[9
y����������_��|�������Sx��aq�4��>x��#��Һ͗E���j�x�J`j���c�1���5
�k60�u�?�ڊ�䥄�'g���*�f{HVJʀ��T��<$Br��!C�=d�sXZLD���X.ۤ�'�pR�=ǆ|���︨|�Io�t �|YM��ra�Ʒk�6�o`�m�u#������!TgP��NtRϨg��'�K��z.����/���F,[j��K_��6(j�شQ��7oc��n�^q�����_���x7��0�JCEj� A7�f���>��;����
H<�8��O�o��1x�����w��1_��*l�\�	��{0s
I�D����/�qC��T���%�jCTi	�!���Nҙ ϰ�e<s�\��̩F8�a�"����߉�,Ѐ3l�l���i�/*��4�Ϭ:�zMr�(-��;ĉrZ�E~�����[z&�KO@P��<s ��ʧ.t�M���0�DM�-*�O�v���� E�I�nV��i��@��=���]z�ܓ���-`f�u�񼨋L
S�68\,`�`��-e����3�@��s^cFQ�x���x��ߏ�� �r���<�������?p<��!��\�9߇��|�/^}�z�<k�X�y�ʄ��XG�5r��X=aa}�t`P��A�K8-�/$lk���	�I�(�TZ==�6��yTu�\�����BTF�B�̤�ڈx�*��I�4�-,��7�m��7H|��Ik|z�Du��c��:g�<�DMD�T%2c�:O�,���Yz��a����W��rY�Ý(?l�-����|,�f�`��$���B�ۅ�>E̺Q�_E�=�s�]���K�'��������-��,����o�{����k/��>�1�Gw�/����'�>
���½Ͻ�_Y�[G�pe��'�f0��O/0̜7?g��o���mA)��1g����T}�������xhUa�;QfL&[_�S��ڡ>��`x_�<0�t��{� è�,7,bY�΋-+�vӓO�,>������]��.����lؤqr.g��&�]�b������٧l�/�T��v��[:i)R�A�:<� BL 'i��~Є�w#$�R��D����~oW����������w�gA�i4� �6�Tk�pÅ�7��,|��O��}�mx�g�/��!�͏~y	�2+ q�����u���j�xiӝ��D;=o�g,��E��$H�6�&-�Vs$�R�g+h)��bf����tR��Lr��-Au��.Ig���WE�I=�(`m�z���Ϲ\�2*��:y��R ؞*�0�U�k5�a�%����DM4��Dݘ9�v#h�c�I��.\	��).���KIU�=+D�={'�Q��P�KБ&eU˴+ޠ|��k����.�-7�u��q����D�q��F�t'� O��|��������g�������0wW��m�7si��M]H62�x#\���n\�B�U�'*�4�{%,�}�l�oZ�����d�*sRQ���PV����=뾹��ĝ,L���3���<m��`�"n�Cz�$4SM4�DWu�a�e���֐�X(����+��v�`kk1z��H��7�zN#�3��͘U8ai���`�2�w�#�w�����{���^z����[n�?�W�\��G��(W���nfY��,�����m����K�Ͻ�����?|���G���x.�����{�}a��5{~��L�!�d�`�0-�?B�q#k�^놿1�"�N���M�Sy�u�Ɂ�Ե�q�+&y���J.���WJ�wf_X�Y?���v�p!{�f��8��$wE�����76��pi��f�>	Zπä
K��w��k"N��SYE�-�P�>\(�b�<�b�������xAR�)v�_�cQo��;n�&��tE
�7i)]l�e���Ղ~ǻn�������v�>hv�+��
���`�x7·\s��;�K�4���G�ؓO�w����#�^�Ë��b��s�hé6�d�䬙���]��Ѐ��`*JbؒZ�T��}'m&�~R�6��Zq	�O�򕚧HFD�F��h��尤&�~����[Ʀ4�2 �-�m����}m9�NcN���&�IZ�0��%�Tc�X~�T��/��?�1�����B�_�B}	��U��L/���1�:&�����&�h�ǴZ�O$^�ۓ�����28�b+��^���r���M�V�:ʌ˾X&G�T�V���׫�7�D�	6����ַ��n^�ΓŬ�G^~�{��گ��
�^�Iv ����d̕����o��/� ?z�q��S���O?ϼq�l̮��������y$t�$s�q���c^M���m�CM���#�����<��ʄ�jKv�9��X��wH)�3�ge��������`VřZ��G���r�|��ޢ4_mw>�����bxsf;�eB�E-�!-���+uxb2�y�CJe8��ijóA�yU_�����[�b���B^/�Հo�ñ%��a���춛����}Nl�B�I�*�қ�)Sһ��\U����צnȘ�:V�����l)�3�hl_�؝p�;n8Z�+�`�����Q�����,���t#���O�?�§�W_�y�}���͇�^�G{��r��r�ȃ�݃w�X#x-d���6���[�Wi1㋾����<J�$�āZJ��o<.;1��*n��so�)��d���C��� i�MYf(��~���%_cE�M�zv�� �=������з��('׷�7ןf��2ా� ��J��S���͈G�Ŗ7N��O�2�7ZZ���0�6�
c�>	���?!h�0�3lp�Z�W^Š�w�4:"�8�g�#��;C%�I���.¾��"p`��"ZRL��m-C��
���]�|����y���㿀�<�(���'ᑗ_�׎�`��`oc��5z�p����7|ç��ᕦ\~!�2M��4 ��W*��@��V6r��gL�W�cL�o���'����?�&��~(k��<-��T�N�HկU_F�4�j`�����B�%�r׎�Ȥ�M�t���X�q�M�e�]]S��z�����O@0zCB�as$����ҴP64ް���*��� ��:B�H�KcF�ش'�h����cz{�������~j!��˄}�d�*�8�6�������f<��&�� "8�![L�,Z�D�B�i���QI6�Z�,~Z���S����R�0h��؃�Q8b�1<���5ޫ�ˬض}|ޢqIԏ&��3�痰\�)�^���_�%�}��p��A�k�v�I�;,^����^<yc�W^����������>'�� �^�pp�5�4�����y�VI5�0]�Wh���%���і*�6ϥ����j������d�Kʯ�־�.bU�T�?C*�m.w��{+�0`i��9X��6���P=��)t�=����Yp�ަ]��Y��F�㸑&ƴ��r�$c
�����P?W�>���ᇲIr�������J�קs-���h�d�<�u�� ��x��&:�����6��d����m���ܚ����z`	C��
���k�1D����D+>R)��ڳ��;��؂لK��A=���J��%C،~��2�kuJ��pg*�,�n�ʇ{)�}Z�C��M�n�f�����<��JX��a���1a�]�����n�ۿ�%��/~�x�e������~~�����.��\���0�u��{0Ψ�b~!}���]�^� ���e
�JZ�+S���-\��B�F@2O����QNȍ7�k�$76��C�x�����\V�窑���~��ץC�}��P�@iox�Hl]�p���CY�qX�
8��bs��'���d��Ko���b">�0�h�PM|K�}��;��;�
�^�Flβ��iY�gʓ�I�軜���zAA�U!RʸP"�1�;�'�`�h��$P�K^�%�~�m�|��k�*��8*ԡW�E�e��l�/l��ު���n�����������!�����߽�q����.å�ػp���X���D���6��g�逋���x���;��-��cBT�5=ƅ^5�j�B%��V��_�� ���v%��.�gE$��Ј)"(+���7CI�;��ҟ�]j�c
��M�]!p�g/Y��73��Ҁ\���:����6J��-ژ�D�a_4�r.���R�-q�h
�P�ȑ��R�ň�{%��Sbm��b��&��Ձ)�>����9���C��k,?��@�8 �zV�?%�Pz�Gu���'�w�E2ۖ��
�Ȳ���T.�N�]zܖ.}�v�œ�t�9_�H~(��a:��2��� ���ƣ�kѷl}e�:J�ܠ�j)O�;��̍?�{����������կ�5���bf��xܬ����fZ��Wކ'_~��i����=�=/^��|%��z=\��V��p��J�q
�Y�������		z��'���੻J�]��.��k�նPiB坭��ڦ6���a� �dò@y/�71^�@���4�F��A։<�MUR����	P���e�ӗ}dG���]���5uLCMUX�i��jfrG�K~�ٗ�=]D^0�qEmN�c���9��F>2Kc`�DǑiF`���gjm�m2���'
d�r�L_\�6)3m+�R^�2_
��h����E%Y'�b@m���wlO��TQ!lq=�����x�3��צ4�5b���E�������01�^Li��u� ��k���x\�Y�+�s&���&�������`}t�Ƽ$pρ�7!@F���szХ]�//�< zjc�+`'�=dԊ0��㕐n���|7|���_�W�\�o?�0��w��]�//��h�"�����E4~#����;��u�89��}��;ph�uF�����Z�|jX�r!زz�N)�0#��txC<ZJ���$�/�@%C��'����I��k|�H0aㄗ��Xub����K"�VC�"�<0d���Z3,��=��dq����qQ:#�*'͗��t�O�`�ާ۔��ĵ5|�5�P/Ĝ�!��Tɻ��&�[���E��5��9_��ƣ���S���	��isT����}$��Z���`��_�� ���_�'^zn��� "�����[4i��R0 ��" k�֕#o�q�|_���7n?����z�Y���������+o��f˙���}�ɣu�9f{���
���S�A0m=
�	WM�L�>R�$���;���"��=R"��U���*S�ePD�Y�0<J��!ݓp�I)3X̢�x���pv�Q�a�a�P��s޻(���P�@հ�|!dD ��1��ge�]N�t�/t,�94/p�F�p��2U�b/"�M+s��g���yn;�u��n?�rǚ�i��4��s�4��^��5~��gc�M�C{���H��Xİ~}2i]?.%�h�r�l��牸�	O��?ٳ��K����Ȟ�/�(>[�1R D���-�̔��X����r���ڟ����o�u�����k�M�/��t��x�������#?����,�ʬd��ഷ��¾w�q ��qЩ�3���6bZ���\,;��	KE)���aЀtY=�b�Y]$g>��*��JDN����r~���+®�%:1��f�ۨޙ%����6 ���B��m]2��8Bh�Š�[��xG�
|����A�
ASIc6��JE���8�R�K��lBJ���0�tx~�w��U��f����&��:��q�Pbqg�Ǧa�ԅ����Z�R���A(�c�q"Ɇ�ĥ�*�84hV9�����S7]�m����XpY�Iē�i�6�ح7�]�`���K�3�r�{��J�x�J��C��EQ�ΒFC���&&�@����S��2_�������>	x����˗��>��'����}�2,�3�{�d�o���4+y�60�W�8��-|(�XĆ�W�`(���O�f����8��!@z	L�`�$�<*�q�G�wlq�����` 誔�G<%M,�q�:.�U-L�P�
�עqGv��c�`_��������#�}|��tG�S���������Y�L/c�:���� ����k�T~�C�Iר9Ee��9e�k����z|�������YI �[H��j����?3]�]�۟ᦃ���0|�w�|~��S����=�<���pio��k������}k�����r�QC���+�;0��H��Z����f��T�j PzG�5���&#XCH/u [O����QV<�~�}�U-����֟4�&�ք�~cU�L �w U?�z�m�yV(s1�u5V�B��D�<����5XH����	��7�PI�I���؉�HZ�/��#�9Y�Y���o��,��, ����+�Dg�6���ğ�����<�g��C~H�]���>��8(p}�Y��b���aഴ�q>�����~���]��(BT7&lg:G�J�bB}\�Uۨ0�";k�I%�����P�����<�8���O�������p�;o����E��_�?��^��Ͽ�6\��_�J4rr���功p�#�Eg��n@�Ѝ�㈯%	�nL~m$��)QU�z���H)v_k��ęԘ�|ޥ�OM7|���^OҔc!��Vc�(�i���Q���&�;;�l�s+�;�b6E��0���b1����$�v̑�냏��J!���$��i��.=k�8i�4*l�i]�d��� X�'5�:�ɴt�gc,�u��i>�l��%_o�o��w�Y˼�*<o6/vR�L��׾�I�W:�-r�V���kL����}ܸ=&����v�H��좼���o���e�U*��F9d8� ���y�XI�2��5��s��=?~��X".hºh[�HB�p�� 6^Ao ݿ������9�[/�}��;��4<���������!���V�_��5�\�vnc���S���5�Q�'�k�X�zy�!~� �����k,4����d�diR��@��N}RI�@��.K\(�`��;O݀|�灃~g�V��!������CJ��Dg��0��i[M����f?vkq�6����2j֯��a�ؕRj4pH�@.��Sh�S�� B˄���#,�K������l1o��~���g�O�} �K�"��R���4��d{Q���Bm�_9;Ӌ+<p��7�����󟁗^y~��c�?�)|牧ṣ�����Y{�?ݮ@Ĭ�W��NØ6X��EC��Λ �E�OV�0��+ �(6�9�Va��`���������"XZ�0a��*�A� y0�l��9�Dl�"{1`r>��*1��z֥H;��8B�0tmIP�3���Oa�2ٗb�� A���ޛ�u]gb�>��7  $� �	��$j EQ�-�'9��ݶ�ʮ�+����JURɟ�Kw��*���v�]���v$Wڃ$��LQ�� RA� ��sv���k��޻��=�.�x���Ϟ�Z�Z{�kE�P4�T��C/��-=��"U6}��H �J����Zr�����6B1X��X�۟,L0�Ii3̏��cF���w�I:i��S=#onEۤsD�:�CH�n�����x8�"C��ܡ���q�3�g�$�:�'3�Yn�>�u��j��U��0r�ghi�LF�)OjJ�=����O�NP���6�Y��`��J���F�8�8�o=�8�z���kO���*�`�@�}[L�f<d0\Y6�p�(���'֊"86�>,���ZKz���}!��\�J�}�H�|�=��ſ��>s������1Lb��Q�b�o2�*Ɲ�.���v�!��,NO1��B���SKG�rG��3�1�h�"��� �~�5@� GϐMɟ�8�ߴ�s�������9>���e[z�q�ܮY�4�P��>f%�&���S��+��Y�B
�<��i�trTm�L�D�hHo�~^�:�e���)4E��� �OF��٨����<���V1�I���'�92��i������y�A,1��8hW��{�������(O�P-���u��;'O�w�܏�,4
a}�J�8���0�
��+�Q������5�헸f�n\s�"|���c�����z�'��%�c����%\d��s�CQ��<�õ�yL�v5����9#j�J�M�%�"�����[�D�I��c(1��/�H�U#7��V��_"u���{0J��zUzX��] �����7����6dD�M�V���G>�MM�� �	��'��'�W}Ö���4:H�,�(���_��4�M�J,2�*)_�K��Kے�4����ޠ/|t���w����ࢭ���5(�X0p6���DJ8M���2�'��Fio0^՛Bn��?иh�.\t�����p����O_�w|Ğ�;�\���sQ4���+�ʕ�3&��mL�|}W8�s��
�����0�ыR;�:?��FF �=�r�h�X ������ٌ��;dU�JD�i@]n��h� ��+�~ �5OA:����B|A��N���L���"]�� ܱ@V�Ta�m�5���^�4��nv��r��R��=󃷰�_����.3�����Zw&'�U�Z�4΋zu����3��%-��8�[kz�x\0�5&)ch�7�� �+����^���y�u��R��Ij��Ew]A�I�H'�3(���L1j�4wꍮA��$ק��D��<�����������H֍Ҧ�k!�=�_���-�/��8�3ߦ�;g+>hT��;�n�l,}}��z��it���%�z��Su��N��:�k��v֠n�`G�8�mrz ��(W�x*(r���O�D*�"�1֣�yC�gQ��sSk;�rp�(��^I�aT�k�p�Ϲ�q�˂�Ǒ�(���i��He�C�|�Q��fdW��K�(���!��g��c�?/���0��g,u���W�2����~N˙/q�T�;�n ݅U�o�3kӒ����d�fc<5�^Sk!c�干A��)}��&�k��q=��̵�L�Utep��" C�m�4Rg:�i�F�0��?6�aL˨��>?O�9�Bd	���*ɇ������]�=墘�~������O���_�����c�\8U�z���
�56o_'���QU(��}(�`�j,6/]�g?.߻_������o�GO=����a<���xwP�����A��3���E��4�Q�jҸ�irn���,hk�ǔ��P&@<77���k�
UH+��~TZ��!����ˈ'����^�{�%+袨��Y�h&B����߰�h{~�?�%q$�Mik�|Y�R;E��xuhW��j�+��jhh>�^A�q:{h-��^EǞ:[������l���C܊�ТIo�m��|*����=a�
J����5�>ye!poَ��z���C�Νw��O߀��fi �MD�#dL Q�n��	�f�q}�1���
�~��/9o��w=~�k����④�⁧��Ͼ�WN�²	���Y�xZ-ۓp���D����ᾔ����/�v�N�.?SM"�k��s��e�"�)�
��H��8C�f����a(�4-�R8��\LM�U�x/���qi�dxQ���$���b���b�\	�(�u���d�]	�P�n��ih��|��Z�/aX1%?�yخ�f~��Q�I�,��bm��x{�"���F�$D@x�����I̳�N��!ePS[�k�,� d�A�*2�����Fy�\�p�.��d�7/Ĵ�	��4�8�|���CF属m�sgD� $��$�m����Y���E@i�!�
�8�$ÌCmt ��Q;���Y�t���5)�s�.m�`�X�~�r�I_g�����t��L�� q}����%{�c8	�S@$�(*P��25���T��:�V�5�P�T"�K�o�|"9pk(8v0N�~�2A���C.G'�i�BпyI���S�^�d\���nY���X%
cuWff}�-G�q�F��sХe~I���_�1�f�:0�$�mF��T�gC���{�L� ���\3�9|jқ�l��N>yZ:f�_HF��lL)u8�P:�8L��d��d�s��(Z�s�==����*�V\�%-��a8�h�*���5���Ŀ��Q�x�C����]vz˅� f�9j�w��U��fJ#)�$�Lu��c���lKW�݃�{v�?��3x�cx詣���x��c8���z~�ї�:���E9��#�s�R��f;0ES/Smͷ����mG��e����ރ! 5�%�	�ςh�h�n�`��D��$�]*qҦ���'n���)6�u+t��"�gp�oT�3��4��2�c`ŭ�f�`��L����@Wi�X������Ï�oD�����Yb�3:F����bPk�\(p����?�w��}���7]}��ͣ�M�j �F��h�s�����<�"�P��^7���;q�G��ڙD�=�`7_����[��;��ǟĽG��#/Û� �8]��7�C���@4u��؂�iyCg�}��4)�[�R�["Y�n����59�b�R/Mi��x�e�_@։�hۦ��� �5H��*wg���-�PnR4�V��Z-�#��`����h��?�W��൫ �RRﶥ�QW:庼�g4��}�u�|��������LU���,7_��	��@���τ0��
�)[���z�1�#a���P����P��f���n���L�:���F��� .bMIF06���V�s��Sm�������(���<Mf��'Cka�zDj��G��t���#d����%|�b����>"^p0`�t��띒W���R�f��|���B�+�P'�����#�t��:�0~��Bn�\�~����|ZLI�߄k��2ż,��2�i�*��P��"G!��5�U7d˙�*3�ь'�5�9��Z��������a���򦻂��v/�k��0c�M|��ӊ88m"�O��+!����Dm_C7����Q�;<[{�_�H���r��|� |��gp��g�k�����w��>,g3W+��;@k�����������#
������԰cԣ�y�|�e����;��˯��'�ď�}O�~�Xn�ӽ9��&r��������iK���ə�G��E�B��4񀄉E�>R0x�p���IC�b�]V ���OQϸC�C�zE�ı/�/Qd�$i���_�CӴ�s�O�\+�H|n�фa����%���t�(X�N�44�����h��E�axu�תHN�bR��2�'��-�1��«p�xA��s^�]IR-�8�߆�z�g��?��؏߼����A\�sg#��>Ш�t�^;�l�~ŁR����8k�z)2p*��bWL��F�0aB����ԯ.�o�.���~��w��w��wz���x��W��� �v }��ռN'�*/�|t��`g�B�0'�4�6
�Z��JE /a�Kҵ���~&!Iz�-�\PkPSb��%� \�!�x፛1��R]�v5�Ee�n�-|�(��䟴�Y�:�����s��d��D�xZ�p��Z�?���p���?iC⚤�K�'Ƕ�3�l�1 �ғ3����l���ok@'�"y����6F���.��(�#�o�-
�L�A��St&.#i�� �+�9�U=��;34���8�΀�ƹ2��	�.�Hi��L��A�Cn�189)����S�*@P�����r�8(#�Q��7Q���'��p��>�q�b�)�@F��n5�,��D䓤�{=��
p=�oL?W���X=�t�D��j
�b���+T2��-��iS���k֤}��(���M�J�
��s��Duվ�9��#㬊�h�Y�/E���[�XA1Q������\9<�5E4��Q����Kv�S�]�\�璐ܖDG>k�Ɍf4�5���	|վN6�sY�e|��<J��إ-��caN݃�3�!?���2T����A�p�bg�Ф��z���	$�xM�b(%Jo���H���VV��[L��`ܵ?A�v��9tZ5s��F�Y�����C���tӧ�˷܌�/�;Q�M��v��+�X[��� ���{0��QS�~WP�Ng'�Am��`^�q�%���C�qj�4�}�5��O�=�<��?�w�s(����T~���8.������Q۽��W��J�=s0�m�k�嘐��;>9��� �W.$=(Qi�d�mM�tN�=�T[	{0r\�{0*f_�NI*�F�2����V�d�RN����"wP����=�Ֆ�1��Z��W���n��H�w1O�^�(d�F�5�O�H+�&�Ȝܰ���:*_�"��\��/Yn����'F��a�q<j��F�g�)����K��C_�01�QR���#r`�%��l�u�é�s����O�����ᶫᦃ����`q��``v��	h�U�<Za?YI̚���va�T�8vz!=8�^�w�y;��_��qۭ8~�|�%��Ï��W�����6o�b�D�(-�0W�8#��u'�*Z���s�5����!(���CL��󏄬��5���t��8|A��t\&��L�u҂�H�+O����Y0�x�J#��r�"!2��Fl��e�(]����9?�=_Oǻ��N�v}a���;C�@V���`ݿy-�9̟l^��N�W��3�R�g�﹬�$i���rC%<Tȝ�����i��қD�hF3���"uד��n���.�ͭ��Ѯh�(�Y�d5��Ԑ�ַG9����)/�(�o쁧Gx#�橧첱N:pn<����qLq�ʢ��i��F�a=�S&VI�22��1���<�?'
�6�R�|1�ܚ�'�)�s(	�|�1*E������Q��;�������_�zR�״O�C���q�..�E�FGmT����z�t���&�\���pi�a9��×B�;��������R���:M�c������I�!cj����y��cZ��_7��=��f�C����g�G�[��k�K%m�&5�c�����M� M�j�-Q������x)�۟���p�^3K��Gνqh���hF3J�^���*�\�זǒ���c�H��#
��t�����R�ׅ�(�vJ�}i��A�����u�ߨ^�\�>#����o��5�^WӜ)aQ�V�S�6%I�%���T����(����0C��u��K3_K]�(��{[��'?�?��q\r�v�x�%�����c߮�17���l�����ID{=E��s���;*p�m_9�0\�SA�Z:���O�߇#�����v'^}�8���Q|�������ݥ�W�ޢ�s�*M{&:�*�s��D�lߩ��ڕqހw���]��s�J�QN��(Ѿ�n�Cpn����ۉa��{!�P�D9�!���S�4�X��M�dޑv���u�ϵv�������]_'���ϱ܋F���̼�r��h�1��
^Q�֣C���=a�)A-���Cr�Ŝ��}q�<�:JE�"&0�p�Ny�H�)VIrB����i}�d�--W�b�c�8��.D]��PA���[�Po[�k� ���3|�՟a���q���ū�sG��Żwck$J�@*c�wQ.l�ࢶw�)�(�$���zHc����7��0_��;�
�V�c��}��½�ʍ7�'��3��Ǟ�S���7���M��⢽NΔe<CS/��nr��&�Z�1��=����b(jNq��@ǠE:Dx1U�����J�m 5#�+ғ��؄��d�� (ܫ���%X�>�kJs`
�̍@�=a�+8�A0�vt��0A&x���l�V�b���sp�������E�䙜����V�(>U�C�wss�/>]�\P��R�bI�kŽ"ת��\���盒6�R�Ѧ�N&1�FY׌2Ό��3�)R���HV
�c����D�Ʊ9Y�(6�8��������I�Vep����ɹ�^��웗��v-��̣��V�垛Q�Qi(��9�E<���f����.�eDO�NZ:���YR3��̚��B����� ��iCA{S�o�P�omTDl�#�P�5�t�h���N���.������K]��Ѣ/Z�4��I�Iu��V#Ʃ��\��>z_��~Ժ��R�E���t�)�����c��=��B�s����ڂ0�N��(��&O2Z�9*���zJ$P�g���������x�:�P�ãdI�:��fk�M���|�{��hՖm]����1���0�0̸�1��G�̽��0&3���M�C3�,Ep��f�b	g���W_�8])�9��$oٖ#��c_[��yVy����Gn��"�j��tt�m��q�-
M�u>5,�g��ӡ΃�V����u�鸡{0Cy�.m$�G�g�˪��a0�?-���3m$���;�����Fo~Kͳ��%=�$�u�(�,,��K���k�ӗ_��w��B�Ga�D�?�	_�Dx4�`��DW;Zj���Ӕׯv̟������K��;���_{�>�4�y�<����$��P�4�r��
MQ��IA���!�7S��f����H.�^6��ӂ}Y�q���q_n&$	T�]<�H��W�'�>
{2b;��L�r�/r{����ڣ�ܑ6�<]⅏o��S�s�G�u]9�\D����DjX����?mb��B�6c7���(���Q�C�j���dy�Ǩz���PG���M�Q�BvƵɩO�7bIP�twF��G�h�/J�!��]��H谅Bn�y��Π��^w������ණ�3����V�k �\�ݲ�7(
7[{!(�!!$M����~�����&�35mؾ�ǎ�{q�e�7��,~���x੧��ǃo�����rse��a	E���:oP#��}m�mSg��C���k��;��q`�=U��Y��m�mMA��1���*z37}6�4n�^Fj��x�)�����JA@��H�Z��� @�p*__�~�,�H�0����̡��vJ.�A�����h�,�Zɶ��X����?�zF�<* �}pS"�;�O��&wX��AgV�hFS�h-����HZi>Ӭ�$�u�(k<Hd�����=�.VO��F�a�H��<R%5$NF⹢��X�̸<��y�4��kA�������&P�"�C�lDF-����	�Ė{-�E��}6�q�a�\k���rL�ZE8H���P��/Z��]�9r���_�s�Y ��ïaAG{�G	������Ѥ+�~��ґ����:�~O���}��G�D�,iԣ<���`n�f��|���/�4S�����1��wP�r�PgY�z�C�pQ�/��ߖc��g�$,��'��������畭�|�F��<�u�H�51t�|�v�ĜÄ4�=o�3�T�<I~�:��Ǐ3� �5ǘ+�{�(Ê�SG��5�#VH�Q���X��0D`�D��6�,],��J���;�&_�|���,��1\�8�q�ƤI����:���Q�)����0]�����@@Zau>|��NDU��J��R�kl�5c���ǡJ�+u�~��S(���K�8 ^|�U|���o�"n�� n��n���ٹ���� .�v'Q����!U6�~�_�iо�� r�P�%.h������W�w?�Ͼ�"~�����#G������<ʹ�?S�:m�J1�+���Ʃ�p��.��h(B�?[s2�e��o��JIHE��Ȧ�����R�(g�P"d�9��#1�TNϒ�.����0.a���m��2�F2��G�Qf�<�MwJ��Q�K�lU�@��G��A�_��I�Y��֍H�GDwy}H
~i�^O`��8�Q�9�
�8���{�i��A�z��e�2�U� `���� ���4_+b FYۋX\�YU��W�z=��|���ݗ^�y�+0�w�?w�ո撋�8��d^w���@�p�چsU.Du�3�	a~� x��G���x�.�X�=� ������;�>�4����x����Q���\����M=˞-�T���#V9���(Ih�3e�
�d%3 ����&�M`��C!�RA�ڈ��>~G�<]쒡D� �sVU�O.�tx��J�q�Q�ia;�v�3�0�����`��AF������w7BE��UEQ=����k*S�H���"�����$yqD&�f<�C�#�����]x0�O.�����`MYF�θXnL�?��Vy�N0�)d�.l8T�z�D��ϻ��ŧ�=�(
�����W��Fg;���ܦ�㆑
(fMYk�ްQ6D72u��<��Cz#S�b�N�<�E˵F�t���IP��X����:��<_���٥wm��D�d'1�M�͏
�24ߕ"��P���h����Z��!�p�?1e]��Q�A�I�C�9:}�
�bi&4r�S](T#�R�wY�����j��:-�~KO&\/'����)o欔�U�"�(K-c{$eʍEZ���J�jT~�5�C_S9���(�z%�cg��&էܤ��7RJ%iE�b"����u�#[䙟�3Zg�JԖ����F�q�y�?�;�=��X�\�cĮl���s��Kp,�/B��=�s�x�Q�|?�S��� q��\%0Z��?d�0�L̫e��q0�P�g���� �,0wD�.|kᒨ�-Tp�R�߳�.����{����
���R�v�6W���<����j	�=�,����`q�ێ����t��`z����z�h�6"'a��>�C�ߺ�j��6�҂S��}�%��E�rէp����c<����'pףOṷ�Ơ����Cq�:�����+��BRԚ�F9�h�/"yM!F0�����32��H�6tֵRv�s�k��8�|�p$������=�H��srnqI�$d�2j�X%M���P��T�I�H�^/Z��$��m��ޣ���Eఎ���1���i2�ܳaʶ�و�1f��2��B>Rx���B ��:Y��=E���=k|+�l�<��A��c���<�?{�(��h7n��2\w�޻;�mA�DF�,dQ���U�:2��ׁ�EAP�B�=��s���������/�r;����G��s?��o����z8�+Q�M���FƼ^����x��څ�UR��>�I0����kn���0�RK�X6Qs�UHӚ�ʗ�5��W-��$���ěB�EssX�ICUNȷW�܄�ZwK��O�m�/�7u�h1�ƺ��o��ˉY�=�n.��T���r�XX��%��� �Sۗf�[B��H
�/A���<� f�]xP��.�*�]ƚ�9�F�:���&#χX hs��&\S,��U���T�H)�_�+�J3������0�9���.�ɀ���A�L+�P`�.YT�S�xG��h�;#�y9 @�kE�<��i5m�:ْ�/����3.8\�\`���L���μ"랼֎�!�R���-��׎xC`����D�1N0�B�%�?6a����\>qe�� �%j?.�+J�4N����Y#���$����������r,��Lj�7���#g��K�i�	�AnC^�G��sY���08�p��h���䀹SS��Ā4�j���XtӤZ$V��x�z9�w�~��ȉ0^���[K�����"H�umkE���V�����?�ߡ��6!��sP��O{1[m��0&�*�H3M����ڡ��+o�vF�ƹj�nP���ٵ�c��ּ7Fԛ�8�wdYb�w�.�F������S�������	a��ѫ��~�maT�@@ʐ?�I@��h�yR�Ũ&��`ARެT_���t��r-͕�(�|�N+w���&��D%�i�U�b�,Q����bΆ�TP�@U���@���FW'߉p�����
~�W
�N�����	��'������/�u����矇-��_���F�P�N"T�S�x.�ZU��;�Q�HQ�*��Ol݂;�=�/\u���_�G��O�xO��
�y�|П�����g��͵�Zو���9�x�J�y�0��<|<���㡦�x �2�z�}�Dl��>�~S\�.���[��H�H���D&t.Z����3��(ث9����C��d@��Z���F�.-.��8pL��yZ��ٴ$��r_:q�כ{!J��4�O�P�ҡd��t�C8�bn!�Q���7:��_!AQ����y@��FV��\gF��Pc!�����j�ך�/��2��������߉[�����/=�[ѳ!9*'�3�����h6��Io�j��͉�*^Y@��7���mW�{ￏG_|�y�I��O�����hh@��k�Ti:
ƣ��FymA	=���px�=�1,7I��l@R2��sA �)��F�}T�'�=T
}=�A��w�҆���Q{6ۆM0����v��	"G��3�X��e�i�y�u<�j�Ũk����%)�dx _��Q���ׅls&�R�`}�ss=E����+0d����� �����Mv]䌄gh���5#�9���$�Bl�U�w�𖪃��صjgF,����r؇Y���X��߄ �~ls.ℯF�� fw�a���j\�9{R�y���Gg�rD��tƕ���VJ��h��۹�V��AQ[d�n�'��rT�{��dM��@s�
W:��T�:���~c�7�i�x<*>�U�u��w�8Hk��e������ʉ[A|)�	��(Z�A�ݺѡLxes:ϖF�I���u[Wn�2��!�^+-v��o��S��޺���>������R��b6�� ��^����v�\��Bd8	��ِ�Zݑ�?8j8or�s$͛��t�0��B�C���Q��Wb�d�]'���ȶ�:���B�Fr�8#�t_����3D��8����#�݄j�W����s��i#���M1�x9��5ޥ)��6b�2���~+��#WC*���qd�L�9�i��0�UAk6]��X�>�����6l��v���*�$�#LJg��<�l6I���$�с�ő�VjÅD&:������!��)4�Oa.�ඕ!c�V�6ɾ�r��<о2[���Q���u%�;�z�2>}?�{��M����<v�
�wL�y��3]p)n���:�,���4��<��/�Ky�X8�p�
n��l�~�ۙ_{l�+q��{��i<��3��Ǟ�s%>�w/n=x	�p� \�[{��x���W��e!��6�P���x�X��-�@�~Z����x۹�����K7߄7N�����)���������`�졜�(�:��_oI�a��b�H�HA.r����a�*����MG�C�@3�N�/X� �)��s#�.Rg���)��^����c}n)���5��{��g�4��Z�a�q0�B)H�����k1�-�k�"�olJu4֏:Ӣ;p�st���jh3�uJ�c
�������jD���4��`��#�|2
F�nu=)�űcБ�V�_�&� �2ډ��N���j2>���M0�Y����F�b�|�/�H4B��S�?y������������篽�/8��z���m6Y�zڃ	:%�;B�;v� 
e�({�3��Z��Pp��9�����Ż��}Oş����'/����]F�u+��,��]/�67m*�s�	mf �
#J��(6uU��{1��-z�@��U���A�h6r��Ms9�a�S���kN!�-���6>�(ֈ��c��7���$/�}?F�I4�:
�;U�<�݃��i��-���g��Z�~Ծ���3��o'(K�c[�)7��όf���Zz��A1��6;� ��$[5cR�ҰF�G�2
8SG��T�;G0������Yh�re�H�j:ȁ!�M���;2�֕:u���!NO$�H]%r�Ɣ���sR�C�$��±c\J[��(k>��=wR��y�PbR-v���))2I'm��m�����G뙜X��`1]�M���R���F�D~k�3�6,s�C=��\}w]�qү���ʄh��v��p�Bt���E�	�݌	���w����>U�WЇ�T�Oi������C���U\.��i�(��D���1���:�N[g8#����*K�W𴢭��-,9>H�Q��νQ�5�����`s�`�]�g2��/�v���WK�5�rx�+݌�n�d��b�g���%I���tyCr�W�!�e˕���R�7�h8�o�m�&;�i��Ż����uTU�-wƚj���I=ƺ1H�3(�n����	�T���є�U�T�^`���G���1���ퟑ30�{��ถ^?3���Q�;+ՅK5��;�/0��o�{�㍞�ݷ��o^y��u/n޿�|�u���!�ݱ�ơ�8zWp��e�+�s�����%�ȆZ�1đ�k�]��f�Ȝ���q���������/�����	���C���'O���f�n�5߷{0=��,�^(�[Ӧɥ?�g�n���~O�{ߏ��}�8h_+8o����d0��-�μ}yVF 
4�q���Py���v�����$N�� ט�6%�N��g��G���h�ڙK��!g�́#�X�3Q�$6ȓ?3�R"���S]8�o��WZ7�pe,$�#rQ�4���:P�fdR�0P�*�!�0���l��!�
v�viJ�La�淅�E|�<z�����w�Ů�ĕ;w������×�={���� 1�ĉa<v�VG�sU��t�.��>6�}J��0��F�q�B_k@���^�W�z?|����3x���FU��>�{s��eT�A:66�=�[��o���7��B�M�0j�G���4!�[�pn� ������|�DhL�����*j�#&\<��[��'�� B�1R4��$}߫"�/3�����_V�3
� �8 K%������.~�#��7Sf4�u�O�2YA۝q.�E�"ӃX��J6̇���������\����;��׍"Ե?@
*��9�mv��!�O�,D��X&�5�p�4`t�&�`b(�-���u��G�(�Y�p��V.�ʬ!EuP\�ɷ���{$p�/&2���s=4�|��]���8�;�@k���1��&m�K�
�eH�B����Wb�9����b�Νر����*���'O����go��g�<�w��F2Wd��s�0n�*�+�y��ر�Q�hj�&�0K��61�q���-��ٝ�vP�p��+�Ws��a��!T�Sx�S�t�neO�!�n��=�Fw�M�x�崞�,�� >ݬ�����Lp�Z���0�xj���A���B4*��G{���i������6�6[}g��4�1��K�d٤��H��()��R���q��;p*�%��S.�E3+җƥ	m�g3����1e��ʆ&�G���Q�9�i"�6���{��v�C�^'��=.�^_�ß�ֲ�A���Cv�F/�N�v_���7p���ƅ?��w�sW^��؏C���m���ܼ_9=� ��G1-ؖ p|D���:\Oo�6i*�{X���.9o~������v�i�������'�œo���z��Ţߨ'���9�۴�D�(��6HQ�.�jE��h�.��jS�Yx��mYw�s��{��֤��#���'�Sk�zIҨ�L7���^ S̼1�N9GL�=�P�>�ƨ���D:�B�<Þ8c���'m�s^VQ���?�����O�W#ya�2`���� p�t9�ISj�X2�C|D��${�?��R..�g
]��o��zP�9�co`�7�~?~�����6@⋇����ĥ{�b��<��!c3�Υ��<`W�¢��gllS�3�\�3fvӢ��V.���E\���n�����y�(~��sx��[8�o�/�9�e�iG��s�T�:�Y�U�ΡN�J�{9;���斜��Y�A���Rq>Y�����3$o���0�E��;6	eT�s�5I�T�%��FN�CP֪5���E���i�0�n<
���n�R^��BQL>��۪_�Kwҹ�^��rN�3��f��I�L�?�����$�b$O�CtBޠ(��C����u�?�=�։Ď��D��I����Jp�*K�`�����iԚ��CШAk �kt����C��%;�h�K�ꟓ.��W[N�V�t�:Ú렇���ʩ�?�V��񿪱TT��o��ۄ��)~Oz$��R�|{Mj�U�s����T��Ѫ���j�1W8�s�;��_��/ލ��.�s�aބ!�=��[8SQX^�pr0�����ýO>��{/���Z`�T�/���M�m乫$�I;3��;�F�^A�!]�p���D֩�Æ��Aw�Uul:��C�3����Z�o��-��7E�K����|�(;ݴe\�޲yz&t&M�,Dߌ�r�U1�I��"���
nTmZt�p������Ѧ���jץ�L+�����3��hc9D�&F�rot`,�t;"։rΞ1��Rڤ�^p�u��8D�X
߭���l7%�h(vXOH�Յ'�t�&5�>D�s?�?I6�M{�V�'�Z�(^���9�r��6E�4��=��Q�kV^�)�����W^¹w7^t!�|��z�2\t�.l����[�m�j�,���A�J� �2v�X�Q����gh��/�s�|�й�����/܊��w?������������^)|s�P9'^���q�*�?���Y�k��[K���ϻ8�
]!�G�f�{[m��Q1��Y�$�5�Ȫ���l�^����q�9g��o�Rw��
I�)�E8m�q>t�-�\䋍p�$��$�A'oY�|>�.d��Y<
V1��u��
�-�.�U	�FH7	�Q(g�߁N���*�C��]:Ef���-J��
�A��b�%)�&]����{��!���ݻq�U��k��vc�ʡ�y��"4��W��K!I�:T��o6�kR�4��<۽e������uW���?�#���<�(�� �
7/.��s>چq�P��E�>м#�rWk�x �P7!���x<U\;����x��dj'(6�S7��{y-�gZ�pۉ1T�����n�mF93x$�_��%j�:.�I����s{���2����a���ܭB�P��h+���$�!���۪����掟�l��6�6%6�|1t6)�3���FQƦR�����f9�քG�<F��Of���Ǡ{��3V���'��\ͦ�q25�k��b���S+��l���_2�p��DN2�������zN�Q 	/���DY`eQ�~�z���r�WVM�;�^��ЕsPSt;�X�jЄ�EY~]��J�P8oa���䣁��0�������J�f��,��Xzg�{�)�K�7�up01�%z��j��G�qp�y���#��+pI�y������}�ZU� �Mtb��):�CT�z���z���a{���u.n��>�x���K?Ã/��{����}gy˜��e`��U��e�_)���:��V��Њ��O�E�/�6֤o(�6l���ZzP��nd�3��EU�N��T	�Gug^'�G3J��*jm<T���(�\�8O��ɶ�i��$7��Nxb�wg*��w�;��+3Q�qJ���5�(2���[�0^���0)�֕Ѥ?��á��_LQ�M2���hF3ZjE���oN��5-׹�����r�NQ��]��X��ۈ����r��*}�uZ���`;��8ل`m�&�'c`���t�CtSwU�KmJ���}��ΐVKa�}/%y�-w(�eI�ړ��	��^f��n�zK.}|�#דl������,��Y�X�+�)��>�p�>�+�i�����e��P'�o��껸�ſ�ޅ{q�������]��;�氟�7e,��Ƒ�&��+]G��O^~T5��C�����Å�ĥ�m�{v�럽o?���z���ĉw���}�9<[��c��S�3��gJ�e��hT����2uXnF�ɔg�1��5��C��p ,�Xo�w�Am#�ӥ���J�a�p�B�+oB5�y�a6	�ǉ5=��h\G�8S.r{�R�1dfH��K�F�&הb,�b��3���	HNj��h�7I�WDِ[# ]��}�2�Q�I#G�dD���S���mHf#��Y���`�\G�.חDnT2���J�*֞���e3ߏE ����_��t���\�ei I���ě��]�����۶_8x w\{>u�"l�_�����\�oH�W�0��8���o+[Z*��ݩ��޹e�����O]���{?�<�������/��8մk~˼_�&���U��Xm�Wmd���ǘ�U�E'��^�D�X��	*G�>R"��nB��w�3S��%���_����9���F��m����;]鉀O�r��e��^�+���ȅ�3󲆏h�+J˸1�YHG�.F@M
w��w�Y���X������,j �c�̓DA����H�����dF3ꢍ0�'�C�>�V�*��JYEFr�Ӛu�L��u�ߒ��?l|N�B�d�f0"���m[����0��@'j��Ǟ���F��Q��\=e�M�c�N�{(��1k�/�ӣtc���iR+:X�#x�C	��V���� ��Tqr�~3�N��H2�c.�"���YWt�G,�p�������͇��R���ko����A��M7)�گub�e�� 86LS�j���_��6�w�O���z���|�ї��#_��d�|�QU]eP�.l �1�:쥅qIDd��C�5z���c�n�{!~�����o�O�/��'�&�b��n
4K��Wz{���.��Թh�>dC�8!F��^���ʵu}��J���Ll��O��k-0�X�$\ꘅli�T��5=�8l�r]�z�z�f�وo�Bp��@kF�(0��8C��\��+�8�bP?'+�,��ޝ��C�4(�L	���IHsD��­k?��vUaj�!!^Gc�p��ڌf4�����<�d&yFW��4�=��K�c��O��A��n+�[�Ⱦ�|~̟���mg�����s��Q� +26�:�zA�o�n�I��7)6!K�N�{�#��	z�MO?�Ȼ��4�$d���B:"$LB��X���ǸM��V�aU��C��h?E�N/D?��-#��L��A84�Nv�c�r�Q�(�q7�~�N�}������^ķ�{�.⊝��KW]�ۮ9��v���~�y*�h���V���!�Gb{�#d��k�}m���"¾]b�/ėo�~��	����62������
Ke��b�4��Io2�̡ߢ`�˙Bc��_��*�ܞy�A'�.�aB��J�$T�WQ�|V?B��(����하<ÜLY������햦�~|s�k��rN[]�^ΉC��=�	���l>�e�(Z�G��Ev�mX�*K���8��땎�Mᕦ͍��3��b�_>}�=��$H>'���3�l&�����7i�[�.� {ݾ��c�pY���^`����qc��w.���������=t��ۍ����_z)�=;�,�l��5�X	R�%ad0��r����\墇X�0����$<�\�k��-���co�>���:�ǎ��۶��慅��~<��N��F��jQ7��a�X��i[�����&�H�?K��;�V:-��ޗMH��8�i!�V"p ���tlKT�#��*k�yk��pa�i��e:��4Qc��J��/F��������\Hk��ҡ�f��:9O砫�y�AG�=�O���ь>���RY��,0���3b��΋�~N�S�M�D΍��ܗ���:B����M)�/�Pr4�Z�`,U{�S͓�Ё1Go��-��)��N%�䉕��R�:n��2�`��WC��{R���a��\7�=��zQ��G�V��h�vq��'�3,pŹ�����U���`k9p8x�Ÿ�K�����΋��ƠAN}eu��~�X����B�nA�}j�3�Uڝs���<p(mмc"�����u��_�:�r���+S�%���W�Bơ�Y���c��>���F�1���w�����k�ƿ���������[�{�n۳j��³�I]����=!(�JL6b*σ����y��PF��ǧ�x/�|�G�Hڑ�飢�d�E�s+��ИM��6��s�Dw�J�N}�_�ʜ�@�U�7�j7�j����8�+�Z�����X��ຑ�����jM4�B�5R���S.����cF3��YA:a1���fu@��s�����cc��Ha
�o�r��gd6�����.{e�_����j���f�Ӳ� ƫ�'��*��������V�[QmBn����>L��<xW�3�Eɜt�L��V����6YYT؃Q����~}�,�;@k��+
��`8��8<�x�U�v�5��|�-�����o�n<p1n��
\w�~\r�vl���Z6s���
`��$vog`Gj�����`k߬�Wq�������K��}{��w܊G��~��#���������hq�
[�:��ʶϔW2�W�y�C��(�z=�qv���
	�L�9����D�ٖ|a��#��vV����a�y�:��>_�ϴȭ�	�nrZ��`�*�d3ڈ$||ґ"C˴iM+�W�r @�}7E�$��}��+����F@(����_�.$w��ا�w��@�I`�^�*�!�}Y ����ӅK� ��^�F�8����O_�_=�2v��Ю�������#W�ȥ�`��-�æ��A'IE��D���u	'\��[��X[OP]/�߷��x7����x��wஇş��}<�чx~�u�Es���83l^�t��
��2��� C(j�E��h�I�%_������91N���"���NO{Ks̮?5��e(K�"Mc�W�2羴��*�Q�p~�.��=s?OT+�L]T`��$�\��h�7�v��f=��Ԝ�o��A�8�av/gF3���Mc��8R��"]ge�����!�N��j�aJ8-8x��Mő�\���&�4�(d��VY#���4���Ԯ���yc���<���cI�������MFR�oZ�!��P"=G*)�e֔H��]����ji��U���_���_������`ɪ;�݊��_ƛ��/�_i�K��[��?�u& VpJ��u� ���]k�3�u���$v��������[�Q,DJ��rݕ$p>�����z�u ~6�m�n�.����_y9��?�}|��{��܍�O7I��eل7nt�&O�5x�2�WCE'i|",ƝU�N�uU��X9.X�+��|�'���wj��k@�S��J8��q��$��!Pq?�|��K�2�A験g�<��B���k�LT��E��9]Յ;J���A/^iX-��Mі+�
ڥ(+��b����@��H�O��,5������f4���b_|%HH��7$��8o�ƕ���A٠H�?j�� (gO�$��,�=�����vC�~3���	�aF1��l������SV=|Z��$3����_������.�-��(��pk��noC5?����Fe1�q��qh�C'��sa�#��p�I���%<��3��Ǟ��ͳ�/ڃ�>�/9��{/�ֹ����%|�`�C�D���@�	��A��у�_Ťp^��;�9�;�Ʊw�Ɵ�ݽ����sM9���0�X�,�`C��ڪf�X��`�.�6?��ቖ�ҕ6L�GE�3��;��ꕧl���1Mlb�y�ɒ+:phj$V��tM�z�<zFS%�C~י�'4h�{�v͍�ffØ<��o��rs1`hY�X�{���s�A嘑9���CH�~�����%
s큆��Y�w�k�4W=���4�M�~K��~�������O�?�.ۺ?�A����qe*Ν+a�Y)ܽ-Vn���oVS��}Ӿ�Z�{�2�7��AFJ����c;��Wo�w�|��������k�X�-�_�P�kb��3	��=�M=O�K� ��Rw"� �	S��^��k��t�!+���&�.>xP�;Φo�T�4tA���p�".OE�sq+ʲ@Q�V�EU�(8Ee7,�n�`�v�W�U��U�(څx������&Tt�܂t��G�v��y�R�2�ӮFQb�l7��|�RT��2�WIP��{���/�?��ɀD9������d������a��I3,�q�]i��j�J�5�!,�u�@D�R�{��<Er��}xDs3��i��׬���ss8�*S�t
+r�TT�_ђ�E��esnbkġ`ö�|�&��a[�	�Hp�AE�$��~��i�	���T#�Ӕ�,ࡌ�VE卋�C�E��n�C��h-+�����Z�=LGbloH��$�%�2(#@#���@9ɉҴ�.&�Z	]�<�>:�/}�|�ȕ�~Q9=��7m�+l�~.��q�{�q����M�%�C��U�}�H�}��פ�=��r��ӧq�%�}�Wqӥ��_^rQ7l�{�dȌ0�/%������X�&:Ɔ�2g�4��Rرe;��/~��>��g��_;���&E�l�W���ke���4�!��?��_�i�����+W�09�x���+���ܚX��b~F�S��͒����$��)�(�,Ϭ�."Ǭc�uB�Qm�Γ�ݮ��q�02��+lT�ʏCau)��!��)Q��� Qњ��Y��h�#�~��E�Ou���y�yX��@s��.n�Nn�.x��n����^��kF�� 1�<,U�:��ǥm��Z��zOR��u��(�;����QԎ.�:�.0��i>���f��#L�[��bD�t���G�=ݴ�:�J���~�A��}O-�ኁT��:wV�O{%,Ө�Ae�̠�l4������;�#�#�J�^��Xg�*�s�5D�2��S(�P�?�{-�'؞�Kp��`k���Na����]���8s���y�nZ'�Ub�t@TkZ�"S5��F#�	�t���8Q�H}1&h�0*\�D��{\�:XK��O�������&�ZSk���b��9��+��'��y��D�G}������^�����\�_���z��۵��LS�r�>[����|�:�hLІ����B��"�n�w.�9�4u\�ab^|�y��_�*~鋟w�_}4��2�v�+��a�,X�~�iZ�$�h��)�C�<v�i���o�G�, �_�'� (��!Ԏ���ӂS��-b�;��W���O:p(�]��[
�(�!����?�}��iwbB-s45(�"{���^5��A����<#�F(P)xg��D i�;�-+��b���/ٰf�Jn@��=m7��VS�A�Xa������iS��,�ú�#�*<��'�oxWl߁O_���|?�޷�!z6Dp��3!�z�T{ F<5�2�
�Q��
�4�2ǎj����5���}�kرm��?���=,�@�P����m��)���x��sv*&�)7<���*�|K>,���J�p1���ar��L�O��i�~�©�����9)16�um6� �zU�*{���*e���vW���@j�z�{�Z.�ng�+�C*�v��ֻ4�*���
w���N��z��L��X�CY%@���d�i�j�Ni��ԩ���6��E�I3c/r��Ɠ�壱x/�=�t�]Λ4��E��x,<���W&�q~,Rn�>k�[i��[w�W�b�G��8NYj�m�.ʇ�g�t�ӒDk2����{%ʏ��XR��W�l���³��hR��;�����Sg�#�?)_fْe^.[>T��ü`�Ni�����F^v+紩Bopn������E�j�+�5N��Nj��-�/ �3RЭ���<��Q�)�����Q�^{���F�<�'�t�߅򧃵ߘ�Q���*��5���ic��^�j켾4JYI~�I�v^ST�5�e��ljm��É�C���dy�t�k���j2i�*uO&���k��e&���d�K��	[�>��%:���3s����O�u�>��|�y���l>�-� ��uo����م���c\�n���z5k�+����~m��m���cq2V����p㩂l��we�4���tsO���:����+.��{�߿�W��?����&<��4W����)$��\���jś���7[�L�! ��m6�l	��Lm�1%�?;��%#��-��@�o�O��]i�uhS�s�����&�����h�%�UMo^��� �����8��a�Ȑ��Z�
w��	�m�MQF�1�L��7�G����֡Լ��䯫!9u�l��|R�h���B6���^@(�W���1�i�=W��=U�B��o�Ir��q��bO��殘QB���>~WʂBZ��utC��b�	D���\�	9(?Qo�4�����L
}
qm�K��SH����G��]چ�ia}ѹv�$J�Y�a��t�v����it��8:�x��>��ɵ+}6\wt�1��ßf=S]�|��,�(o'�(���Hi͢#%*�u��yʸX�Wqr>B_i�%����}i�*�	|�0?���*^�2g�QȨ]Q9��b�l6^�����vuE��¸��q������6��ڄ�3�I&�t�9>��G��t���Vm#2k��^��l��$Ǖw4U�	��z+�dw�j�\� �ޛ�+�hV�m+�MS���#'�
_O�뎟&˴� ۹���#N�2�W.�t�0��l�D�,��A<Ej���Bv���Ҽ%AI��8-�R{�oa)ʲ������iԋ[p�����������q9'n�h>sp?�ރ�;w6�|��ϵU�5u���x[��k�
��$M�#E��=V#,k�m��7�<����-l��/������✽���u�Dc��=�t�0W��ޏ�X������VBFg�;�Tp̷����5�Ȫ؎�C�&�A����|f#8%�EJ�/R��*.���ߦŗ���Ix��8t����G4YV��g��3�D	 �0��.����i���k(1�h��k]�j�_�?�r}���;*�U���&S��H1�ϴҊ�˔���mo(��b��mkXɛXƉ��}O��=�$�܊;�8�p�ոt�غ0�9շeX��2�*�0b�w�A�@��	��7��:i�jl7J����q������G�>��L�^�'B/}�s=�9���1D	D0�������I�B*��3��� �1��G������A�&�c<`l1uo���P�M�8aŀs��}�"W=����D�qK�(ʺ�'��D��P��k�l���RY�&K\���ʶy�a�r�@��9����3؊S��oyҵK܅��)iJ���"�)jr
y�ʅ�],��RA���;-ƪ��a"%7��z�э��a��6ͨ�@%7��+��4���ߐ&T$�uX�v$*�sO��>F7J�3e�4܅C҄v�rG}�Ц[i��|߯���0OW7��v�R:E��*��w���v��p[�h�T<��ߣ �� �O��Ù��b����v���>
����k������c%�q������w!e��\�M�z��Um	F��kB�n�j��R�}v���ԛB�Eٳ�b��7 h��'M?�is�a�}]6����?gW�N�6����V��i
	~>��6(��nq&(u∟����<���}�G�24�l����������4��F�|�/K%`�lA�qLX�2�[=�/}����VLV�kC�$����3�������	vP0��$�r������س�,�HU` ~-Q�����֙�ہ]K<#Q��Ybe���:�6z�r��M�����O�!����C����]9'0�*�H(FaY��^V1�ѡ\+M�c�[FL1�N��0$���y��!��}p:h��6O��(���^-M�C��z>�����y%�;���Tё
���������f�-�.���Z7�5ȣ��`�t��x���V"�E��.�o~إTY��uh��6⌍���+8}*��S��~h���;#¼s�V�h�n�����c����m�ք�`��ۼ*�RGDX�k�Rc�)�^���pKE�J(^W�ˀoԅ�C���x�Ol�i��� |�pu��ܚQ~�ÓAQEu�.BX�eN�c!ˊ�ĳN#J#��I,NC�Χ�c���q��^��@i+��G��I>*h�����~-}���Mr���ʉ�*���E<��w�l��aMAfN�G,S���,\ �����zqؿ�<��Gb\EO��Yck���_Gk�L��;�7t�7�j(�?����sq׵5��$��Si_������|�e+�����G�z��l޳�%�s�wNv���j��:�T�l"�6���%�(��8Ct�$�(ݫ����z���|�i�y�E��8i������a?ʬ�JG�%�<sh;���%�|��5����ۆ
������X�u��p����?sm����K8�W��������?����W��w\u{�ہ�~�F˰��J�H�l�CT��:�?�tF'�bmϭl_�8�\�����;�o_|��c�"*��V����z$:��"�z�}�eF���=�,�Hwt+y,(L��������X�9��}��h�J�̚�_cZ	7:3�:OR��E��r�bF���7�C�l��FU�����+�/"ՑD�A9��	����H�4k�n��C:YORXP^��u�*�wE ��*�'659F(2~:��v��!�'o�;�$���4�{8�ۆ��zx����G�=�C���g\����������٫M�vTzɃ�p�������F\�`O�����D�Q����x����=��+s��Oi'���"h��E���y��s>�A؆z�+1`�sY���xN���u�8�\"+Qi�Xo��L�Z���^�l�,�%��Hr�^3p#�k��؍M��YS�G5��抭��]���qz`6��9�`כ��%�@gx#��B����.^�O"�d�!��B��v�hfQ����N��P|�ͱ���iu2��˨�H��ȋ6��ɏ:������Zba�3�}T�e	^�\~Xh����ҫQ��w���n&J��1_(_����<f9�O�x�#�D>�/���6UX���υV�Aſ��@h;���3�+�X����=)������>4 n�/�	��	y�ă����>�"{��X�:��,Z\b.�Q��\�KoB��;r��\������3����S�Y9^@'<�B��7؆ӟ�7卉4����F�p��.j��J�A�V@s�+�ѫ�cU&����t-��lߧ��#u�cmԢ�ª|���a���~o�d�gM�3惴AP�8`�9��hb��L=@�\�Ք�\5���Z�lhR�C��>}�9��*���F�v/���6&�X\�	9�d�e���;����XF{^��DmA���aN�m�f��>��>��JTM�LZ|&��wn�b�F���-\qD�F�t�f^@p��'�)F���x���'O�=����Ğm[���E��*�>�&]�-/.�\����y��L����������˰v`t���O��Kx����~�[w�+*���N�`J�O*�ff���f�F�Z��Vȁ��*�yrvr
��Yj).U�<`6i\T���	�	S��աl(>�_y�yY�ot~}��6���L��:e.�\��Lϟꆍ�U�X�:��v���J^����m�N5m�.o|Q:8��t�Ѽ��!u}�y�Fb)<��Ɔ��`z\���y��W���Y��2��`K8�����egMю���R�s�D��}Z��G��"��&���H#�:�&e�j��"�K���QE�#�9�T���}R��4��x��*uɍx^,.�zK�u��i����t�.���ԩH��}�2��A���:�a!�\���,��uVu��������Po��h>(�qf�	q��
sX�B_)��5P�L�5�Ø���-����~}�BWa�ʂ̘&{�O�3s�T�̮k�34O4�i��!�����V��F�(���E��Z�>���W���{���*��S��e��]d��,U�Ȃr��<�S������hS~�6��̗�{�9cU9
��y�ӳIs��S,*��\)G9����L�K�u��� �G���������m/�lѺ�d�q�]��]�|Wm�t���b����I��Ǉs���{���c8��Gq��ݸ��e����g��?��q���?{@��%��}�m1�ŷ��v!�t!�\$Nc��n�������oXTɓ3E{>DC�i����:Tq�V��1"n4	�7�E��`8'�@ߵ�<+X���Z|�)ZLC׾#M���+��E��|nڔ����<Z�&tః��F��5�6e�'&����1�-畕;9��4��)���Iw?�=����Q�N�#���t��1>)�A\��w�<���l����E߀��)W��xօK\�e�U��&�;��K／��4��}�`wo7_����k��#W��3aÖ}��	�pN	�M��[�S`gR�̮���4e^��B�:�\��·.��9�"���\O �ҷ�CJ~$��:z����C�4�( ���FyIңuh� �I8}O�CQ�,.�<���]i嘓$��P*�%����F���7P}�@�<��d�z�l9
����}��|��8�"Q�i���MT�ڵ���d�Y*o���7��Q�(��L�����T�_� Ҙ�jr�:���l@��2�RW��	y<�{�2\�6+�0(��ee���U
�P�5Cs�����,_��f�KMk�P�J	:�G�.�|�sR+h\��×[�qv�ȹ�y����,n���0fAR>�`<�y<B4?�f��s[�ߴ�v��	�p��uX�1sbEW��> ����t�ȵC��q�}��=�i:����P,5�.�����o�ƣ�4W�;����_�v��no��1\ֱ�����S;j���*�ڭ?;�;�P�ۊx�=� ��҄��w�Fk����2{�k0�E*S u֛��z�זG�����Pwj#�V{^'��(��y�9���A�c�	�?��d��c�i]�&Y����S8mN�8�cX>u�E�9^ȶ���	4���b$5�q�Lv�ԣx�HZ��/�[C�7R��B���/���H��-�P-�Hai�����iZ5��n��Ɯ����s�JeӘ�}mN���C�0�;Ș�9섮>2|����FOX��44u�����+.�	,]d��f�������n�(���d��B�.tU2Xv��L�k8�w>2��)������x�����K'Poي9UZ��Des'��YǛY\O�g*����͏�MC՚Z�e�a
�)�:���x�wH׎̃Ah#w�ǧ��\����!U�^>~�M���O��Y[~ݬ#���zy�u���I�%��I`!�?{odّ�����^-ݍn�Kc_3����Y8�Mq�RxdI&�`X�~8��?��?a��V8�r�"�p�B�-+��d2Ds1i��p8��,�C`����Xz��z����̳e޼o�W�U�� ]ｻ�z��wN�<)�z�Z�~�ɑt�p�d���Y��v+��G,�qx4��͌Mqe���1���e㑗�K��s8�Hw��T]���:8��16JWq��uČ6�M�Xv���iA��i��.uRf�G�S	 G��fG���`/��aP�:u�g�O�6�>�z�nB|Ұ��$u��af��JNx����o�w�N!2���:�+���1-s|�ߋa�K���B#N�M�c�D/��5Y:���?L�"�ic�'�J�?t= )�c�\�!:8b�F���)yLԉ#�g^��#֋d���dJ�{�WQLD� /��kO��^��r�@�#�T���/<ږ�cձ�����^�ܦ��R;̐�|��(e��o=6[/�2�U����/_��{��h�F��n�8��9h�m������Ë۰�tӂ��+���f�d�.?�e$�)a��.�L�oW`5�>�է��%LYZ'�S���J;���D>}r@6�,=�q8�C�L,�?����<�9�neę��{�~��{��?=��k�ml�/=x���~
�?y+pߪv"�����+Kv%�or�wQ��k0�Q��s��>����!i�����~XN�<�����bj���&�� �^Z�[������µ<p�<8	�J�i�Zl������N�=��˵n$��8G>��5�>B���t�9R���w�L�Of�+�X�K��	a�2�P�`t����-
��m�1E��L��}�D���o��O���x�&,NP9���R2��9U?�c6¤�;ܼA"D(�����6l� �í-x���ǯ� ����*<yߝ�|�h�����*)��`"���0��V0pk�yd ��8H�|e��e�=�;�k��r\�N�&O�oz��-N7�QT2��"Y��zH��c�Knv�g��v�$��Ɔ�Ax.�Ju^db@E?tFY��μ�2�?����G�n�>�F�K- }��x�(捎J�,R'Nl���I�ur�\��
��\d�1�8g�@l�(��h.P�84KE9� /�{e�����
�e��Rڴ�J�7m�B�*%KBt��;�>�ԠÎ,&��2��3 *O�UƓK_/�^ q4�0U�ƍ���T&���q��"�t���c!5k�C���22�Kb�����V;�t_Ѣ9�b���R'uCx����Uh5���L$6嚔]n��o����Pn�>� K~�;�{VХ�5S�ZN�:�Fm�xy�Z�+��&DŅ�l��=�yC}7�u�J(���5��%�`)���H��∂�k\�w~׬�Oe��3�9ۏfHm%�1�N�r4�S&������>H7Ф7B��u���l�7���>F��Z3�K���7�A׸Id��l2ō���T�9��I��fh&�ր�+��υQ�yC��ӳ�.���^ַ<���n#���K']��6������Q��nx&���7Wx�WF��4Ap��*i�፟M8���yt������|�����\j��O��)�y���������L�E~��mǻ�����8:������ӫ��m������W���O����5T�0��L1q8�:�5��١�Z���ܦw�\j'lH�:�Ȣ8P��Һ��wU�O�	0]Z��}�����`kڭ�+���r�����b���F�@�����~_f˓�>� �����z6��$F�� ���#p ���<b/3�hSBD52�A&���x�}��Je�WCNA�ubg >�'Ϳ�L�O�2�'��1:y��g��xhJ�\ �S�sKn��&.���FӒ]�U	�D��1f�g�Gԇ���'�8G�+jWr�%,L�c�>K�'�\����Ǥ�9��.4WgmM�9ŀ��x�Nl��, �ed��2,��arPm/M���Gut%H��v2W������	����o���Z�iI�5d���7~�M	��X��,F͑�\���Ʉǌ�L����w�j�8o&�I�'���{���I�h��T/Q��]��h��E�y rba�B�(o�����Oat�P(!�610NU�Fͅ�U)�;�8,���V��1��5���o1��WU��h�kP��6�����{�'p��!�6�d���e�	��㱒�&�V���.��*�]ŭ  ��IDAT�͋d�I�*�Uݷ
e�?���\��dʻ����Ʋy6x>�ͮ�Y�'Xv)<]({ɍX��gC؂~�Uq
����9aN���Π�s��������'�9{^�Ʒ�ޅ��?�
�<q�C�J����� ���>��O4�@��pdm욯[�G���O�S:J_�ϐ<c=A A'�i�;t��c!{���������C�<�@w\V)%�1AB�!L/�v4>�k���>���,�pg/�7����PƳ��;�ˁ#0�-]���b?�Ed��CȲs��7+�Y�Y�e̚��	�u �lX���TX/B� {�|�Sfu?{�d,M(�	R�'���% Z��+�j�����Or��&:o�����V_>�8����w��t�S��ކaS�ɛ���z n:z����#�$O�XF�i:��N!	�Sݦ��iS�E/�>�h��X1�t�G�.�z�<�{�"��$�f!���N�o��2����У�|��F�OM�≿?�x/��l��2�8���q���h�� dt
i���V08��7m#������n������s�w2���؂\U��ڸ�]��Hv����\[2�荱�ۄ�,�~8�;���e�u�dJʛX/�s���Ϥz��c>���	������ty��U�!�;$�k���l7�9)/�.�I��N=p1?�:��K(G�>���`�=y�g�2��KvOޯ:��m�紴�2�4m�,�)�0���}�ArH�tޔ;׫����7���nP��	6��+|��W��v��p&s1��iԨ��p*>��Hc|(��"�ڔ�VV��o��9;[�f��1b*T�Y�+����ĈQ"�� �w��1����ҧ�c��F���1�+��|'����� 4ɵ>!�M�_��X�Ԁ�+� ���6}`%k��t�{@u��Y]<-�"��~�-�ʊ�x��r<��g��~���7�g�6;�\�vI�h�&��m�/Hp9t|5M��q��F1b�`P����э~�o��4pA�kc���0��0	�?p���m�����!o�m����ޣ�~�s�eR�w4h�N�ʺ|L8�+�9�x���f<캩Q�)��]b����q�Y����:z�}mYc\��w�/����+��� �Z��׎>�)�����_U0�0]�?��U|}#m�a56`���b�"(9�P
cj�cЏ�8�rD-�FO6�H����z/�҆�;�{�Hz�VG���3��ضtO��5}	Wf�������(L]���T���R����wR�Bu�H6o�~��PƎ�QJg�z�n9rg*M�k����I�0)O(�?�k�9�ᾛT�I��s-������g��9�O���g+�w��ǫ���KA�x|Ԑ2x�%N�")!�*���}�D�|�8{%��IȭJ���V6g�W6/�����_F�K�����sPo��L����L�F�1�+�`� 9��o�-��R�O��5��N�UPZ�
8���WB���4I��˞��{��+����q:�Ti����D�)����G�`�th��)�S	1�=T�&F�\tL��w<^P���y��K;�10p����ɏ}��cs�b�j��~��@"&t�m(�F��i���_�G[l�e���#� ��Ζݶ�6궙i37����1Q����u�M�E���nb�|�Q�u�8�)g)���dDn��K�d�$�wқ��ę%�l�d�w�����L�;��fV͛�?�.@j@8��l*yd�;^!��&0i�z\��>� �|y��sJ>f�g�ɀ��BgV(�����㮔9x��
�O�_�j&B@ܠ�h5�%zb#�G��~����h�E�J]�@U��Dm�o���a��=w��o�n�����ޛ�Ae��� E3 �>����b	�誅�
��ځ3[��1�f��X׈�!K�5)�yV����T�v�sO302
$uǝLJ��?�:RSZ��B���� 1�֓U��	�ӂ]�-�H^jA�G����o�3�U.�a8 "tS���'Ù�I
*[ƛNv�p}q�Tt���<[Xy<[�>�(�~ׄ��u@�Q��:��{̊jq��B]�R����^�q/�.�#U��+��J�{��5T�7K�]d,�Hv��r���� �V�)��8�����(�xLk/;?�0�>�1q�A���#�\8�nrjN�-"��C�0Q	�9�p(9F�<u��c=�Iy�Ӂ�eHcFJ��c-�2هԛw�	Qɂ���Bt�Љ�Ë~����ji�������^��w�����)�c���1����9�
��G����`q�[�=���C��K[�އg����K�/���{�<lmo=�;j�~�8�z��s�Mp������^�n���{5:��_��p�����j�Z�)�򋟇o��*���o��cbd�p�eećAwqҙ�!���V�p�p��\q��)�C��%{�I: �y�JTl�����z!d��S-ȶ��nYt9�ucT�N~��! �b�$9b�<8VU^��|�p����A)��K�ʐq�tT��"<QaA�$2cM���x��d��x!R�7����m��V��' t��~S���S�>�c�tf)G)��Ҭ��^湢�����\�9�˰�"ۯS2߷�������ޞ�;<�5��:`�CX�Qy��5��P"����������ﵝV�on��<U!=��hh�Q�5��V'���I.;i�sFi��'+��|�b�>+�^��,�+<���g�`f�7�)H�f@��@9��FB���y&)>G���h����G$}�Q��2ïk��Y�;�7�ѽk�n2C��=w��?v
���$<x�	�v<���.����[�ί��o�Y�L�j ���M�h>��>����a���h�h�+sR�	dEm{�e�(=C�����d.��	H��Cđ�I� �q����f�}X����<��{��?`�esF�(!s�:�M������ ��r�[>���k2��O�6�>Sz'�N!��0��
a�@���,3�왢�Rܡ��Έ�F2���CQ!g�6qS��c�3��a܂��[D����g�>{���Mp��xW�p��x��3�pW�����bq�1�k�fQ��U��������|��O�f#������j\s�]G�q��]����]7�M� <�}�v�f1N8W�:g���FITȀI���\lڥ�O`�ҁ<`I�v	;\\̳!L^�>1���h �&��*F4
j��]� �CFH*UP��8�Y�B�:q� ��wkQǎ/J^�L}:|��T����]N�7�ܞ���+Zў�ލǋw$E���ʇ2~,`'�3<�����K���;y�d�Z�$�6d,s��p�g��Ѐ
j9�r�f'c��s��^U�4�5�:π��~R)xt٩�g�.@s>��TG2���lp������N{b��lދթH����:b���KFB�'K���� �.�m1�����W� �qK{o�m�XH� +鳇�!����O�?���
����NÅj�� �z3z�7���<����Kp��m�5����_�������	k�I�DB��An�g;�����Qyn���g������%�7�z]�Z��\UerM�ާz���P�1�q�{��I;9K�P�1��%�6�?��F���M�GE9hF��&]�������Z��8SԠ
GZ���$��v�=쓐#��&I���UG}�6F���F:����| +�$x0D8��q�<'|���]��9�W-ThE��?����J�rd}Q�Q��D��(�ݘ��h98dq<�&ʵNi�s$�K����-�^��)=J:�� �c���ʯ�p���sL�a�d��iq�����A���̈́$J)�@�������)8��Y�*�����CMK �D	�v��^^��O�x�W�ڀ����zm���Б
��C~�2���w��ϝ�~����������c�܎_�1�P4��@�f�c9D\7�`#^�!��GKk��w.\����o����a��:Q;�mi���V֎�е��
{�uF9�%����ZTֽR^�EaY����V�k�4�ns�м8�]d��ų��Āz�����(��=��5��޹�6*�׿����R�|rN 9G� 5�����q�u�>]# �_#@UK��h�!\p0���.���vJ���Q��S�_y�<v�p��&4�}���T�&��96��6�MĻ����l8Þ���N���ma��~����������n�Xt�PgU����{5WeJư��]]#։ͮ�Q.�w]�=�F(���9}NG����尒8�I��9Y� |Zk!7�N�P�s9.bo+ �wc��
���.V��Z@���]��c�Τ5���$JK��<�F΂W>�B�����X� ��jG"��Ma\Mlu�-^It��kE�������AG>�C#-xIF'sdH����e��b�4�ē��y�t�C��؁�_Z@oTx�5�"��u�G�L�_,;r��$�<^�ę���~q��z�����컼��5��^ �
a�#��b^$A69��'7^��i^�/�ɒ1�	F�R�����H���o�Q"k*L�A�ߡ���n69���q�?���q�IR`�ƨ�f:�3�1��=����x���5l0�Z-��דv���sk�����<=��{�~����~�G�?�ʗ��kO��Cd<�� {�8���ӭ#v|�;�˟<�����+h*�NǚZ ^���LeK�$G'�'H6��)=":�I!&~&#��GүJ�`�	�B��zY*�h>v�*%�KM�k�w���I��H�@s�~o�<,����lP��9�RG�t� m����E��Se#�}�lEC�Y�=9`��=���cQ���֪�s�%!��~����Ȳ�ޱ�i��Y�U����j�d~�c��G˼Ʋ\�.w��;��-�X�v6�:Ē\�N�l6��	D��*m���mD���k���m�w�ήq���gTlC�o��iR/`�$�]Nuc�Z^�t�;��z.;��,���yS7�ID�I9-&�z,^�h�&FuN0����o֩�q��Zu4-lװ�3��!�}�������Cp�m��Z5�5�Q���右�a��	�J&y�&4����q#:e�ְQNy�t�P���Mx�ŗ�^�b���.P�\S�1��y�]eVQ�o�c��.r����r�w�cޯ�����{+�5]�e�y#p0in�-�⏦�U��l�!&}:~�J>�u(z�[�N��4��z8)o��c"�7s�1j�>	�7�}�u�*�ϱ���B�'|	���aAgq�I�I"'H��"��T��1��9W�|�/��Q3N��Q6�ݥA�L��w�0�c82Ã'��_����s�<�~��mC8���g��]w��k��F�d���Z�n��[ǂ��
1�|i�O���7~ί����~Y��F�^�ae�I���^�nҾ �w���J���d���}1+���^V`	�L��F���~�}��A�x62�>DC#m�T�z.�t�jLW}D��>��5����ʹע�q�	���^U����3�cŋ$ ����e�����/187)�=��SV±:l$�m@<�yA���Kڶ�T�j�/u%W	0���e���2W,�G�f77����������2&F%��d���&t]���$%���3Nd
.�1S���KO����%�6Aީ%��f4PT ���b����W\@��V���G����`�Y�MXX��Q�$����Ѧ�Hz����;�qC!��6jA5�3o�M�h}����]�Y��������[��A)�Ωߓ˥��V��k�J� >+G�if�cDw���W��4Ѹ/N������u�٩2�q	����$/�3�Ǹu8����z ��W��_wM{kr��4�M`��P�n�������?���~�G��i;s���,�6o�ih�7�H� \�b���q޻8��ݿ�>8����ش� �:*�	��x��;���/���.D���KCE!G�ث��.J7��������K"AlpŃ���	%>f�=y���w8��?G/���q7�T��/Jl�y��K�=\�mI�A���*'�U�k��$���
{6��&�a��D37�wKM|���`�~�����1�������
��bj�!�=��P�0n��N��f�}Ȁ����N{��� �1f'�@���1M�
��tg����)]Z��'�ۼ�X${d_�kћ:����E9-�P>����&�V�d���y��P�i�̚h������8��* $s ��:\���VV%r��E���c��x$���Mm?�_8��&q�_��ૄ�����&7���q��t�Dr�4!�s �ۅ5�<���ʥN�i8�
�q/�@��x���&F0Ge�M�!A{~|�F����a[<��U��ܴ���4���w��&��O=O>t�yõ����}f;֭�<b���ⴡ#���a/ThC���P�6%V�xس������-�맟���L�p�x�:���Y_N�M�H��׉�k0Y�E��-�|O�g���5�J�'N=S(�n)_[\d�&g��ʃH�	N�lu�h�>�7G$��#pT�'~SaE���q[�0 �������P�r�ɓ��4ah�T�#MS�#�C͔k��0��d6�:-�sv�@�P��h�!�ڜG�o�a
��i��[��/>q|����;n��7�	^��H���G�1<UȒ'�Zb��F�p80>�D9��a5��������}~��o�o|�{p�@5�0#�P���@�ѹѠ�'<1��@�&>=]�&q��."K���*VX�C6P0���3q?���r��"G�N/�7P�w_�ŷ9󚤚d�
��DL���p�k�z\���������>�<*�(
����9�h#)%�_Q|��^�Dz����YI^�5����EQ�.�j�$��� :5�J �W�.��4���x쌠X+:l����g�=��,h~�_��Wz�EpF���YM�ĉ�9��ZG�3Y%�(��{��]��R�N��.P����{B�-<�E����@�@}S��4��<רG�yIG�:��tޞ����������gN��'���$[j���
���ae�x�Sd��t�P��:O���R_s��矌���(*����/�V����������Kx��w`k��1�Vjh#:�.?{ya	C�Ђd��Q�'^~mlT�3��O^{^���1����߅_|��Vk���jP[iX��5y�nx䶛�믾��ap4�\t�.����|%wP�ne�#����_�A�4�ޡ蒔�`V�4c��Nʀ�9:zS^p����K�Nb��21�LRo�^Bz0ʁ��8.cPn�8!8w�b���Ġ�Ie0�K �AYN���`��sz�]k-�e�>���+�ض��J�a�R��I�+:�S���:�����w���M���Km��c��\�sS����u3%`��u������&m�n���Tp�E�Bя��s��$o���p�o�\�l���dve"�Nm��}ߊdd"��[�滊8p^ӏ�x�.!�Rg$κ�[�h�Q>�e��U���Gz�c��1���)�"il��#\	w�`�z��� |�5���Lp�P:�C�+�o�p ]��l��[]F;p|}>q����z�>������f��x��ڟ���a���M�;�]^��f�(:�vj:*��?��&�@1��s��^z~�Ͼ	�����ґMbTR�r�����L��;�c�'䖴��tbѬ�}���t3�e�<���S���ݒ/�����0��x�Y�p�%}F�ˁ��)�F�֌\:�V���ș�P2��[�	�A�v�6�|�J;��bF&y��J�@��#b�H��2i�1���k�N�ק�;�Z,`Gc8��~� ����>�0<|�p��{�1V���7�ą�&D�{d���L^���%�,{ 6(����[���o�<�}��+���~�`#��#�B��]<���|�P�I5�4= ���+�e����L�&�t2��ǣ1�z?�������览Ѻ�L�O#$&��<�I@�#�����k�Y��;�k� &��xAc?A�6u$�y�(^H n�M��m�ID���Y-��IYb�+�/L��q�D!�{���Sn`�#�|7�ZN[�h�t�p���NSQ
&��ƅ��ᔂ:O:@�� �/�w���c�37�t��c(�$-���]�bw���7G/R�&u%� ��e����+��4	㤨no(�t>yQ0�����27'j��8}������2�0��b���/�G��:����6^��vC��x��Ƣ��.�b>I�7��pjz����l��[�����lĝ��Ql҃�0gqͲ�C�~�������������(�c�ex�6��Fr� �82�Z��P�a4���f�	��_��o���_y�10�����b��:ڂ|����/�ުFU��g=�t]�u�Sw8(��?�W��� ��~M9�3r�Q];�Q��0 ����ttK:R�Z�K�YI�̾7��+I$�Oq�P.,ql�����n��B�.�X''fJ��^8�F������k}#�����ح��N��Q�s��C��@d��6N���ɉ��] �@�u����]�Y��Km������Wg����8�]�}4'�f��7!�=��#y���cȑ��7s�hօ��|�2ġ<	��!B������o��V��PVd��;��9��^��.ϥ�[f���J�����L��Y���1y�<G��an��R
CV�T~Q(��$-k8�3D������Q�\���&�}!lzE;�7J�c�y} �~;|�੏��{o��M܀�ՄQ<�>D�	u�Q�R��`QF���a<!�a��Q=���n�y�������|���ނ��߂z}�M��k6(���w�����#���z8��wx���S���]�@iԳ�Fw}F�I����rސ��d�3���*�b�+12�A"^��v���9pd�שj�EC��4��H8�5�^,���Ǥ.K��C,�T@��{�����	��'M�L6i��OVN�ed�OK��4r����_k����g~����������� ��7�_|���S���;�u��?Km<j��h�9�O���f��i�J���� t� duA��_��>��~���?�|������c�P���-��"�2D,���0�ԟ�h�G9����k�y�R����Sy��/Q�tn:�9�mj+�����d�Piש85>�t��
Q�ҺS3��Jv/^�\]�3�m�Õ�wM9�S���c��K��aر�aC%
E%����%N=j������gx�v�����>�O*[ʳ@������Z��Kj��g	�k�g������`P,�Q�&/h�օ[r�;ޠg���~��XrRg�oS���,�M��J�-w4��V䩃g�U3�yR�����,d
2?�q^��?��=�5�@R��w��Ah�����a~ ��P������Y��'�#HלtH��w�U\�P%�JF/��(��R��3h���o��7v�}I]a0 ������������ֆ`U\1����#�H.�0�T���`�7*�D��������ÿ�M�~�8|��{B@ðt��CڽU���p,ߧ���	}䍥u�Ld����)$��q��ķ:[G�E���^��n�?�I1���t=|�JG�tx �eӂ�2kw\�:�^���7�P��">���&��-��ұ�G�:���9��7�W�I�)�|���@��@&����<`=���݈������q�iaL��S��k��t�m1��z����0�m��۳'�wz�UAd�a��7`�M��pF�j�\�����n3i�"'���>��E8�7�	�{�K�a�0 K�[�Dґ{o�Pϻ�+盺
��(��y��+_Ӽ�?�:k0)�����mИb��Q��R���t�������,�I.�g�M:�w~���ݡÅ���Z��3n�]ڂ��,<~��W�x���)��ƛ��7���6��6� �]�H1��69�i�f�k�ۦ5�zu|x5��<^�4���~ ���g�G~g���67�����G��<й��Kc1*��k�T�t�$�&Z�K{HGF����)_~�I�����:
����lyLoƔۈ{�	;��1��
�����ns��k�I�G0dZw�y�D��W�	�䡥�Tr�Iz�lbH*O��a�d�p�T2�,DPMw>�/��@&�/��Lj7�12�����9̡��������Q�{z�5*�w��[@1�	��[n��|�c�? �|NYk��nC�/�������8���l�d5&�K�H-G��"�Y���4�{��v��=Ͽ�|�����/�^?wFk_��7�?=�-N��,d��VԠ��D_���{���[R���H�X���$o�Z��$���t��S�4�� F>�����'�#H=��J�J?4Z[�8W��q��hע3�f�4�n��@8�L,���Cx�A�X�m4]Z<И���$�(�#��q WJ��^y�P����3[,5�s�޴y�ST7��~��~8+9�W	Y��yy���E��$gH�?W����dTｘh:�h�e��e�w��rl�ӈ\f��M�/�y ��&Nl���f>�ɿZ9�ѣp�GSL4��(kW����w�o
��`nriZ�U޻c�����N�/�f�����S.&��/��ޟ�鿅I��!�:_$zS�Zq�hj9�*��骮kXLh�A}���]��Ro(;�»�����|�'�[��F'�Ae�ûmk3@�Dk$�� 	JT���י*ۄ���Ǉu;����u��������o��w�:n�X���������ƛ�����ó��������,�b�>��P:A�mzQI�J� M����|7uN�<��.�hc*�-��UǪLg��^��t}7�<��되ϕzGvҳ��OGc}�0�J�8�;�{&�H��x���30�q�ţ�XG�w��op�����>�T�a� ����\_g2Ik�&�CtiZy!�+�����ЧVtxh�Ma�{��j�Mj	�H"���!�%�?�|����x{��H�YBh ���ӼB����I$�8���Gs̃@������Y�e�A��&���$�&��B�E)�_?g���h����>�[&�{������G]2��'�#����SX*;�rQ4<���5�xL��0ju���ym>q�]�O>
O�{;�}�1�\����35�o��������|B-|44ܐB����bC����e�C:b�4���1\oÛ�?|���矃�����nu���Ga��9F`��I6�1Xs�#<sۊ�UwD�͈K����_��Oz��]��t����'G������Hᒪ��X���y��6<�yMW��G��k��"�23$���b�0&�����ѷ����j���]��t����.�R�]���9���-1�Sxd�����ܟ4����M�"=�3��@�����CT��B�'9ǋ9X��������a0u�o\�� y};~O�||�4<�q��曃ӆm�v; ���
�g��'%��?e�L��lgqffP����y92�iW-(��!<���}���k��W_�W�o�����`�p؂� 4�X]�<,��`�P�Y�*4��[��+�N�Ue6fc�pE�4�Ǫ��dR����Ʀ؇si�1���8�g��ԑm�z����i-�ߕd��qS/^�<�E@��������A�k�3Vސ�L�8���.�a������C*�������ɓ{�|����h���;Z��d>�E�&�r�k����.F��dq(�&��%�8v$<o��睎1\�*�n�ǚ���^�i:�r~ԜF��܈��_]RU�Is��_�#o��ɀ��>ɛ�@�O4���!����)��r�.�AW��).�vId
V�	;P�G�p�-7@�AVxs~4���'��G��ς�l�u����1���7�RJ���щ*��#B�m�PP��񼂁k����6�O_}��{^�/=�(��Y�i�����<
��||����2Ն�sg$�p�I�1��T�O��<K�Kڮ��rS_�)�)�Ԗ��=��ё��S����`.Z�SVN��}��f{�ǆsxl��2��/6�ǽ�yE^��qVO�Z���>P���z�V�7����B�X��{���սIFpJsQ^Z�
+:�t�󨯻�Ʒ-�w���Eh>��O�-�O�u�c��r-��y���U�H�%�^��#��CV\EI�^��N&��ӶT8d,ٷF#?K��g��>S�ג�1f����k�|���1�����)C0@v���x�#}��#�`ˆ�(8&�������-�o�0a�c݌��p�������'z��:��v��iܖjp�#��`!��n@ux�b�����D�6�Uذ`u�@��0ּ�`{�?}�mx��Vy�Ux��W�ݑ�����A�c�(p����<G�X`�?�iuT7�\W2��c;Y��z�zK�R([^�¶ʡ#�S�f=H1�Vύ��*FR�t^�R�C@.�'a�YiY�\NB���<��f	~
�_�>5������Z =dYywK��(L:�H�	TzFv�FK��]�7;Ns�=B�Q�Z.�jR!`A	$8Cs��tr�d���	��'EB�2Q�.==-�>����`/98�N�w�p=�£��K�?��666P�B��Q �	Q6���\4�9B
�<��x��<�_��g�N2Ǳ�+��U*���wv�7߆������2���Gp�㕍!���h(�h����*$C�%M<��"���V���0�v}&XDRCu��@�c�&w6r��T0�sUgCS{���H�Ӹ�p�� 1�B7�p�N�n��~/"�����rV*R^-�����4�)��قJ�i:Uq?>5(�u'N
�󺙎��A�,�_`r^O���a�+:�����yӛY��+�O��v�c���ӝ.��,ʣSj�=d��d���� 0��G���̔F�R\��0��FBQ%r�هTh~WP^	�W��ct;5�3G2zA4#%�V�p������b.V��)JY�r�8̯A�k@�E�b����N��#�p����1#6˓�%�r~t~���������p���ƈiC�T�o>�1�:h84�p�H�8�n�ʡ5D l`��n��8����կ�>v
��*�5,P�?Wmy*x���g�e�� 3�%�����A�? �ɽ�O��.�u�|��#N?�bv�J�eeM��p%>�&�ض�j�q\��Hu`��Jᗰ���q�����k%�Aj��C���۹�����xv��u��@�`���e�
+�cE�h7�q����>���d���m��p�l�AW���Pr�;h�rbO4=�[l�8+�d��ʲ�I�k�$sHM��������> �li�h���'�1}vuƲ���U��bW΂pLV?�w�,�!�;���soH�A�)#Q)^�����Dwi��q3�Sw����������|#�����G��UH{��+�&OZ�8�47t��Q6�%�z�7�ZBؖ�J�����[��W^����������:w����X�f�d�Њ�^sx4��M�&�>� �*t�����Z��X$��H�].t��~�p,�����m�e��E�����?�f"��,��̛���m���h�Nf�+]ŹC�5Kc�� ����d�L6��%7���K@M���<{Q'�JHM��f�хF�͒	�c�Җ-ɓ��/Y��!&;=��3��x;͂'����V�*���``�3����<y��O=��/�y��plml]��f��Z"i���8U�����C\5k�Z���L4NFg��A�6��Ν�Ͽ�.��3?������������#��i(ʇ7� .��&�%ј��*>C��Hq��@�Řb���-)	j� ��o��f��X@�Z�KP��A,>O�OIC�OZ�tx_-�.�	�T;�wi�;Y���P�z$A1�����T�Gh% y �+)� �䙂R�1b(�Y�0^ъVt�i�\�g,�dC�}Y�u�NW�*�fzʠ�}��)�ȭ���s-8_�ݼ� ��er�WL��D�e�|>��:uwC�`��8�d��NPY�ĩ�%x�%8��\'J���f#��zL4��Eՠ4��ӎ�Q7��T��)EJȌjx��{����w-�]��Q��n��ww.���Pq��|��Sb��&D�F>�#����hh�\t��YX��X<(:�7>����/���u�x�ۤ!A�	�[�l��r�񨽶!��N7TlX2J�$-��N�^�ʲ0���L�L���=6���y,Q�:2ڤ�9��2�
�k�C��_=ԙcv�͵��Te�OB��a��N�O�� @�}9:n�8s����H�ɳ�\'�E_��E+ZѕA%yQx
�At�\�ߜ`����)�'�����䟔Y��N�n���H�Y�p�G����԰"P�����Q��X��kn�mє��!^�!ME��1��y�(�̛<�{d�l��J�蜮�`�4��kFCQ�ǣ�յ���7��0��-kk���'��{�[�;a#��N����g��H\ni8�y����.媱��5��_8�;D:oVq����9x��7����}x����s�a��ԪJ��X����ӭT�s:�%n��am�9Bl���ֶW8�N�xQ�H����o�甬� c�NC*���a%�=$,Kv-WteP�,�	����)K:Bũ�.�r�`��x�2��N�UHiB(^��Đ�'��fR�ӥ�jcZg�TW!�M�&�%�g@��MÆ5@�_0󣇧Ln�L^N�S���fw��#ص3�!|��;���O=t?<p�68�~���Q���W���=3�O@�EwOZR$�������+�d���Z9|��E��0|��W���"<��8�*}H���C-��Th��F����%C(F�`�'!uu_Qy�	�����d}���}+<�RS����a����S�G�pyыU!�R@�{�/OD��y�2V�0ԍ oM"��yb��ctVڝ�p-)Ѥ�t�3UJM�C���֭������ce�\ъ�F��Oj*�A�֯���{���,=P�X���"���N$m+uM�yZ��r�� E�\����C8W���uԁ䷞�b�*Ν��xN_3�k�l6��p�+�#5����t�����&�8a�l/���|1�(����Uψ6)��NE.dG������h�/N\��u�G�.��Z��/��ȥ-��1����������t�Uk���0�jMr�pbz$Ӊ/J��7�w��p��??~�ux���1|�?��I,J�L9y�M��b�� �ȕ*��������w܆i7D}0ū�ҩh���?ȱ9�[��D���9�9�Hڢ��I͌ҕ�c���ĵXo��E;�$&��m���f���("9��H�۰=���|{W�"R���w�Δ<'󘃎���<M�s9̾_ъV�g��)�LW��bz*�@�������)��.F|O�O����9zVۚ�|�Ͼ�8��ф��~& ��N캜h��r�`��kZ٤f$�b	ḽ����7�֔�i�ON�ȳ���DY�.�>���U���q�Ё�0T���j��N�}��l�����ۏ��N���.x����o�M��_�	X�	
��qH��ڒ��mF�֎��-�C::��щV5�	k+0�E�O�|?|�5���_�o=�:�v�\h���AfX�Ǵסl�(�=�#Dt���w{$'6�'�j��ӣ���K]���ٔz��ԵcK梣$�7)�${a��ʜ�8z�7A]�2pB�ϗ�.�k�m��*Xs�����zV���"�:aҹ������^'��w�"ey>�{�/�Ǵ��މ�$Iä/�k�5N^ȏ��4r�@�eG;7���&x�0�z���#��=w�g~ ?� �}�T��<BL
X�'k�H۴���K��	[���7keF��Q��p����q���z~����^����<|��w�l��=���z�7�G�c�^���Cǣ1�D Q��ܲX��(/���D]�s�~���lO�s��j�&:$I%��Y�j�&�,I�$�tkH��zj�2�ߤޣX�8oj����ѷ� t;;u�9)#gq�f|��[�_gd7�!�jD�����4��o��T;u�*�a��X��G���pЪ>��83r�a�a�}�N���O��s�����V�w4�ik��B;`&�<$S8�?6�'e��u���l�s$&��T�Q�u%;�6�I�" G0F	���sm��GY�2d暞�j+�L����Sf�%7k����Nؐ-���A�ј�I�C����-�:�m��R(l���:٨OCh4�'�..uĝ���?�Y�m��i��pus�
�q:��DL�5��w�p�8�85�X=4��Fc��ن�[z�m�	��b@�w���"�At�'g���."=���s6�N����ε���r����W98~d��ᣘ}¯��%hcN�Z��uk����{d�̅�pdz���E>�ߜV��l�q"��iIaNd�v�`>T�hc�n�F�y��aƀ���'�B�[!��U�7����ߣ]"F�����O��тE�l��D��/{_��p"��iCK�띞�a�u�I��"�����y ?Z%]��̊V����ʔf&�ƀ6��QIt��;;R��!�bcR�T�X�(GÂ�����-<��'�N�:�U�<�Zl�'��]�e�5�2	F��S�Yp�#`������I�s��E���%�y�*#�N���E_�~'�5�PD�|ժ �:ᜰ���A���Ȇ����M��a4�c�����'�>��> 7ۄ���yݿ�cK����0��/���i5���#q`�m$U�2��c�t��썚��<����-������w>�Kk��5��7nZ}gM�6�h�)i�'b8��Υ� D��������=U��>*�j�si>y�~���\V��H�,��*�ːaWJ!e͂�ֹ��Û�ʊy��;�[@��5�)�/��A�v�h㕨�A�B��+�J�i��)�V���s���(hJf�eЄN6}ה�G!/c ��n���fҐ1��ఒwM</��ѦP�Hׂ����֥�p��§O�_�����G�[o���L����>�u4�e��C�x�ώ��1h3ą����eß�f�=�l��b��Tl�.����=��k���3��@]`}�Thi��|ڃ��C0ި�G�!'�&^Z����0�B��3)0|������2A�w�r�s�ƃ���=�ɮSځ��MNu��sn��S9�rB/�\����گ�9~�,����$z�N^B�)*a�$���1h��N�w>����O*u6]��1)_N�e9����[.�Vt�I$<7��ǽ�3��"dY!%kf���"�3yNa��m3uzK�z��J��1{:Q�u��ΨY�+/5��p۹�Y�K�@S��r�����	4d�#G������aB�{*=��6fi$���;i���+1H�,�z������9壕F���EGp��%�Mcְ.���"�7��ⲩ*X�C���ĨՉ���@�����`��P�1ҟ�G7�@����@�Լ�bX�i��>�#[����wA߫Z��i��l�J�z�n�9>/��)/��*Tq�����l�X���}�-��IY/RLWN^W,D��D��%]��A���, I��]���e��y�dN㹰�F�n��[�Re]3��4��H��I���)=7�9��,��/��:�͊����Ė]�]�t��l�xY�3g]�ٴ$CR�Ե_�����Q	�p��� ��L1eO�
#s�y���FdvĴ(�,�s������� ��zC�R�Em���B����2c";���]�C~u�O_ӱ����wt�l(�&b���3x����ۀݷ[}bg�"�q|~����S�ă������-�߾�S�T!�qHǢs�_��z�WD=Ǜ����pR�5����u*SCc+8w�,|��W����}��O~
�n_��z�/6���M�~��M��.�x�)6���P�Ɂ�����E-�@:���S?�k�t�bv.��k�͉�ޥ)k:$��%��I�Pk=I1
�"�/'�݌6��ːY�MPCd*9�,�v}�.4�v�#x`Y;i�����IHvI#��Ҏ��M�����`a�#"B� O�L�<'��n:Y���!i����m�]xL
��1 o��C�����#����9	�=t�̃��]7�c��0��^H��4��q�d�̡+��NAX�H1�o�5�}����;q�g��^�h���������[/<����>�smY.�|�6PZt˸�2��JX���t6x���I��f?�0_�]A8(���:�𼼙wn�&�a2��;�o����U����@*��_�~g%*]R%���l��
��]r�ܲNH+��栉5�1�����X�]H����2���b~qı�.s�j'j��o����s�W���� �=-�����F~�9'��1M��>y�TMd��q�E���4�@.;�`EWM�7'ó>C�4�z/Y��[N�mU�!K�<uY��y�<AX,���%�9	��4?�c# ��P��&cl|��1q^:���T� �ٰ���w��VתLt�hȤ�����d7X\�H��>F\T:��1CEftI�1o�5v�y�lPŰ�������"æ+r�<+]R�K՞X�]�i�I��vҼ��+X�u�Tr�E���W��iM�Y#.�k);�'�߅rpҫ�'��c2a�mK)����h��>�/�v������Yz���>^8<2oB�Wt�S�9�Rx������"ˀ�4}/_0�v|FA3�ym��"�,�G��[PWT��aq��&��N � fHD���:S��bR�I��S���x;>Ӏ���TM�6��O�?���x��������w��O=���6���M�\[WW���3�i�U�@���e�݀T"�bhD�:Tx<��q�m��/O��N�[��3�K�_}�G���?ٺ ���w�Z;Ҫ@�*;��Qw��c�LXgA�f�bl��iT����MF7��7z/�d�� �=����#�I9*�lT�?�Ð��v��}�t���µϴ f��GW[�eQ�n�Y�"��㈮����:]�	q��!�>�<��墼S�3A_�w]�K�O	ʵO��&қtbWK�._�$@�c�M̏�R�V3w��mC:�~������Gp[���.��c��~���MX���:�������rT�b(s�,b�4�W)X��*C��օ�Ä>��7陳���ނo��&|����/�?��-��[�� ��F'��W�e�!,:p��hb'$_+}%��pyS��e]�<ϡ$
4���\'<!FKIA"s0[��*� ���ά���Ō������|S�f����Q>MS"�Gw'�/{r�2����!��76�n^W���d��Â�� ��q�h#4[�,��|w0�`	d���cE+��\���7��t3�iH�\4�^�f@��餴a3ID7գ��=���ny��O�gݎ�#c:l1v�7����g�Ӓ���L�y]���1�
fv���-3�[��*ggQN$C$�-JN9D�r#v_�7"�0��F�e8��-������]�|������G���h~�����Bc�0���h���ss��U�������z	�Z����xl+�"�������&�g�=��Q�!�g\7���\~���Q\<k�h��R´�O�QS�&t�"�S/�b�S�������Q�v����/e��*�}
�`t��RQ.���B�K,����Sc����8�9h�r��"� ���I����3�I��{Q~Y��P�~���Lx���'���±���,|�W����m�iL%/d�j=��9�+����$��{����2p٢�*E���vC�|g�z��wV��W��;x�@2�	O��C��;�[l�R��rGM���p|ܵ	�0<���}	6���=?�����'�G���\���f���m��4N���8 6�z��H�I�����LH	0q	��p<�{�?�g_�)|�W��^~^9w��1�9T�����m_q�^Ee��$Cy��1�,�'�)���<��!�T#4�t�=��LI�ANW�9�N.�ǀ�~2}̹��Z�d2��{���z�$���{e��/]�:h��:��C�m�z�Q�u���ŏPI��!�p�v�Q�B����AY�Ԋ��h!A�����q9���7��V�E���[�1�̝($�8����Dj�8��ã@U�t���En�	Kv�:4�Oj?I������v���4<~���_��w�n���#�vZ���v>��	��G��qq6�+��h
\�x/�����h�jA�����[o��}����^�������A�Cn���4��������iW\8&%0\�� ���肠F1��f��A�|W^g�M�3 Q����Ǩ��8�⟾wR^c�W`��	
A�}��y��BÖ�~9�7��M,K��H;tp����@b���q�\�+�S瞼�w��"��~�������~�nR�"�D��g��4���]")�GS�=������g��x�u����h�v�v��7����lL�3��e��yN�<#�RO?�U+�K-��K2�!r�dN��!����$/�l�2��4i��(��`+�����]�K#�y�!���p���Jؠ�+�kRШ��˼�}��t�D�)��.ּ�����xC�u�uOi�t�R��,�;���q!�������cΏ#C;�x��:�E�� u���z�|����hT���7��#G�kpM5�����j�1����&��j���ۑ�S����(U�}�jo�8z48������+v����:W��K;p��g�;�պC�Qe~5I��c��m�Y�)}�Q%=�$��c{����3����ܦ�_��*�${#�H�@���z~����a�K�d��ف:��a��h+BW�)���),9�Xͅ��2��1���u;dl����1ɦ5i�AR�V Y�>��G)-I����͐�4<և�V��yh�"s��^�>�cl_�	�Ҕ��g���+�v9�i���}��-^'g��dC�r�|��b}a7*=����ޣ��R�s��%SЇP�m���a	6���u͘�7`6���Y�Ɏ���.
��s��NJ�4��B��n ~L��q���p��u�<��)���{���.�����I���%��	�nǵ�b�Mn��G��`�F|C�>�_Eϑ�>ؐۻ��%x�����}���͗^�W>�����RW~Ӭ�A��6qM��Q+��`x4����~�?��z$xZIH�=�d�������T�i.)?(]Iۦ�~F�}�SΥv����A�mT	���,;��i��ԑ�{+�R}{��\�f3٧��g���2�k�(��u���?����w"�4�2[T�S����[{ڏ�8k�%Q*_ߜ�1td���)� ����zyW(-yBBl�Po��'Y=��B�95���9t��7�����v����]����w�x ~�S�����?
G|-��裸[?.�ڰ��qu��EC��`��QX�D'j�-d:66o��5~����v��s��k�������6�aFvc�޳�n�`hA�@"����>>W��q�#R��jObS������_���j��B��߉��0q��:����D��Sb�<��a7���_�=Q.�D��!8. '�h������lVN��^_n��t���x�`�c�)��Q���v�G��t���Hw��uquo��d�xg�遦��4���s�f�g�f=;}b:Пδ��tfb����:3M�|�4'�w�&���X�'������4߀2~R��B�)�v�i����T#`91ؤ��2ڤ����6i��e��ul�~�`|�d�5}:1d��Q5����ʖ`�KV)&7��#��K�\/����C�4��K1�F� ژ�q!�E2�]��vlև�ޥm��a}�F]�'.����c�ণk�ڥQ����]����;�&�E!j�� ���������k��$����~�r���6l��w,/�,�8���WLϽ���\w�3��c��&y���|�i����.yC�i���2�i�����t֐q����t�L�&O���3̼i���n��J7@�M���l��H�uzՎOn.-*��݉�U�$��N�f�U3�Ĩ%s�ixl��^��I��̸��i��W^}�`�6��Tѯ�t��C�)_�j��{��]h�xk��w8��&�o���KP�2�(mb4/�?�%P�S�s򡜧��h�`����y4J�#Py�Eu�9������h`>Km�i:�!�1~kR���5�������0�k�@��뮅_�����8�y��pݱM6�O��ٚ���E����(���brio�$Kk0�
Lk0>>y�Tۄr�mu��^?_�����߄�;g�5�������S���ÆY�X�t�NƊ.Ʈl����ǒ��À^?�ːR���%��Z��4�.ez!��{� I'����H��u�q+���P���Qվ4�KBr�WW��~g���;�<jnVQB�F�Kή�	/�!$����'�B8�AP�<����Pj8�݃M��U���0����TD{&'�����J��l�V��/i�$�6P�1)����v�n�����_~�	�����O��ê;��0�i�������b$�H�i�,��4�n�F� �������{���߀�=�<�����8o��D��nCH.�My���lī4��`�D������%�4	5�+7�&��R�k���J
O�Nʞ���,�&���>d�P��dEt��p,(���va���L���h�&�23����:l0��N�^)#�ɬ`/�2�^�y[g��,�=��[yWtœ�|�}��䲋���̙�D<������4���rN�t��
�mL��䖏�S���9M��V�&-�v袛wv��N0i_�熦xuQv$-��F��w�2DK
�z@4�9���<&�����2�4� Z���w C�I\���&:���Mpp����6\�G����&�u�Ywb��q�1��;o�z� �谶Q�j��;5�1J�a=��h��1
Q$7��a��zͱ���F`���U�m���1���dgq���H4IΕ�,�Ї7E{�&��8A�U9�dFVf9J�����'�j�MA���]i�O�>l:��zjh�"��:w���MIdDI�j�0=[&Nc�*N��g���\��ɼ_.��X`3ײpUV�ޛ��7�e�{EW'M�#��|6-�}�k��M��x:������[o�)�m��3|�a`��aղL6I�"`��B�U�W��Cs���TcJs�@�m��:���&��_'�$�l�R�Ԩ�a`�[Z�5���rX<���-������n����ዟxN�x���uX�q;;ٌ�����"�����`�u�����8���-n��P���\�W�~���+�x�?��ۖi���+�e��ѧ	:be;��fr�i�~[�"�t5��,�����L��N+���)��'g�2P��B�4j]�Pi�\y�i�K�r�Z�c�O遉�,�7IYd�v��;��2��Y��Ɠ�k ��z`��lx���;B�� ;�8��Q8YQWQ7�^���QoV��$P���<�lTޔ��ԟt����h ���2 �CbL�ce�ҥqj����ȝ6nO�l��vl�Ɨ~~����ןho����kL�YM0�q�T����m���!/^!��B�eL@H02����|�������=���?o�\ �y�:���0�����G��� &�cSa�X���0Ԧ���7�"�.XEJY noW�K���Q��[���ߕ��|�&ァQ@��c�(�g���o�H���rܐ;�\��54�\��I���P�NJݠՙ��B:z��oNHe�c3=�4���l*݊V��M��&��H��Y��;��=�\Uءgl�N+��4rl�Z~��LX<���c_�O����|4BL?�yC��dd�40��'��Ŧ]�q���^;׍D*�<ջ���0�>1�J4f�`x���
B���#Ó{_���8F�
u��E���78�h\��2G}Ʉw׫!<r������X������T�5t�'H�N��z��֡i��o������ҭ�#V���ۡ�����`�2sHf1�h3�G��Z���F�J�x�F��EW"S�Nx\���6�N(��ӼD��"*�>u��풴f�7�k'��ϓ�\�^�"J���O˟��X9r ��ξJ]���V��������x��8t����>zek6���)h;s ��ѫg.�ih��˻�<��S0��efI?�IԵ��$�%w�s@�����.���؈珴��6��/|����p͑at�nu���jck+�Bt�డΣ�#4�X�:@tԈ��U������k�����Yx����w��n��:� ��Q��]p͌C��hIhB�khB�k4Jg!5����E�d�@�A���0�^�g��
�w�%����X·0��/�:w�:���p��T�1�d�y(�(�B��}X����q%�C��"2/�;���s�0�8�aw�>�$;���J!�>စ�J�,
k�n��d�E��$R/P��{ �a���m%�����3�e
\7�d��1������颟�w��k0[;��n���o�Mx��0���ѥ�%Ec+��+FZ��4�a�C;�g��b�]�������m�8�#����}�S�K?}���K�{O���; �x��0�MЖч�
�Bl�00$Oo�x�N�4���fa����kM2�	�:���J�������{-{8�^�,�W��d�25�$ ����#bdi;�C+\�V�}�E�ᨯ|*��.�Y�-���+Jǻ�t�n��Hq���)��%�>�)ޙYOy������V����H<�}�+�r'�֛���y��|h�y��aQ]�?�HK�U��tݲp)�X	�%�^��U:1�ͣ�t.S=���`M���?��eF��ӥTd���!�҃��T��F�#7�9�����M�P�G�����t^�� n�����%�nX�Vp��6�>{N=��cu,��u�V'�Խ�¦}.��j�ϝ�9�M����C&p�u�sѡ?~��6��<|ǽp�ջ\��V�\�~�����7z�?<���#�e�(M�\EeIww��x_�C���m��4@�����(t4�tMO�NcR�K����JU�/�ǲ���J��W��^'���AF�2{/m'�͝;O��(���B$3�M3\+۟�bj�t�	�&��hE���~uu��SV���6��7�p��`.��~����>I�+�?{�%�����J��pYu@��9U�ݙ�*��$�O�[&�/	02�w(��gz�_�h�k�z���6�k�ғ�����2�y�8��6F=G�N����B�46�"�;Y��X�p-E:���u�2���`.^�p	~���g�=�����/¹�����ذ�4
K6�]�kE�(�Ձ��)�]�Q�����m��71cƊ���o}/����\��^$��_%;����o-�ȡ�5jĐ��T8TU�Q��¦�逶�\<�zi?�ܴ�M��fzEk������Bz-<} �j�qڳG�H} ����.�S %�X��&�PI�?h��x�P��Y�'*���P��`�v�$���V��_�<4]�ɴj#���J��H�{JV��l$�d��8�~��z���n���W��[nj��C��v,�#�Аi8��P�D�Eo�p���G0�����{�ܖ]�ak�s��ʼ)�N�3�BR,")�P2e���,*�bH�eHV'� 0$���G	`�IdH�b˔lQT�D�M�g���7�|�޳svYm�}�=�~�k�5�{�9���k���<*;��߹O��,|����?�<�<��9�m��NT�Qmx~+��,����2�$h �c�����xB�@MV��'��E����,��4����ԵŎ)��"����#Æ V� � �shLµb]�(���04W�Ce��p�5՞���t�K���\�h|Z�9Ϩ����<�4�Z�d�w�c�iT��͛�
|�	�O�/pH�{6�L��s0�zƦ
?�!8�1迲y��F�@1 ���B�y�䁣dh��3:���4�s��t���[�r�M�1~�L��mb<J=�*	�ǳ�5ܿ��~i,�KS�'PY��BBe/0f��S6&ge�(�C<g8�D�Oq��!$ǚ�Χy�
�ʠN>`����[���f��3�S|��S�({GhR��a�o�~6������=���ـ���������@��݂��AĤ�r�g���!����-�^7�ބ�/�e��Y˧3�@|o�x�� T�ty0�� �vw��)�g3_1f���o�&6bJg�bE9e��u�Tk��+g�L&���!�i���]�G���Z.��HT	H���Cc�0-��	����B�>�M 9���T�y	�ʐv:�Z9������\������1k߻����q'[�l�G�4}K�<�����Q9<wA؀ҍ�*�w,m\Y��e#�2�\�ب�č��%5(S����;����F�����(�rL��Oߥ�TbK'e\6JF�r�W��M�~��l�u�>ZSZ]�	�𣃘yK2�~o�i]�2����)�;�GJ��g�����b�e��Jb\����%��rlT@�QLX<�!�_���L+�����/�\��	f'
�P�� 7���� M4ڠ�1?��x�]��(w����Wy1i�^�py�y����������y����VN��vf����;��f�8�B��Mp7P���:*˩J�����n$����^�MU��Y!6�+Ģ�����?����)a�OB����;�Y����?���ByJ:�n�Եv%��൑�]4����r.v�S�{!:d3��2�@��-��ټ�2�&��S	�Y��:�Wg5����s��Pi��I#w!4;�~x�FB,F�p��	�v�������_�h�A�cl!�ih��8Y.<Ȋ����l�u��F����|����O��=��G���ʓuX35�ox�(Ե���"Σ�p�v-�b�O�Cf�"HL�i�B�]Xh��Jf��T���ۂ`V=������T�����ও:y�|�<�$��(�'��*�.�%��1���Dq��_U�G�*7U2��W�R<J��mN�F�g�^��0���H�i���85��H#�4RF�2Hʜ|"j�ܧ��+e����OM�{[��C�ǃ�>��1���2����yo4B��x&�¸)�2��=�E�.�!�Ӥ�
g�ي;6z��B<���gp�	� ������֜o����mcz.�*���QZ��=������ވc���v���U�;��_����:q���n�o~�m����������ǵ4���>��5��c��Um^zǝPن���������>�>���S�J�C�VF
AE�+=�h�,?o�1�_,[c?�s���͈a@߉a�+|w\tTD���y��C��K�h�������Z��'�\]�����(��4�H+����\�j���Gݡ���q�O�)�q�#��SֿI��H��Jwvp����2��5�������1�͞#f����{(*=�Y�5����HC�[NzF��ăv1�ݶ���r�]W_��O}�^��/ހ 
XY�{4��a\$� �x�%S���;y,>������-x楗�s��.����_�18k�`Z��F�G&n�Md�e�X.��OM��!�-�tɩЀ���%��}i&��t?U��RP�+u�S�޵o�<b�{��~`�T������äD�:
�''7hp���EFw�x݋aYi�?F�ı�����R.��F5��a�?NlM3�"6�h'1#e:UЙ�aw��,�4���cJ]�?�Ӛt���k	d�C�@���w�<�<g���I�$���3�7�B<�a��D��p��u����1����H�G��nh�Aުض(�kV��Z��{S��yma{gz����߂���}x������:4�54-`X���x��+A����W��2,P�\Ö�Q��>��B.���	�t)�MT������$�3��2��:6�$:�ȿ��3�#/(�����-�t�Me}G��0H[��cM5�/�~� ���2|��Dw��D�G�E�\����V�C\�n��F�!��@򓻉���{{r���X���,ߞ
�l�.	���H���dQ�����fv�%����Xi��Vw��e�Pb�ryc�*A��k���2Ķ�9L䔔N�pjm��4�^8����0�u0�������g��xj�4v�N�N`�jN���b�X�a����Ji?������=�Ҭ�z��̡����c�J�%u݊��l8�o�r�v��p�uo��nF�HY�D�}�ū��c/������3"M75JҎȟ)<�A�,t�:��-v�$$JO�d�B���1����e��T�O����'�Iy��׹����O�(��W�#�4�eL�n����1��8��7�ӓ��4W�}��p0%c���:fF�CE��`�-yL9�<�goX�m��B�]�^Tމg9�?��2���Y�q��μ� �fw�|�pթ` Ѹ���q��h��6���U�^�,�x5��f�t0��� ����?��߄/?�(�pq�7& ���rۈ�}�WmT��o\ڕ/��sq�3��Ubb}�	`��:�  �Tҽe�a���|W�;�&��\˱x����^�����	�H��^e�+ĕ� �c������SF�;tㅽ�^7�F�[K�2-}�
�@<���v/נ��m=�m8�JV����p�[�i��#������E{Ж��}ՠ�yBP�Ya��	�vM����'�:�.��0�
�CĆ!W\�c����r��q-B�voZ ��/��y�����=�>��v��7ڨϜ��q�dx�\pQ�&x�΍�b���5/�XD�ؖr��eUb�?���|7TZ����Q�������2CP�a�F"�`�!:c:w)R%F]~��C)��;D�!ž��iC&�ʰ`đ�8�Ĵ�-lV��`_6��P:�H#]^��n S!��R��Ä.�TS�L=��3�Ѣ�+J�ko1��uZ�e�e#�H����x�0s%�� �wi��vff:56nAg��lRUp�-o�����t��xy�&�Z���V\�<�vW���h;����v�]o���o0��kk�hy�뎛`{6m�9�ީ?ވ���}���o����Sm�6�P�V��f�Sm�c;|�D/ �3H[����;���Ia�8��� �=�ʫ�̅`�O����s�=+C���ځ�J��͌�;����0�}|����X��ŗQ7�O^a?	���������"��:�7�����&{v��\�ϛ���;Nh��)#�4�P*�'��7��i=*�w�ɧr��3VV����Cp������0�8����=|:��4m��;v7������(a^�ɣ����O:�7��N���S-ގ�	�����Ou�r�n���o��vyMw |�i�������><�ҫ�Թ�pq֦rbՙ͐v�2C�A&&�3�K�5�T���J�S�x��o+=������%
d����NǠɁC'�vb̂l�Nw8�-����ɐ:�ÔҞ�+YE��$C��$���:���zM���4��l�-`X�60�P����r	��Sc�!�/�Dm4��Tq"�'ڲ����˲gh��Ӊ�t���n�<u<���(m`O3MV1�εeXj�=%e��lUǯ�.L%Ga����EH)�����x���6^�x�}�,\w���]^�x�6|��K���'^!�"1�隄{���l���x�����������k��l5��uX�l��^+a����2��g&�U>��.�b�b�+z"�.�ص��Rw逓Ŧ�ä�a����trRE$j�K�)�,�}��ey�$R $�6�]�/�C愣n��@$���
�u���~�˚�k2������^8�����[bđp�)�����v��Nм	i�@��F�xR�k�E㬞8�#_��-�C\O��7�N&	j����:��m���5 G{�V������l�X���d�h�O)������'b�� 5�gJ�,A��u��Y�ky1/��ъ%�bIc�M�\���6(N��ȋ��G+����+��[�:<����W���If2(��w>���ڼg���7	{���=��~��������V���'`�Fo��\.5q�!�/�geX��4A&oe��[�?������{eĎ���;pb�ǟ�󵅵�ê�D�o��]!hz!m/�.��SZ����ACBi=�S���R�b[�t��&��5rNM����z����0	u[ő�*%i�2>����8��X2��xTP��/SH˓��θ�p�߱��)&��b����yTz����#�4ҒD�W��:-����6�`��k2�K�I���>q#7S�/���멖��\��l�W�;Z^����,�DVNw���S{�C� ^5�(��k�c�W_�s��pũI�+Qn@�v������6Q�  ���+�#_:��У���.|�;�Ó/�6̉MX�X�5�q��\E����sN^֩�ڔ�פ�X�z�'"G�3�H���H_���T�A4��!�ʣ$*g��eZ6�2����ǹJq�|W��}���H��:��*�W�j�OC��ri���^i_����1�7+Sj� �C�J@�����9o����џI:�*W�z�3YX+�+w�+.A�)�h�.��Z�cN�	t�G3"*.mXM\�m���Yx�.��]8�z�1x��o��ӨP�G���JF�X���Km��<{�ux����k<y�w�;O�����]�	��MXoa�Z��_M�[��&he��w�EEh]�ʇ�7���.�r�-ƭ`�i�܂]c�&-�S�c�_��2�s�n��C__�!����6��ST[��7�
��b�T&�f	��Y�'��Q<�&]��᱘uV�Տ ��\�����ƚS���S��H�[n��t�[���9�C�d��PY�[nFi����8��'��ڳΔ6����ZH;}^�5F��%�,Y
o�7��F����6E9GG`�����z)���#m@���<�m���0��B���d]��$�B�	R�I�+�RE�7��d\�N�	^9j8q����:�����wR�>4��{���6<;��W:�G �
�ܟh,b��]ūx��x6�y0o�����w�	�����S;���g+6��Z2�WĢ�U�����̷����&��-7�ٯL��<$`稂I��=O>3�Q6�ý�1�&2W��b���5���p���G-�p=�S�1;�)�@�d ��ҙ#��s���o�pQ{�|��d�8�ռ����4�w��Nc�%6�fAoEħ�m�v6��"ްR	�%�(���F�Q�)�&���'ף!��W��Ky��A����
�K��ʟ)t��5&���˙���z������OO`�*�3-r:}��)� >j2uᾓ��,�ޔ��hLI��+jc|o��<�nEn��Q����3��/����_:C���}
y�%xϕ��%�f�#8u�����Е	�:���X���_�{�������}��LO����ؓ���-?�;�#���H!�0&%|�
�I���7��9J�C�)!�su�U�i^]�#�Ó���!r�2�d� �x�rJ����)�ǐև귰؜R������q'�뫴�"�䳜�����t�}'�w�DN,b�i'�yM��1�o�8���o��%����:�`��&Ȟ��Z�bZ�1�Z�Mu|�j�p6&i-)&��F�<��wL������w��r�U൅^/g�v\�&�*�X�y��K���<���c��e��CO���^���j���8}֪P���kц����$��\W~C9��
K^EJ3y��Zv�VJ�.�8���l'Mo>p�p�J��?�a�:H�<G����h�  8�wQ&�>�0����R�Ok�4��%c5v����Pꁃ�Ubw��Y�u���OO�'�x�UM�G�O�4�Hǉ���!'�Ҙ�{���c�F�[K��U�&��P�±�V-?���ko鮴��>�`��R#��=p�r[��3/���:X:~�� �������;e���ښ�l��_�ʆp3;:�h��n ��m��А���F<b�\�ch��g�Kp�z�
��uײ�q�����뮀�\u%<��k���p��P��)QN�Q�pJ��f־�n��w�o8u`{��I4� n�V�;�s����^4t^;jSQ��=E�u�s��9��/�^�Pf,�P��V�R�2IiT%�o�5��a�dd�i�����;�_&{]j�UG%�R��x'�䩌_�.�Sץ92}ױ��4�H#EB��0k�?ҩGbu�Ec�ǞB�~6ϪE��Q�|���4�_#�S�AE��Ñ��I�Y#�m��Z�%[�kZF��H�A����m�� ��<ۺ�g_?��s���o�%8�D��U֧�D�AZ䉰���Y������?�U����ۯ���ԓuظ�M5��� /;L�.Pc|�^�"^�r˚J������܃ai��O�����Y�=�8��
�iX���e}1�a��Ê�������t�8�����6`#���t���p��j���P��1��ʴ�GT"9��#:���������EI�f�cL6	�L���G%�I��0 Or�;�\��	���s��������'�t�N\����n���xw��\<O��
�����g�y �}�yxew��(W^�7q�g>^�`�+Q *����g��t�с��7Qb�+����"���VZ�*����pW92�t-&($Ńw�G� �.�O뒇�<s��p��4R�YTj^*���
<n��쳠-y��=v�'�h�6'Gi�K����0�h�@kŵ�V΍���h�N��؞أ��:��vK���]�����Ta�'�_qg�	L�A"����"-��u.�촏OG�#�o4�`����wm��*��8�<��!�qZ�!�&��De��2 ��2[T��������7^_z�pױ��)>���$1X�,�y21.����F���:�����Lw��NE3SX=�c(�V���?�<�̋09q��x����C�y�#Ö�ZΠ���M������'$ψ���U�VP��fQ�ۗ/i�F:>dFb��F:�d;��ĝ�>��*+�!_�:��]ƃ������0)���r��@(�=�uJДA?cY�W�Ȭ�KJ'k�6&�߿>t�{���nXo&n��	W�^�ݺ=�\��6^�ǟ�����{��^~���NZ9e�JX3�6��G��� �M+2�_e�ʀ�o��k��[B(o����=�(3j^�����sZqw���﹔�蹐�H6%�u�};L"}���b��"��a�B�Gc�%�gn�`դ�0t�1F��1,�R�~P	2t�J�/;��禳XD�,e�ÿ_7�����}Rؐ�f!��@Y�)��S0��of�\�ň�$EZ�]y7��2�
.nV�{_�&�t���?�~8醥-<�s=<�p~k���C�G��|�{߅'/\�󦆵�P�� ��lF��ַ����z�{��w�q��x�
��a7��Q�8qE0/7���/�����y��	��c	�7y�F��l�)4�x�>+���p�u��� ������q�4����ҝ�S��ke�BW��HFV�D�����#�4�A���O#	��=�y�8���q��ʡ]��� �P�j�o]J���I#+��Oǫ^K�Sn�MC�%v����Q�t������Lὖ���J2 %�\�_��'Ν߁�w�½����
K+N�U�����\�<�|a#�%|��
9�q2`�t ��2O0pʼ6����p�u�Î����6�Y<��J�n�V:�U��e�KI�V���n��z�͑陈���W.�p}���E�̗�
�l֕���)%?4�)2Ҿ�uL2{�o�F����U&���AFwǹ�Kj"=�J[%����r���[�����y2��lLf�W!#���#���w�n#�4��4�qT~m��W�,CC�pyx���XWz���R�z��ƽW��J��ex��X�bI9�;�}*����a�E�%"�����Z���d�����W���v+��:^;W�+�������W���~�;��߽���C����N�k�`6��U(�QWo���3>�Xژh�QU@p>2��`��cاEV�#�yt�$��J�]{0&�n��Ȗ��I��O��]AgZ*�|.�L�'�(��|��4��L��-��9lI֗z$F�'�"�=|m�����0t���`G��p��wެ�E�\�n��Tن����)�t�!ڈ~D����R`x��ݥ�<KJT���������0\��$?15ɏ�*�
|:K<��L��'n���qw�l�i^�T�?�o�� �����M�ºWx��-���?��=��Ǟ��g�%�`�lq
���TA�ں]��1ۄ]�Fq��b9e�����H7[X�dQ��3�n@��4����T�Zlew�s��sn(K$�\.Q���LxZ�k �y��j�h��q�s�s$: ʇ�&���w,��{Ʌm��ä�\�^�U9��uY_���W�H�o�.�G���1���1�N���}�Z��XZ��Ae�6m,[`I=i��F*QѻЀ0�E���dn���|q-�b�-��D/��хL�"	��	�OK�%� G���*D���2��pbE}�K��?枢eC��� ��QJKER�{��Dy�rfi�R�@R��z1KMH��V;~�Ex��7z�f����2S�{�q�r�,�UY��{��'-�@��zX.E�0RN�&��S��O_}5��s���W����s��˼pۇ~Yô�ᮛ��kO�����$/
�X_�}+7���|��g`w�k\5�z��U%�Q%�0p�p'G��q){X��2�F7�db�i!͘(���>'�r��dp�I��<�H+)G�_�!��g{%��3@ʱ&^��6c8o�Q^�4'�Bg]�nmH�4�H���n�~ǲ�ŋ�Oqh�Qq9�-�^9�Z���E#v֦�b�{�x�������Ae��HLq � ��o�l��g/<Lt�=ſF�b�su}�ۤL�eIX���Q颽ya���@I�V֨<>ڝL���������?�a���7]s��f����/��}|��߅�{	��T��`k�G1gT�8D�� l�>��T�^P^W�h����W^6"��}��Ju��?}ݩ$��)zn��,nh���y�{ u%]�bSN=��.ʏ(|$J�L^g��,�`�!Q�Q�kwb^|�y㹬4;���$��!r��{�NH�AW Y'J��%���!���٫��5�r8X$�>x�eq�^Β����B�&�A�Z�`9e	����J���	#�F @|�w���?����<���p����.:�m8Y�ub��w����p�ɓ�����Sxu{^8��6�S�t׬4M�ƿ�^i��F�3b��5�ZmT�=آ�?�D���j˸�1���C����	��ה���_��! y�	��lC�%�4�O1P��?��d�lpފW���TK�f�E+̮�D*����wՖ��{9�I�4�AWܳ�\V�Ϋ�Ej���ԉ]��XW�⪛6�Fi�cF~;Z�LF%oTj-�(�'*���ᯈ�!)(L�J���6�Ě1�h�(�a�U-Y��=\{�
�+j�7�z�`����^�N���3��=��I!z����ᨈK[h���7|~��'��Ȧ;7�<� ����$�T`�-�����Ix;����(�	��`��*X�*�����Ymp[`�]W�HQ�zc{7�>��pp�L�8�኎�Wyy}����:*u�X�T�R�IY� \�9��QlN(&�����
VU��(�٨Vzڔ��\�C�o�!I(%`�Z霋m�}�Z�*��2�?�{�ѨR��&Z�χ�֩�	秙��R�4�H#u-w˩���d�l^r�V��h�+�y]���vE{���/�K/�@6��_�`a��I��2�u��y�ǰ�# xj��H�I���F#�p��AQ[��i`6����]����s��7�Wll¤�����6�xqf-ƾzN �@���t�	y!FAPA�ջ?����\�#�<�r�Z���,WUZ����y/L���*�"��C~�v���!�ʞA�Պ�{0�,=ܐ�K�Ɵ�K��^�8N�m)�-A�G�!^B��^7p߁l)��H��W�-e��T+h6�h		,`(򵬀iq:���k I����&�0�s�T,�f��G�E-_=�8%'~{�f��������'�fϜ?ͬ�:�Ԁj��I7~����ۡ��?7���  Z���#�c���9>�ƈ0�'%R���U�� ��$P
jm�c���W�:,�����3���4i_�Z�� ���A ��z�������J�U!�d�ǅ,�.p(�b�:7�����-�<ˑ@	���<�/���S#�4�A�\���ni�zJ� ����KOR�!����og����[���Ր��G񍐃��H���RU@�7�2�+��*^xbA����eo`��ɻ�v�ԍu����.^�[O� �4]q�E���Xi�H�u��1n���(`�F�F���N��+\*��3(��V���s��o};�O�i;��0��H�R=1_!?�NP9v�zx���a�8ٯ}0��}�X6�Q]]�pv:�����>�k��ʔL�IW���HCu�r�cB�#t�+N�K Z�&奂��*S��e�S$��<�2�U�@l���9����pi�	��p�Fh!��Sn9o��בw�B"*�+�h�1�H#�Ue�޴K�WGs �|m���x�,���W��] 	և'��zH�+��PJ�" �`L�Sp�>o��{0�+����Xo�Y�ï�ES�X������L�.�pu0�>9���T�P�K��$x���n7��W�D�Ry6�yD$(�c/&`�&ك��d���D��e�$c^�����K������]�򒤪�w�b*B��{�`�z�g$W�=�NC�g����ˤ}���dಡ�8F:D��P�
�� ւ���)?(^/��3�J��"���eo��1�U�����P���Æb��ܐgw/�����CL���O�o)�Nѻ�'h R	`P+O4<80�H�䵃	�I��,���u�-�;��C�D�*�Gs�ac:�W͚Up��}֌�$� xB>��4�Jd"9L�,�{�c����i�ta����������-���ޗ�<px:#@6�J�,��DI�,r�Vȧg1�Y�'c;*?G�r��ӫb�+�5f��7�p��(���o�ISPXWŶ*�^iU�4����~˘L^�3B��/�ѧO� ��W�rN�[��C��18�e��eTc�%�i`����+�����?�����2��Vv���l�#����*�Sa:�jr���F�2�
�����0����v�濿x~���|�{az��,V�&� �h7��6�.�X��'l04p�M]��/� �_� מ>0u�#��P�Ů������૏>��+�u3�7D	c���/�h�J	��˳B�֒~�z���c2%���xB}G����r�P7<2�-D���k*<eeNGJfRu}�Au�^z�db�u#u��I}������n��F:�4��ƑY?搵�/�V
9�d��hS���t�[_M)5�[ۻ����2&<���2"`����h��Ҹt{0U؟i�%�?댅k�}m�vp`���	�z���pX�DEy?���j��y�%38����&��S�N����~
����,��d���$�P�	�H���E�z��O�`�kጪ�$�d���,g����cڌɥD�me2��a�ԣ�u\ǅX8�6H˔7����������/��خ�3�2��}���>�s����R��aF���sHXK۵�Gd@�C�6��n�a{�Z�Ƞ �[��?y�.��K�P��jB���*��ėw��Z��E��x�l����"Ubm�;��<�,Eީ��:`c��w�����R	eeb�<'d�O�xĳ�w�	�%�$"p��}��tӆOP�Ě/⧼�0ư��ȧud
cm��s �P*y�p���JBD��qA�^y�͇�b�>�U�y�q��a(�E�8J��VN���5�H#]:�=Hl�W�)8���r���p��V�9x'+���|�R���(�׋\��%�8n��A���yd�����!�67�E6�L���9ø藀p��1s�Al)�q�?�UUV���?��^8�~�4�lM��_��W��'��_������`�.�p����5�kf���2��{��5Q�e�T� VLB1�r�O`�=`����o|���/~fל��NZYmF��˂y�nl���ï��Z��}���"\{�j��p0f�F�t�7���^����/��ں��Q�5 �߽��I��\���Tj�?�P�Ƚ&����:����b5ʓ6)�"e�����!e<[��x<����O�:�s	�<�*�!�]�\&VyY9'�]�P��)�Nx�I�!�/ќ�Rq�i��.Wr�R��:�����k)[(�g%�"T�O\I����\�jm����-�	����-���9��b�|ߌk���۴t:_I��_�C\��)E�ω�������폈� �9�'�`(>�+2���:�N�O�-�f���d�'o�,�7P�
�͔-�Ee�}���m�!v�R����$��nbK?�QVx����������qS�&#e�+t~�&+�
��aD)$��d��2\�E6�ţ�Bf�8�Ir�3��kD��PJ垣����=�	�2�����������u��U(Ģ4�8�y[����;�2J�k:��|�f�C�+%)���#�I0�|�?�!�*�nb:�b�,4TM��,��2��H�f�#T*Y���(ܽ,����>41�������Wxm�*�\���R����j��E��$#���zU�s0�TX��3p�2e�d�w�ڎ���|g�_���|W�w,7�~y�P 4]�%NRFMQ{��M�(�4"��"~/��(/�)�<p�F��
DL���敔�q�LXLŅ����D�:��~�f!��9ӧM>�s�޻�J��A�x��H#]~��{��g�;��ϥ %8&�*T�X���8���Ԡ�ń;Z	_ﶕ�!Vz�8M�2�K}�����5w���q��C�f�J��n��e�+���-��� �"@� :Ў���3�`<
AƢ�w�2���_�Q��'����?��_x��'~��z�܀Y�D<��	׀8��3�p����5N34Seg��.-���2n�Y�v��M��.�Z�F�ag�<�|�s_����`��+�^�!8�f�.�J6��~R�$ud(T2�q�0�v�����yg����[�$�8��vZ���_~�;w�-���#���Ȥ�$O��2�;-B�@m��r���������Vȟ<��b�F�C�8���㇝���\f1�m�/��2+�?�?
�M� �
N���՝�u�
���i���,�~Fm�y�bI�b�]���4�H�=��a{��)�krb���4HF��o��&)�YJ�c��]E�(�E�<�}��$#�*�[��P:�5�?!�Ԃ�Ƽ=�Lv2a�Է,�=�k�y��=�u
d�b�NS��������������gC�'�ݸ'���3�N�k`�F`_�бĦ@V�6����T�swQ���@�>q�Y�':r�%�	(�4&e�Ƣ}ăjXx��4��S��f�����.8J㏬O��ҨIʝ����\1�1�}uLU�?��g�$˕Ri>:}U7�-�y�h�����cA9?����꣊�@wFd^��]��$�ʎ3���a��V�pyP���A�S��Ġ��>wć�#�4����a	@�'�i�:��V�ʋ��*�5�sd߲\�"����l�Zp"`��*�
G�
*n�$=N_�
�ד���]�\+i��Nq��d��AL�琅�-;�x��L�i�D�i@Z[�$A�(��7�_������R\�U�هW?��r:��|a�����J���3'@�B�-���T:�jZ՝�#�4��)���~��AҸ�'x��\͙b�֘.6%x�B�՟�z�z8�3�a���y�J۠���ʥ[F=��%� ΒT���~�y�^3����&��ҕ�)��tp��6j��C��ݿ��믅�^\��	�'N¤�@U��S�W��E�~<R�,U�W�7�F̚����)��m"�;f�}~ak�n���/���/��Ξ�Ϟ���5��'�:6~p�Y��jc;�֠��B�a�!�!3��s�M�&�{_�4����c?o�����*o\b������矃O}�;�[m���W�+�Pa� �d,����R{3)ega.)�^RN.	qR ���錀��J=���z����9b�����{�0(��?�a�iTB����<ø����T#�6��5#�4�>Ҳ3�CT���z��zѭ�J�R�l��K�B�v���{%��]U�~g2
�C�=�J�2N�(��%V�,{O���͠�bl[��fc�/�A�z �h��7��E�Y�APy����	Lҏ<��N ڸ�����3F��W���K���p/K�KTB���ۃ�r�|�N�g�Mu!y��Ky��T��Iʐ�#�E�	�I���_�B�ӱ2}�W2���%��OeD�3�����T���t�*�~��_���x�uxu=;�,v96�[��IHzh�-/�^�4��=�t�@1mT'���>緌'����b�"תg���UA��B��VƕH�ę�D%�\'1��t���zg �`4 Q	��T����&W.O,�[�	�̌������{v��I*^E��`�ȥ�%H?����Q�Y -Qw�-������@Q�dLt�B����v/�K�����äGf�$�1�v���|�a:�H#�t�)p��J��{�Ivu N��x�0���}�h�k��uIS[�nԫ�Kd����Ͼ�C��D��1~�ȃ�u�
�����۰m��G=��C�NL��n����	q�ث^+RFV"_�C�����o�����`��X��®���%i���:	A�����[��(�TVnik�O����)�C�V���?g����|�ѧ�o��;�=w��|���/��}>{��p~��ڤ&~���o{�G	TL��Me�{N�+�x6�%3�Iŗ�-פ�J�P_s�|Y���Zӂ����Ś�4��~�����e(u)���L���2�H#���%���c�<�3�B}�<������fۈ��sk#|�@��E�z.��i�aۃI�V�Y>Qo�L� ��ʰ
�� �"eQF�\��j��6������q���ƶ��`��V�0�
��l&f��������3����6I��L���ƀU��~�K��P��{0y2o3Vꉀ?��df��5#�Hwԍ�{��.½�sLh9�}�ń��W�ɾ\��
���:����_�ŝw"b����<��g
ߖ̽�YI�))2ճ���
#!*E	 �tc^��,hB '㪈q�N�5t�4$�v�Մ�I#�� �FteR�Zē<��)\QɈ���*��Y���9$aA����K�"� ��K��G�i�ߡ�2��K�E�;h�(�F��\Ҕ����3�V[O2�D=y�2�X�Gɪ�8��i��VDv��y����=])冎���*��e�M���I���L%�H���s�u�+}���'�<��P��wZ	��S.*u����|.$Ri�l�w��в�j!/Lj����&̚�!bw6�z���h�����{"�"�A�ְ��Nڙx�Q����h+翴r"�h�2����%�2;��
��0��ڢ�������j�_wW�8�%gN�w�^�{��e�|�pjc.^��zv6�����mx�&� =f�)(r�7�h3)4t��R��,l���iHI͠G٢lD!��s�Ψ?6h�[�e$�Y�ǊHt����#�J2IER�L�+��%)t�LP�g:Y��10 ��4�H#-C�P\��+��t�σ�)��Z��T������G���nכ܈�B��\?�2��_�K�pr#�h\7�Z�}����`*z��(b~�U�=��5G}G�e�B^P�"0���I�`l)'��t�>���$9ʽ�(]$CX]6�I�ŭQ�7�����A���d+�M�E��1#�BE�ᆨ���u����@{�Ǘ��GAv*��X�)�~��"�-n�������r�5W�,��ɻ����*�R�P|�5&(p �T� &�7*	���P�e�pu2�w���P�@��c�r2��òBh�P�w�[|��Q+w�:J:Ў�) ����X��9UiE}W��9E>���� �-��|�L�v��p3a,�{�m�
d��ڶ��y��ώVc��X��i>ɣ�S�:�+\Y�}U�5�u$���E$�q�Yu�nөFQ�Ba+ȿ�K�%J��mh����f߃���[c�x����i�ڀ�����fU eDR�'Y#�[G:�����L�/˲���c��ƨ4�7�+$�|��i\!�,�	�Y�E�=d)��	���J�ƹw��(uE:$������ ὒ�փ �Ok�g��*��,�\�"��l|�	F����!~�
��_=�@6��<rH��o���q U��g�������k��Y������\��<�/wȲ�;^�u!�x��<�ϩW3i�9w�A>�&A���b�^o��`��2GÏ/�A]���l��uH~{6Ҟc��'�X����l�MTI4�Y-eY�G�� 3*H��`d�9�sPqx`�W��r�g,3yW5M�$�r��������h0�ޒ����ȋ��٧)]���K~*��E�������*ϡ��q�l�.����F::tИ��?��|�t��҂5�rLQ��M����U��\j�c�5*}	�L���҄�s�iiy璚�p�E}d�gN�f8�. 򂞃�� ������n�&��.zκ]�A�-��9ĺ��Ke ���
�_d�{0���F�SCi\KX��'I8��� S��CUgu6X�Ǽ����-A9�Ɛ%1�0$;�,�4�������6�����5��Ϥt��7�x`D]cلD��;'a#�Й����r��:�9��:�b�;��j��e��Q%'�j%�^�?<u�d��mi����]�������=p���J�]�,�~�H6 �xg�15��$�Aj8����9��d�.U�I�ܫ"4�4��ߴX�X���l�dqO��!M\)��*�h@d:]�G�X��qX<�)5]f#T���� hP�j��*�?��v��Pu%�.�K�&^�����ґo�zi%�$���l\�B��\E�E7�U亊�h�@�)�;Yǥ~����,�P���j$��$��g���">���#>j���"n@��.�z\��󐼺IT>���9ɪ�G���sϧY;wn%�%�_p�y�i��]�ڋ"{���9$, +OE�$���ގ4R'Yؓ�O���^���;�r��x��@
N�q�6!~�T����"^�(j�\����wB��e�3�>��Kԧd������κ��F�e�Y�M�9bȤ�/"p���=��OE#��G9_��#J$�e��P����>�Q�\�a��r�ֲ��2�6�j��w��A��)��5���`�,<l�l����Wy06�����,���ş������s�	�5Օ�ڄH�cI$5���+�U!�L$��� ��WA��6	����썘�j-�QJ�7��ju4A�4���b0�Z�*}r	��ʹ{6�nBw�hC��m�����E��� � ��3첵(�] �E֙E��`h9���<{��Yp,�H���RG����F��x�N�@X��E���9c�SPt	5��iJd���_y�U��XW�#���He�CD��!�<�Y\ϳ<H`��0�!����.�Ăċa���` V|EdT,
g�zǡ$�Q	A����Y��Jv6nr�43�NB�\E2����8��2I��l�7�j'��h��M���Pf���/H����V'��vJ���
ܶl���U�D�j�4�_�`Y�1h����wQ{C��T���O�5��;a���1��.ۮk��,@C�H�,A�I���Bz{�Be���TC��}�L�3QR�)EB��Q�A�f\�����J��R��(�n�J�w�lN�$��\��޲�) =Y�))��x��>�m'h���S.��&.g��L֩
$������@�">�^p<�iX��J�t�Vѳ�Rk�4�!c?�ܽ�n�u'���o�?}��Mn3��r5z�Qu�jU�TL����$�W��TS�@�l0'�C�6JGI��ZF��l���� ˖a��,mN|���E�yN�MR"��.7T_9RP�
�S��,%j��P��J��0�d�#-K��;�~����F���<#�޴�\~Xsz	+\�481D�I�2�4��a���i@R2R/���o�$���H�$���T>�<��1�Tx�9(�sDbT��&a�T�p1n�ٴAV���c�L{��2��u��̔r��~BC#t
���b	=x|��
ը��jt��`P��4�����\"^���,
G�\~P-�c���$h��
+"cQ�eo#S��3�_/��'e�B��3��\�r"��הl���#(�q�S_��ʀ�UqJ�H���b��W��ah�/ER~Z$�~�=���a�}}a9����Ž��м�+��9ڤ���x�zK\�9^�Q������pE�4��)(�܁�����q�ϒX"^��y��\�RiH]��L�ⴏ"�`�����P�%�CĘ �Z��N,���{0�Wr(6���+~�KCa|'o4�� x�=��R��D���c�k�m���g�� "��+j���x�PB�Qe��i������t�?!����Hd��GB=pIӶ�M eEy,�>Ϙ?DJ�hGa�Y�R�{��yN�V�g2��ȶs:ɞ8�kn=ԛ}Q�OO)�*Ď)�씩r2=Ũ���rp\i���k�7bb���P.{�_� ��)��I�=�vƁN�)���3lL�
��i��3d�y(+A�Ư�S���`� � o��` (C�j���m@���{�pw<��������+�ʟ���E�0����-W�Lڰ>$��](�/�7��֖�`�\G)I��2<H{�^eY�����"�%� .��BŤ���t�'���K�b��t���Y�>��<7gi���:UV�g9��wCx������A�1�#a:�����ҕΐx]�a���XPW��m?Hr!��tr��QX���lbܗ�eA~MZ^�X����Z��tQ�/�"}X�'-dU�R>,J�I�o�)�H�\�.r��BH�-��x(�4y�&���%2�f��I�@c��gu��G� ��>Qq���">��Jg#���'VU;/TU����.Ȱ߄0�=��4-��N��i��Y�G�_1@�:Bq��)�z�LO�ڃH�)V����%:�ƲO6A�ޔd�'��*�΀��T?B%=wN ]�1��H��ׇlLw(.Z�G��e�q�H^Xg�|t����~6�_)�e�1�/.YG���c1�&�n>�3.8��
F:$tąWq�`��ht�K��Z%
�9M�1꩓�Qa�����=�S�6��P��	L���3�x��"ͽ43X5N��ޛ(����c˲�/�┟�f�xnW�m�T����=�үq�����5h֍߃�63�c�L<(��8�R9Sp��e'��Њ�+O��2�¢ы�W���"��}~��<Q����Y+y�p�h>mv!l�v��[}�?�c�H:��8�	@`���c���F+�z�X5Y����r�W	�TY,	�m�b�_� N�n��|	H�]�oqದp0�AN	�K���Dyd�e*��I|b��M��$ �P0��a���IB2+��W����v�w�5����v5��\%`4�0q� �ງ���Q�<���I��ئ�*�6���  �n�	�3f0ݺk�)\����<	�\{5����\�[�P���;��kg����W^�sU�|�dЋN,L�b�+[0Ѿ�8�7_T3����dLl��.S>lM��*��g|U�!Wc\��Ӭ�_�f���F�%�+���xM�/x�=L�^~Ƨ|�'�(]�G���Q[�3�M��_�u"�kG��U	�*J��c$�q����B�6���cQ��i��6>3��>6�R�%~PI��N����r��=�%@4����/�V�Uʶt�
m1��u'%i$����6�<1�!�nHV��G{Ҳ��n?ںː�OI��L��P,�(f*���dӇ)�Y �ٕ[�P��6�Qq��B%���p�kلkk�|B�G}*S�i�V��/�8T������h�[j"����M��V�)GN�f�%�۝��X�����������(Kc����&31|�|�-�&�,�6�����(_u�CSz"I�ɹ�����m7D�4t���@��þ����s��+�t�.y2"y�G�o�s�hU���J��,�7I[�5�V!����F���A��C���TLg��g�����pt� +��;si%��VϠ<S>��i�a~;&	L�̥��Y� �<H�-0ا��G�"2��6a�Ƞb�{T��?GM���cҰ9V�ֵ���G�x�� �￸��ߠD>MH��a�1�X��Mav��h__��	��>	o�����I�L*o����������W^�'_zv�O���? [�Y���Z���[3���Ԧo���'`+t�F����B�F��-�|��`�Lc�u*=��?�6ڻ�Va?&�G�3�Hh ��Bي�F?�Ŕ\>��-����n�6��'fE��q�H�����Qb�!��\G���7�r�6T�����`���M�T��n��<����m��q�K 	t��Fʼp$��V�᯼ �O�޻o�V��R樂�J���"辧T>=�d�2/Y��L���f<�N�r��[8�Ӊ��sfl�����"�X��EƟ��<������D��� d|a,D�T+<������=�ؙ��m?g�p���zݵ�����;o��t�)�����O�ɵM�� ���h��Fm�ƫ/��/����{���p���S�����t�m�z�?i󛸻�+��v�U�#P8�U'��ه\T~y���B�2��4�b�L�����)����r;e�6J�<lcJ˽����@2� ��:Fun��0M�f�v�A�&��f@)&'�����`����Ut�-0c��0v�&����^��}�_j7v�8fp���t90n��^ۘNe-�L)�t���u��˔c��JtP�����2���\)�O�8x�pT⧸~b=�	��+�;�R�C�6���Q_�W��ѩ:E�~�p�8z�yC��"����#ĵ�Ni�!�XU�57�[e�_*m���]�x��4a	*ɵ�E���䲕ꧥ�
���J¾!�!y�r�A����.�A�f��LՍc���W��.x����e�2��"#kÈz2�m`�HF���q�eKA���yP*}��E�D;�Cr'�O2���G3m1����]��ݱ��K:�.9h^�!�� x/����� �ٌ�E&���>��#���}�V�ߥ8">kHMG^��&j'+����2�(���d>s�&�~�����p|W^{��#,�w���/s�B_:{?}|�7��CO�i
>jD��6�-�>l��5��7z�Fl���VB}p-;l�غA��@b�F41��<-q��Mw��y(�9y�10�r7�P�-Aaa+�����w���|��SgNP�8k0�j�i�Xn��1�<]TO��B̶$a�Հ��<��}	�*p�ƽ��]�	�Lۿ�γ�c��N��;o��v�5p�o��<	7\}5\u�$��l@�b�ڍ'��.\܆�/\�'^x��Y�������^�g�m��Y�u���;\�*��Y[��JM�~,]��Q�mfR\*�A��r6�i�G���}�B����N�I����_� ���K����K���R�/s�hӏϐ�0$�e<��T����!��A���x+#�K��I"���W�NgM���I�i��T
���p���y�a���2����Rg���)N���,XY��{%�h]i*)Ӊ pV��s��&-���j�eZ�o2 ���a*flg���#U�˕ A�6L2���@��\�>�����)*�g;�i&�Vװ5Lw,LN���7�0����LpqeqAH K����8�4�d�9q���%6����v��.\����7���6x�n���x#���i8�.��l��`!:�mV��ڠ�=��g6O�[�p�;w�����׶v���_�o�?|��'��O>ϵ cj��N*�m��Ͱcz>�	 ��Sl���\:�'�g@9�+Ǐ�P�`'��k���'0Y#$X��uɊRRcĸ�yE�t�*h��҆��h����Hs!꟟��u���"q���=�H��
�mJ��%k�4�Bd ����/f������0���&@���P|���h/F�T��^Ӹ�-R�}��|����vRRd�Id��)����[�6y��e������J6��wa�Ҩ�
�x��-sDפ-�FG�T�o���x3���'�9/���'ǐ�=U����Rܧ7�u�|��HX����R�<�Amc(+	�D�4V	��o�ۉ�R�ZDT�^����0�/�T��^��t"��t��w�H�s �"�ˈ�Y3ٺ+:���:GE�и�I*�Ӣg�$��c?�r@:ekE��PO~}��HK�M~����!�t�cOr�*ǔJ� ���'�J��&J�iu��>�����u+���z�������%�	�����R�y'�Y�@��b�����ަ�4B�a�9:w�{�|�O�pr���ݦ
�7�4�>������wJ�@J)_��Cפ�}gP�J�׍��.�z����z�����o���x�as6'-onƠH�!��h�x<qr�9}���ػ?>���m�CO>�z���OýϾ��y�S'�ޓ�͠��nƥ_7|�=H�_�g'{�\$(l|kثu��e͉�!Ո��(���Ŭd0�M��d��;��=S���8���v��ǲaU����QϘ߫ǈ!Fir�P<TĆ���� ܶ�6q�ȸ�[g7O���e7���h)�������ω�|#�H{#iaYz�9�+����i�}߽�T�?{��x0$�w��8�I�jI[g)ƓFR6��]�3�j9��X7�Rl���.�k���~;|�������3�¿��7��W_���⹾a��q��Z5���O��`&X<B��lm�D"��&��1vwaz��������O��pf��l˹�h��l����͖��B#�n��gg>�F���'N�o=��6o����/��|���~�k��Nզ�&��L9O^`&T��L�D�@� ���>���G4�jSZ�61�&�v��z�1
��0�}�G�&�U#��j��N�oE>�ꜻo�c��b�J���Ǝ������+����{��G)��G��� ���w��k�^���+�
	g�P-������:������ }ɦO�a�W,�ۀu3�g��"Kv1��B}#l
��3����t]��=�)�,UyH��(�Z���J
ᄑ=U���^:tZ�׏r3���J�$5�� 0�Ps��H`�TE���nQ�)e�Gˏ�2؊�˴%s�+���G�v�#ҡ�DgjW�2��ܙɀ��"�T��h3��C�97�I�4YjC�蓉sR�%�弯�h��^u��/m�����M�wsz	gϴ��K����aP�Y�_��>0������usY�������Q��}��Q�9�,�%��R  �h�|TX��dN����ҁ�'a͈�g�X�Rc�"�q�U�3�� ��w���ly���{����ì��ٹ�p�������^��҃�7�W@|Y�|~��`]��N�>��s��o�'����o��5��fS�ݙ�Ň*x�@H��*��6�)㽩ՓU��\	o~�5�c�}'l���c��?��?�?��a��8���{e�{0uā�sÆ$�B��hܓ�j]�4⸎���C�'ۃq?ɹ��	�l�Mh���r�<�kb����c��D=�W ��C{�}-��:���.}J
�cP�G��a���b����~k����]��X����p/k`L��7< �Z�:�J۪daT:-u��A�v7��>z� S<]V*��M�Dm�E��	�LjB�@B,��_���m�hʍ�]�����ҏ|�x㕰�B���;o�~�mo���>����d̜k+,�B��W� ��2j��B�Z#������l<�M<�4�ສ�_��G���'�ƫNC�8������iĊ�݂r�'�m�NG&�	�ڗ��뮃���-��w��٧?��)��q
�d����i�Gb��v��8��4�B�����s%6C@��ˑ�(,.�_e�\�Y�E�NH�,�&m�D�aT��r�P(NXt���d�u�io�����r�} ��}��ݼM#G�[��3#����PK��NؑF���煈��SZ�Vi�Q�e���u�+X?��sQ��걀�R9gӻ���;�Z�����~�$��us��q	,��-$��G����YA;��
9E�֬9���$|�8Ҋ/#��n�@��3�\#��CX�e��/�_��Q�h㉹�x�[i�M��T�).�橑�\����U�,�C����S�T-d�ޒ˥�̸��?�d�x3�X����cu���w���ci�G�Jd̧{�b��F�L׮Kk�F��=~3���J�:�
�2|�!�L�I��<F��ȷ�k�|.���=�C,���(�q�g��n9y����Q���=9�����	��v��o��� _}q^����]������ж�= �*u�3k�q��k�]���43��/��N��_�ٟ�������L��Z�M�oq�b��
#G]���;�]�Y��S�z[G���pׯ� ���W������o���6�ԱuU{n�ť��`�%��q���z@2e0XWs�2�p��u�ۇ���W���$b[���e^���q���1m鉐Z�Vmd�y��H{��ʩ8�#�%X�˗߱~�l^�h�����pX���ޱ������4��GPchbc*w4��y�5ܸ�����w��,�K���J��p��Ku�$�:��-:�8Ȟ'_q��z!�w[��RC՛�9<�iֶ����G�?��OÕ�"���Ŭi�b��b��O.l������7*X����>��\R���e`��M� ��[˷wZ�p>�֛�?��O���v'���;BFt�u�
P����&h�9�&�0F]:��h}�mo�����������?�yxpg�k��9���4U���c���`�u�|:�*��BS��Q R�f	4����g�~S��	�� �9OGh�� FNU�Q��w�q�F��F�B��g��q�P}�D��, ���a�>D�������c���3�����	�e���W�]
MiYZ���,�'BL�V	��߸�v*[��<�+#Fi��C8��|-�5�}��X��ڷ�d��O�٭��#�����VO2-B$:5��'�8�p�g`��O�I�&Ie�����ēM�j�.�e�����ܺ�2X.��)�s�8~P4J����H
;�3�Nf�!���G!��4%op��G��f���1hc��Z�K�XXēe�i�Z�\���2^"6�Ra�"�e2_���C�a��Sn��d,�m�^eK��l���V�*zE��g�!�F ��Ĩ�"��$*�I�B�7)PF%%�t�!�e�����a<,Ʒ�w���F��2A��W%շ̦e�zų�i�\���ܼ�İ%�F�XG�[�4�HM��\&��T�[��>��,!t ��[�(+ ���5�(�V	��w�^��H|�a�iyF��$Xi��`�f�vgp��?��O��~�0iv vvB:�]��������g���O�W_}f'k�ǭ����sn�fV� ���4O��S�m�̆�;p�ق_�����~�������^ϛXVR��B��ܻ��{��G�9������r��O�ȇ�ݷ����~�{߅g&�PM6�D�Ӈ�&��Q/�y�G}�u	�<�\�rA��0*�Er&I:��R�K���?'�w��tjV׽�D�YX�>��������8��k1G�� #:x%D�ܡ���p�3I����_Fn���2���;��ZP���Bw1��,t�R�d�<���Y�-�J�d`(�ǕJ�����}�� �NrR_ 1���)S0,�?�JJ�Si�Ѓ����ŁZ��hw.�n����O}ά�y��-h����MW��~�?��c�x⇵]d��lq�6 �	��ΐ��rx�aܝ6P����M��}�g����ᴋ�7��e#"�~K��yc���W�� y�"-e���+l�?s=����,��;����}��������v[��[S��MIP��`EP@5ʻ��/d���j�v����-��7��[N0m��P	+Yc�mE���4Dyvd憡���9�r;��x�^WZ&�11���Y�T1Yz��F�߄�a�ƒ���Fi��Iى�d���f�ͻSFꔾ�(Û��؋}IA�!O�ub�8ꧨ�YX:��V����9�j��V%�聝C�%b弗�Ą�O-��ٔ[�(�ֶT!���#�����Х
)>K��M�i#��Q.��gF��q��Z���\D�e%Ws6�1����e=z�EE[�8��M�Y��8��T/ �&&����btԽw����b��%jFA�e���Xל�`��<�7���2��1zi���iɹ���R��
�,i��5r����q�8�H�VqaK1鐅�; �� �Tb�LQMk�X�K���2:9ٸ��B�^������?�P�p�4Z�B0fW��z�M������_�YS�}��[7�:B�5�!��`\����J��z�`:m`m{n?}��_���;��nhz1�?i��'a��L:,�^���*&%6~�+Y�6�	�~�[���7û�~7�o�����ً0�؄z�o�`꼢WuH�<��|u��>��XR�$����ܠ4�����_wI�&��<��d�8.�WBJ�-�`���u���"�H��3��ѐs�C�Գ�-�!�	:�R��)�������N�Is)�8�J�cy�'|KVRA�O��eH�>�杞���؄
p&���ߺ�>�)��J?z�TR���E��m���V�MV5���|����� ������n}Y��o|����+_��Y�h� �48�'8��og���Դ}b��uM�K����_��'~�a�]u���Zop�xU��E+j�L��N4䰑wR��t��6"fP�<}�֛��~��~������g�����UU����i����	�"���,�5Rz)�<]�UZ)�b_�.�&�
�Úx��];� ւ���dq�j��9�Gbn� n�f� ��z1���W���ǺWXװr��-�J�Τ�A�����Fi$I6��z�9(ڛ�Q`\x���9ʤ���eʴ��9
��j��cM�#�W���K����.���F)i9�򦂘L��@TL��:�Ȇ>~���w9|dj�L�W�����9I���c��6�+�+*� ^dm�$�I�&�C���~��oa��!K?�jR^��U)�(*�R2�<�oĸ�F%�0B�2�eD��U��vo�N��,d��BI�\)���l���Ѩc��F���(4��~�d�:E}�H�S�B��`T��XT]�MX�o����ޓ�.�45��G?��'`ܵ�:�/�,ujs~�#����'��I�3[A��h�XP�Yi��V3��B�u�L[>ַw��o�����pǵo ����G6JLCl��v*z{0R��W@�����*nRL���F������o�����o��{
.�5��fP��J�����o��e�>���(�y��1uYW������,��z�(C�j 5��Տ1�,7����<��(�J"94��?4�/��K���BK^����{l��ze���|kmQ:��_�;%���>_$=��{�%xbe���.�{1��BRHTXʍ`b�x:�ӛ��Fʍ腣��-�|�[�B�b,���CT��f�c�y��W�	l�,�&�j�Z������X&(���(�i3���ܲ�	�ï�2����.�So@!� �@E#�rC�"�
�\��
YU�\)D���g�M��ˮ�Ϲ���O=����՚� � �+�FJ��f�
���J�]��)�*C�b�J*E�cp��`b�dK$�� 	Ѣխ�z���{���Ú�������������s����ַ�^{o������x�p��������E�3��#Q'��U*��&�m-����ǡv,<��fI���3T�h�0y ON������J�1b��'ұ:]#����T����JCTr��*�+7�Ř����Y�ϣ��� 9��q30\�E��$)α�w)$:�zV���[�� !�3q�W����_5�U�)kU֛.�g����>7�L����4���z�T_�)���6�S��c��B>���o4&�v)���Bwh��sG���;Y5�4[���d�HGQ�i�`�=��@|�)���X^j������o���>uO�}�kJVY���fT��ɉ��,6����YŊ��Z$SQk4�z��oc2<Q��4�jEe։BV+��͇/-de̹{��j@� I���x�$+M�.���	�
&��C�-�o,lE�t8�����Y�'r+�:�v'���ħeIR�:�]��ܔ.p�x�����I�`[�}�139v�Рn�a �.�Iy��T�=��4�*�{���E^���Z��1
��6[��Ԣ�.2�F=���<4��2���ue����A=1����-��3����o�ѳ`�?���܍��k����G��ق�̍�-�5+P��b��צ4��q�}ϭ�\��x�}�?���Koiis�g-҇:�!X�WڅwL�{]���$Z��Z���B�O���niy����������|�`yÍ`�1���+q�)攮N��i����|���㍑��Zž4�%I��_%�I�m)Mw�����إ���-���}����*��`�aP�s@ �דF�4�69�����uxY�������MulV����B"��U��Xg��ٞ!��D �7��E���_w�x#�{�4ؽ=� T��pL�wm�����݂�_@DbH�p���n�凞t����EW���������6���|e8�9px�a�h� D��b�ApW�,��§�mlz'��	]V��ݳ-�����9x��g����`ov{�;Ν%����ǖ('U��Z�4�fz`�^��q��;�qNz+�2���M�*�U;}��&&�F[ӥ�t�Q���R��L��$�*�����E�(�vD��qp��㈳)
/:�5��~�Yg]�R���n������>�D6�W+�46�*�2ᇸ[�/�1�{�����b+��dT#��yZ���i�{����Mx6����'�A���-�>�}����r�(0�y��	�T���速�j7��� ��\���p�ᩀ�[��h,�8m���t��Z�ISejg��<m#�=f\6K��;A��KX.�`�lu��i�e���״�NS��V��z�r�����SD��tv�u�q���jj��;���2���xϵj3��OɎ@�Jk��pju]c8�zQ�3$/�@�亴X�QF���N��C߼�ƟR0Ll�-�L�İ GK:	r:F�X�<N��5���=��G�c߯�E���(��Y�C9l�S���E'-հύ�O�n}�S<3x�5��5����F�k݁�[���^g�#��ۖɠ����}�������^���{rM��	���9;n�u�0�%\�k)�|^v�9�;����+����N _�?�\��X���E	a$ʗ��$����E�l�Λ����]�	�����IX�:UK�r��$��t��v�ף"M'�?6�e�y��|ϭE���]�(z�"������@��r�ү���9�9ՐG/�v<�V����z�%;?��^�>÷�FX8�a�8��\�j�3�pW��US�1��A��*'o�c��r�:��A�ĝ��I��
�� d�#` �����_:y�؇b�44�42 WO[��tLp�G�G6a����O���� IV/ ��(��p.s��G=�,�����=۵t� +^̰�_����V�ϗ����ģ���;����k`�`�����]��>{�Y���;��^f���7�V@����v�s	 �կ�:��M(2b�aU%]�<I�d�?m�m��������t�ix���!���_�;m��]���0Vb�V�"���
�����4�C_c_�j[���P 4l�`J��\y�����:+x)���I�'�S�x��#b�i�LTk��,��{*�F��'�F+�R/%�/�E��g�ݎ���1c�\���<�D��}��fC�e����UQN������,�b>%?�0?O�]Dy�;W�� MƩ��&ځ�pW#����cŘ�x�∸�^���k2<�G��y�����2n.}_H�DZN��)+�rq��Q}4�4��a�1�q%�t�U&ӯ>���auY8�Lf,�x��z���2$�W�q��Ӥ��.�l�>�6K�Gd���;he
��u�xA�<]�!����n|v��xA֘�κ{a�%��K��I�'���l��D6dl�BS��C՗P6��r;BDQ�wi�}�c��3��\̓T]Q	Ga���#��$$��u�fL�Q%囶�Wa�W'��gK�!�
RH�,�d���IR!P�ǖ��M<F��9�dپ�k��vp��|սw��7����S�G��~�Ix�J�f�v������7�7
�ou��g��]����.�&"/�{�u�?�6i��qC$"��B�U���T�9J9�>��$&��RW5��5���4��n qz��O��x۪�[,�.�)*h���1��J�R7!\g����Q�&1��P�ǘ�~Z�>�н2��v��m�-�X�:=:E)�r��c�g%��w�Y�%�U�>(�;zatq�<���H8�Lf,�hN�'WkM#j��ӗnNN��y�HǢL���K�KW���Ӳ���
�R�O�?=l��S%�}��eOč��ش7g�@������Wc��q����Y �若�$�"uя�4��*�!�aQ am��l,g���w��7�'0�S0Vk�L6�B���y����b��pB������@�HiƆ���wק�-\���[����Ax՝�,ܵ){�P�U�6��x]J,˓P�{<��?�P c����� ��ʭ�5�{ۭ��/�_�� ~��E��9�n�X<hB�6��kg�f��b��-щ:�F�RtV4h�k02�@��Xפ�1���F�/4|Ez&b��~�C:������Ja���?Ě5��S��7A��v������m�(�A�)1�RH�|�6u-L��:M��	Xa��M�'c���� V���R@�U�ar(	~4��7��giav
]�:~����/�iHK���B���9�	�L�ՉTʔ��h�r����� LE�4�� =��y�+�Um���G)ʉ��Fv����i�h����Ux����s8y���S+�f�/����y�����+q&ZE������"�C�D���K���Qq����w�g�����ѽp��l�nAQ毩PX�q�1�0@<~��F�&Qb8��u�VI:n�>d����v��	]��W�x����Q=eq���~Ɍ��ƪ���f �j����ƀ���.|��+d�կ� H�OVA��t��*�$]Ł�S��Njڑ(>Bt�pS�/}��L#�BD�j�fٺ'
BNa��c�(�=D��2Je��~�}e��P_Y���ߡ�c�3[ì�t�X"�_C
 ��3%��w�S�� ���ʛ�_sa�"��
�'	Aa��	k#�y��T���K��'�7N�6Ie��B0��J$5�w)�4�M���_����HJ�~!�EOcz̊�Aw�(�Q_��=b���m�&'��{{p����!x�7�:#��k��\\T��3�¯�������$<j�X͠n?݉�l���Ĉ�l ��D[C�R7Ou�P6b=�i�����e�H*�k4B}���1�q�-֕��%4)!0����ƂA�F��x��V°=�d��bX��3��u���4E�H����C��s.)џ{^�Q�w�o�n�%���۴�9Z��Y���^&yN��~}!?�
e��r��!�72~�K�����Lwl��TW��'ڝ7φ�L��h]���
y$X��$t����5����2���\�+�?V�Q��W�]*�A�!)C��w�=���Q��ӧ�y~2�'\��U�1��-�����ף����J]��4��wް௯���'靺���;�Sx��^�`{��V5j"ϛ
�����Z3q�����8����xj���+�TK��}��;F4Kx����Ǿ�;���O4�Ѥ^��J��C(ӵY��j��L�aU��{��z�+�nU��M�Nc����H�NV��SƁ�Na]�}7���{.��jՖ�	��1�.^�����)c������X;���_����Š'��!�W'2�>����R�oNkI�]���+9p�"0%��Pёҕ��t� �ǅ���n�/�ېz����Z�yC����SO���S�Sᑍ7����0��`sn��?*#�/.f��.�>�c�B6˒4��J�Ts��Y,X^Z«ϝ������N���=l\@A�N�@ �󮩗�*��tw��4u���t��+�2P���pL��.��R9��6�r��N���-����/å�+{	KRc�H�&M��o�<<����G�e`v�Kc�p7��,�ޘ��D% ي���qm�簡�u~'�5^��r�SӸ0�@4�n,���{�ᩯR��k *�!Jβ�8�0�X:̏�ǘ~ͽ�3���N�~�* B�ꎙ�z�у!��ر�/�B�����e�q��
��a��
/�q�Av]@#B1.a��ptPhE�rA}IՔQCJ�0�2�W|����H�o��[zȧ�#5��5Pul�Y>�{~`h�;�k�p�0{�8f�NIad��l�ep�sm��p^y��W����_�l���w���%�۪�������;���������e�/\���ԭ>�ʢ���QW��-��9�)�9v�e|ar�Q��io��Ӥ&��+�%e/ 2U�TϹ^�l���S^��p�A�"©=)�&�������A�K�XE���-c��U*
�����T��ca��u���c�1V�-�qJsJ:��g�������}�U|>�k��00�rc��̈E�&-ۘ�d�_��g���[��k�Ѐ��~���s��cֈ�Ye���Y-^%�ܳ&����YEjU�&��������������m����E��.(�^�ȭ��!���m�������f��?���g���_o�,|}�B�.��p!ۆ��.(t�������w|�s��?�	��V[�;U$$�lXyp�J��I����R)����;(֢��h��	]vI^شiV(�3ISlT�j9 �_J�d(�7�Î�|�r�'}��W��[�k��dTƫ��Q*�p�6�3�4�9QV�.=�����V����'�A+��RT�ľ{���-Ƈ)�-��l�!Z��J^�>�3�	�ƹ��6t
{h�����L���ڤW����>��D�J�U4$zLr��K�7~�p�-g�}kb�6��C�W�B��}_��������+��K�ȓO��?�yx�g��/����?w�p��Vx��=w��Μ���T�e &x�+�o$-s�A�&�۲�~l����u��O����`g�
w�� ��Ea��B�4'M*����c�j՛2�E��@l�� �:v`�8���įeC�R
���
Ӏ�Z� �%hc4�QYJ�U_��^A/ږ�w*貥sj(�/�T��'��g!�j����a�Kb����D)��|��#-;���wl[K�Szs2>�o�͆��BZ��{�4F��پ�i�>'��5(�юQVwʷ����T2^,���]t1�����a��0�;Q�µ��y� �<�G���X���\J���#R���|�nxh���\��a�&�"�dtP�y8J"O��qv��Xz���i���rj^�0�MY�|6��V�'��]��y.jaL���v	��^u�9���/��^z_��,�}*Q�ë,�g�p�V�yٽ/���=���s���vn�����@�kP9���=�Z�u���l;�Q��J���`�kJ8�>;�q���&µl���:
Q�Nh�<����j������a,��XO\�|�0�X�^[*_�fCeգ�O��{�^��1r�����#�L�*=bh!W*w�qӨ��x���� u��Z��OʣS�2͛�kI_�闥z��Т��cE:2cƝ�kD��s�Ks�m��CX'��o86=��%������J���#n���7广^��#�)p�^��mxVX�[�U+N��U�{\=��"����+�T���5�9�Ҋ��{u���W���pn���UvްQq��D��5\�Mm[ua/_���� ������(<��s�Y��Sm�n���fx��w���w���m�C֘��w{*YP�%�Q}
�z?��7��=�(|�ҥ��ƯkUx�qE�O_�p����{�X�����`���2��Y� �6a�f#\|��%jII�����~��Szf�zC:�CV�����懾������vEb=#¦�b��Ou��ͦto�oD,)E<�$��[���d��t�HB� ��kMzrU4
[��@#@�<
'g�������4��`H��K�L�c�����(1�%)t��@C�2��X�S�\�,���߇�|�b݄��e*|e���P��ȋ�8 �?��`��	���%hE�?m���廰�p���{�[_�PKO<�C6�r&>w��ZA}iw	��{������࣏<�]ރ��ƱeㅹKZG@�������.���{Ϟ����Nx�_���~��hw�y�&����7f	[s�/�>�/�×.x<�0n7Z�=O�5/�S��.����B��-�oU�P�0�SZ�s�M����L^���yt��JH�Z�eg@ӱT8�x�����Q�=Mɔ�On�pr�a�(���7�m�����臭���iS0L�U I�qK*����[�ߙ:Ҝ�i�*�71��!�D\�i�ޢm�:��=+��/����
��"zFȽ�C�}���z�ꑋ���Ϥ��<�XF��P�c�s[��K��"��t�RYyG�(��Q.(�c���<_伡�q>�sI_�[�K�}�fI�xyfN}��F�xx�<�t?A�m�Zі�ʦ.��Z�:T�X���#�V��ݿ��փ�E�^���Mu�����0����\�&
�MK����,M9��.�u��&�>����ѩ�.C��o��;��)�C�g�A�_xk�{p�Ռ��Mo�׿�A0�W�0��i%�N0|��������O�,<�p���'+�!���mF	��M�y�"ጌMm�(SPFg��Q�,�B�v�$o׃�Ǆ��
]~������Iy��
T+�m04��l���Ȯ\�J�JGm����t��m1���6@���!�?7�G�ܧæ��5tR_jD?H'9������%�g�1�a����8�dY%��)�7~����]����Ò}���8Ju��=:���u�ĵ�M2cH���?�z���[�I:nf�R��T�@�7�o�=+JW�bȱ����sۑ�~1e2��G�/ɣd�auz���&�1�'a}�9���<8}�\�m�_�|�k�V���gV_g��)��u�i���B�)���c?�لM)U��$�1�U�m/\a_GLj��0���:0	h�'�,ݩꗮ�����^v����^�'l/\�8����5�3_�'������o��_�<� x��4�1vf=��c���8��E���;Ϟ��Ϟ�7}Ń�7�n?{s8��9�ˆ��������<p�m��oy���P�8��
.�<�j�7	Wu�<Է!n81B��U� i��g��F���ICQ��8�x�9@�-��F��:!_���p^i~2��}��Y��:��a� ������G�d���(�8S�E.��ǴϪ����&�ҟ�'p$�D��<p4AԊ2�8�iZ�B�O�W�$L9�z�<�jȥJaΓ���.ń��Nc����A�`�#\
$�!�ˍ#<pk��4A����G��*�~�D�Q�����V�Ϸ~���ne�U�4����(�h�jXT|��/�O��}�k�<�
�-��v�z�,jg@XFLg���~Y�kxro��3�އ�~������+���f����r����G�]#� M�����w��������{�1^��Y���\7ZW�Q�͵{��@���'�Ć�.��TZ�s �E���@���"����؎��ۋv,����'�a��g?Ĭ!�)��hE]����������|̒�ci!��;��iZ<�<[���Ɔ��q�@��O��h�@��0��� ��I:NWQH� ��d,Bt$.͉U��&)u�4�l`JٓiX{(��.����D�4b��$�Pt2*�Y�]L�\��3�}��k*��O|�	=S��+�K0��2^J�I2K��),���M�Ux\�Ć2`�N_��k}ji�j�
��v���=x�;��_���x���Bԫu����8j�׿�~����g����l�nW!��!��Q6T#X�y�&�M��ӍK��Yl�)���0XS]aD^��3"�O�V�z݄�� -�����,�m<�J��(��`�)���'h��&6N�)���f��B���,�/a������`�c���*�Lщ�8���\?��%��p۫<d�5���6��]�)]��c��.&[V1HpX��I���n��E#�w����͵C�R�����7|�d�(�!��4�M����=��&�t�����fLxkѹ�P=0�BL+@>��lp��Ӿ#U���Ĳ��J��5b&x�y�k��tuw	��x��M�sL�D|�!ug�nu������O�;����?
ϵ���f[n��jƧ�-b>{�a�����/^�O<{�����O�և�����mo��uk�����C ���*�k������~|�K�~�1�����S�o!!��5j�Iԑi�mQ�fS�)P(ۜH�P�"���C\:����M��z�7o���f3���IC%:7�.�*�bj�5���������[��8 PƎ�f����O�٘@��\�緒Gǫ��+d�S��kX,*N?m�O��Bt\(m���G{�@_�������V۸�Ǭ�
�ؑc�~X�L�3NȔ��m �vS[�>(��H��@��qc)��O�J���! ��ʶ#��s5a
�(,  ��IDAT'�?dc��߫୯���_�U��]�pc�����*�m���vZ����į�������;���N�Ж�.±��$	��eQ�ߖ3w��8����������(|����o~���uw����r�R�\+��^�[^������m���z�� Gc�6[q���*�#�ӄh���rJ���8�qq����2�����-:Ҁ�IɎ��/��מ��Q�Ć�K��~�mD3^��$���l�o4�3�u}bި�����;�u���S=��C�V�Q
jw_f�v=�=g��;D��R��.WH�i;$��2�G�O�
A����*�t P^��(v_�A^P�̻ܳR��#��ѨBuq:f��)ֿh��d
Z�冶\�r~�h�F��6����U&+���հH�T�4ۭ��g^�pۙ3��J$@�E�=�S8vZ��_�b������-��;
㣁x=%@G�Q���d�z�zY-�+tY�f���R�����챉/j��Hf�_���p�Yt\�x��Q���s}��=���ոƝ����jz0���X�8o�bØ�7uO�~~��)N�"�p�Q���I8*!�	V�g?�qC�b]�X��HF�#�V�6�H�^�PWe�A-�#�6:O�N�\�x�'��^W���CS�n�P�w� �KQ�0�h��� �1��s�4`��3�+n�u>ҍ�����o{�s�f4�&�A�s��khZ:��x�鯽��?_�W��|��i�u�]��kU)�U�1���Z�ٙAs������'�����O<?�?�:3�ff��K��XA�Y�;��Sg��3o��̿w�_���d1_\+k0�c43�v�q�z�'g�v�:5fFk0XD8����*�z
RE���%�u�xU��d�^v]u�|�����ڷ�",c�qPK_K���`��#�j��a������M��/�Z���1K��<p�\E�p,�k 
�2+И��k��ڴo�)缡�+��4������F<qآ�R3�x��v:HƋ;��	4����B�F���32�s1g����.�>c8�2��G��,=�\z/M=L����� ��GJ�ղY�b���������v+�[!�XF!����<�`�z�]i_�Ŀ�u����&<��
�Sg���-�����|�簉m
�U��:L�@��5�`��w�������?�������^����B�L�&����;�Û^�r�����uB�=��Q	�e�a�h�����c�MQ����G�(�m�ci<�,+vG1��<$`�&�s��*�_�-��X��Z�	
�\����:q"J���%?ͧ_��);��Ij]'\�]�pXu�9®r��*e�7�t���\�p=��,��0ڨ%��:�I�J:ie�����G?<	�J�i�������<�!g�A�v�	�1�֡�O�I��.�KU�ġ2�_���(jbq����6�zo��&�ے����}�9#�h6�!��,�v6^���9����!���@�D	m�
wO��N��n,��z�1�N��$�����U����^o-��jb㚴+bA&Fb��Un�$'xg�u���g����wd�D�´r�R�,�:��Ƕ��t<f�l��zs�=K��]e��'�fA�I∹���Q����NB64(�c��=��%,�w�Շ.��1��x��L��m�6ʞ��[-�q����g��=�6�Ũ�iW�M��ۊ)�?;���[�0�z�A���	�/�&�!��4q��b��������7~=�1kb�U�Bۇv`Va��<�<��w����������T����l�k���M���Rם�����گy���^XX��~~������?���F�$�O�'��Z���z��_�<��_��<sf�ڟ�a�3�Q�9+�=����	��I8��7�'���od���3�P(�ЭxF�/�5�8�q�:��O�˟4�7+m�����Y,����`��sJ�՜\��3Q���]��wy�I��z��0�:���xˀH�[Tc���� -RdlT�9dwN����4V6�r�X�y�@FwN
:�z���� e��nX:V�]��^�����`F��B
$�HHsI���ch:�,��힪�7�����|�����q@�f~r��RZı\��}gN���38h��z1_�N<��v��m��_z7��o~��m���+tԈ��uK�;���kKۈ�HKJ�O�"�����Á7؆'�^������Fم�����2��<=��kOVh�0�����*��~.�S8���w��*v������J`�2�Z����f�����k�C���#��<@�`RO��Y��r�F���i���q�V�d���Jg�%EgG����&h$CNW��q�(���1;�҅�\;�p�X08%N_����*�b(��g�2�aH��P�ǐ�D�,��J�����/��K�w�y�Ӿ��k�ȯJ�lt��;feݭ�Y�c=41�A��r��(��B˓��mL#"�W�ݽn�3��g}H�>+�6ݟ�ǥ�	�(jӴX;�Er� V0z����z5�L4�)y#D��P���ha{{+ƈ\*�V�r6����̷����<u�
Q74.��� @�|*ZN�������G,��i"�0���}�ب�XQ���r�C������jntc�y6"��+�/��W�V�:ø<-��8������c;%��=�5�JzKN��ї���߰�d�vL(�+��njc��Wɧ/N���gC��4�9��o�Xj�R��]Ȏ($ �NG�-��wl�Ј������LĐ�dX;�衙D�'��;ڜ	W�<d?e�b��hY��N&b(�`���.�>�w�&҃�?����*�i���d�ˣqk�qm�&1�@D]-�c�z����\�o�����7�
�..�46:r�5Z:[Ꮮz~�g~���/�՝��RAؘ�k@s�v
�d��6����[ ^F=�m^���칶���O>�e�[����}����_|�n�pI��t��3���+^��x������m<�\��aE����'�&���o�� �ݦ����>�:/�ǥ�	z��*��%*�St��ƈN�@]�Qw�s)�V�CI��&];b|��V��0́#LNd	�ZmTf�	�^X�{&8��ɢGj���A�?� ��}.\�M`d�������A	�M/�2'^����?!|�79��-�G���8�>� ��}�K��W���W��K�K�$�4|Q�7('kR�2���e��r��=��PA:|��l �#�(-W�d~.n�G*�>pn8�vy�9!���yn�3xvw	��}��>	Ϸ��=ˈ\t��?�T����9e;��*��Ћu�.��ކ?�z����9���M�g_�20�!"���͞?i�w�Ο��O�.}�-B�z6#j��K��_ba\�e��=;;]r��4��xD��<=)đ��GY`;����#R2���|B^0U`���ӈ�jBRC5�3lt.�d��|C��8p_��R����ڒAF~v r3����7Ҹ��R�����}�\ʝ�s(�\��y�<�O��[�N�~��36������v(�J�3���7ƴu_Y�����o1W�͵�� ��P���-��|�干��I��1C��/h6L�H?f頶ʄx`�	m]D�Oh2XDX��I��PO٤l+ɰ>���4ޟݷ��{����du8����q�p�)�6�����8e��b�I�T��>�Dg���@����� ҨfAl/��x�I��=ְ~��b�0,����&w��σ;��Gt��u�:�� h�x�2���/���]�9���gq�3s=Y�ަ�ٓ>�Y;���|�V��3��0�F��;CTbhM �3K�$t��>���#����Y�d���NF�'8����Ur�q��B����H��?��ߥ����%az�+蠔m}8���k�F�]����T�{���Hs�fLi�2JuN��B�c�b����'�z�Е~/aؾ:�0l��P«S�^I��?�ϕ�����/��+΁�8c��R>����e��(�q�|_�)�!u�3�u�l�dK&�h@X�N�$���5�:K�@�`�k�O~=�f�1��i�^��6�숷��$�	� Dg<jd���$X�Yr�vԂ^�����I���2��t�:��i�ɩF�T���Þ�\�5�Xm	�K�&��_��^xŽw����^L/9�N�k0�9��3���ԯ����no���M�n��_�k�aɺN�'�ذ����H����`��N�����?���?����+o���ǗѦ��'<)p�����W< �|��"l�u'W~]����Yn+�gr���#��Ķ�o��}'�TZg�BÞ�q/<���[	qx�`cz�0����:y��Ķi���,K�D��I2�w���&�1��!*����I�o���Mw�!���c6?7l��I;�>́�Wl�M�j`��Ƙ�f����咎)NA��!�\�yJ�.�!vF_%dG�W:�Ы��:*8�3�
��Zd.(c��9���ԙ1-
�Q51���ZQҘ�I�b��3]��8����,V��@��������4U����hsź���`|��w{a�W��B���X�o������w��?��|�a�5�f����<ƘEP0���y�O���	-6���Y���r b�[� �l��6��_؃�����[nm���ea(.3����ixi6>�'O�u�&x�V��j띌L��������!��
�{l|5��OB�씣�G�9#v�K��P15�]c,�:����3���G�3h�� ��[rBx�T�P2�8C��S�|�ˀ|��wVV��8�&�=%�^��˻�T�!�R*+s�գ��>�K�r���O�lP����|r�ʵsn�գo���)є�W.M陬W�}���{^F��a�T�[RT[V�̚Xfv예�;'h���!�tI���5���UUV	cd�Լrt�u(�K�,�F1r8��{��Y)#�c�!,Z�T@�ĤOh&d���s3�[%�j�!�8V����wJ�f�3�O�2���;A7��{c�f��#��ق�~�c��W�θ�(���X������m�c/\���ܟB讍�C�S�y�s�wH]g�a)그���T�ec��kQW�x���s�$�/׉á����TJn����}�ޙ���H臰&�aR�m�3-�0Ԟ�O���O����lg�N�P�Θ��3:y)2�����W��16�����,���n;���2~IW�����#�?�R�R�S�¾|��ۏ^Xz�+��}�Җ�/ջO�*�-+�b��	w O	Y�w���C�����,K]���QϜ*_Q?�s��)���u��4��X�M��G\���ϭ~�)�2=�@�p�5��#��m�ϣ�*<���zL��1W�Bpj�DCؗt4��<�>ڂguw�|�'�R���V�pļ�g�^�����+��?}����p�E]�q�2aƅ*br#�7T/ eG����+͕�7�P5����=������x������w���f��#�I�!<j�<x�]p�Ԏ�Dk�y��[��񴒸N�m�t&٥�/��w�\�L�^��?�!Eb%�Z�f�8DT�k$I�o�c� $n|ȭs�#�d����P��Xq�<��I���c$#x�\���*��KӘ�㨋��X�#��Ra�+T���f����l�7�σ'�0D�3����i�Ճ�L�U���f�{�o������8�T�)9{�*"�ʤ5�i�/�hX�ȃ�uW�ɿq�!왱��	-EZ�-�i_�X� ��%���G��W��^��%�c�c|A�K��� ������V�o�s�Z�?�j�F�R�P��:FC��^c�������; �%z�,<`�vM�n0��'�w�c�Co�V��\;���{�n������=���wܰ�䎹��"��i$����!p��`f��oWPh�6T%�I,rA ���34}b��0
�/ϙ�d8>}���Z����K�d��3Vڤ,���	��2��rt��得��~��I����+M3Ds����)uOey��R�z��q����X��N�qJ=J�Tޘ8�Y:�}(SaܜJy})^����M��*�d"[�gm��+��R,��efێ�0i2 Rx��+4������C�,��%?'��M���*�?jef��]��r����--�;N�Aě+���q�$y�l�٢�f�M�&=��I��u�W��B4w�qW�o��s���}���_�	��Qot�N_�9��[烟�Bh-B�<������KzC_*_�}�mP��v����~�Q;<:�O�e)���7U�5-���·X�'#��zx���:��z�:V)�A?��9�0�������:����3ê|{Y.�����eC6W�>[j�U1l�+����c�S#�w��Rߥ���ֿ�ߎ�K4���������W��ˏ�?C4�^/!,ٰ�ߨ�"̩�Vzxa�ږ��A�]��z�j��F`!�[h�V䪢d:,U=�e��LEiY�N&$�m�'���"����G�(1.�O�SANձBtZ��d�5�RO9�I���p���#xCE#��(�;�,�r��{�x�iX�T`��K�4���۶.3_Ve� v�f��>h�v���x�q��⮈iڼ�z��;������7�k��|5�;��+�+J��go��n}|�G��Z�Cע�9��Pg$�	&sњBcI"���G�t��z�*Zᨛ�)9�$�,�p,��E��'�S:�r�M����#�Dm��m�uc��'� �����t3 k�*��8Uf�z���J�h-q��U>��;q���RzL+�+�_Nc�BWh���b��r�Q0'��O�;:�!.���C�-���%%>d�������@��f�D�6�<�Ֆ"�|D�ğl�5t�,��\߀�8ǘn�4,J�-��ah���\1�Z� d����_.�{�BħM��:�Y-�ß�|�`OW�K�mp����82����*# ���R�-t��-�Q^-�rFH��[s����|��n�>�hd��9^�<�� �u�� �\�U�[c�G�;)�Zё�'sF�a� �l��l#M,���@���t��l>�m��]rP|x3!�7�H^2B=K?��祹S2���5�c�i�ra��n�Ci�g9�]��U2���l�c�H:KF�\]ruO��b�q3uN���%\Jϥ�,X�*׈�5���-�L�l�N������xٔN�Jez]��F �}͟�f���M�|6ğ���5{���	\��O��Q%�nf�,d$��U׊ze���+�[6�Y�O�B�NP���.��{#�����wk�\���я�k^���B<Bي�4P?3������)x��~����|�;�צ��`JǼ���1K��eq^��
uC�2��H���b��&u&�)Qp��b�p�#�:��ζ�c��}�O�Z�X�hH��ߕ��
؃&��iK]���Ҷ9��a��31�b�Ma�!�9Î�gH���xCa�5�]�c�]��m�/�G�w��i>+�c�֤[rs[���LYw�x�n��-u�yY�J�Yo���o�ɤ���s>ň�{�[����I� �S�A�w�(~�\�������cs�S�Dq�;��ݟ^�� �N���S�	}�+�r\Խ6��gv���g��'�+�V�g/� ��g��6���c�*���x��	5�  �7��T5\��u,K�n��g����._������W~�=m>�p
��GZõ�;�^|ǋ�y�_�̆u+�f��R}k|�NDhC�KM��G���2=>M.� ��s�V[�`oi���ե�Fې��q�xjH��t����Je[��&��*�"1G���0�:��w�eM>���p?H�´��U%ɫ\|����qW�xCWϱ'6ҁ��z��c�.��ݲ�2sWJ�����;+���
�`0�[��ݨi}"C�
��2��d$\P���@"B��U"�-����3�d��hL��tV�����+���m�b;�1=�ޑְ�A�{�~c�(6� �9E)����X۠�SƝd��p��s��-7��ut���V�)	�d�]��K���W�̝�E�|A��u.}%@6LE��ĺ�^
�]ݜ�����6��|������S��e�:���:I�q��kx���y�	29Fqd`뤳�F����؉��c85ѫ���� �ʑ�!�'=GZ��#8u�F i��8n���Qm7�7�c������+{��G <1���@^kr/�Īq�
�]�	�� ¥��,���<�'�eku���ra2�d@��d���89#g��s�C�~�6��i��8�:��U�z���4h�=�+�Lq��QTn�Ǝ�>z���E
�tZ����0�R_�+ߡ8y�����K ઃR����0Ļr�|֥�����_@����k(4З����
�h"���ԊO�=^7��U6��@��ψ�KkD�*u1�M|��,��aC�lF*u<�'}_�k&mХ\ާOÿ����k�������]��R�;ޚ��54�����$��_�%�R��yM�3F�LH�m,H,z��hN���&Վ�XҟӓJP�6����w(��w��`k��Iu5]�U���9CHf�n#�3�ɹ!���4cFቾ8�Lo��0�T<�䔱�4���'�<�t��[��:E�=���wct��Y��)/�Si=ցU��E}����ߖ��9�_���K�_�Ї6�G��@o�r1���Ԟ ?���k��mn���L_ga�M�58��B:�ce46Ը,�zy��k|"p	ffMO�J���M�(����&n�Ř�5��ҩ_jp���_ݩ�O ���V�П_�\�Qz�A2���{ঝ��/�Cw���V��������m��ϫ�	�������<[��&�7��)���p]�	��TS���wDߒ����>O=��Hd�Rj��w��9<x�6h{m�[ 1_�cT���K#��[�&RU�����4~Ř(����ݞ����o�$Xw#:W��*�b�+�3}r�BZ?(�R|#���"Շ�p���ڏ%��3�4-�[�,F�un�
c��i����o� ����7فw�w3N���r�5: O`�7��b��tJG�@JI��A �)1:G_%N*UUT���w[L
�oEM��dRd#�'��1�2W<_g��XV�S��Rű�q�RV�9�&�-���H!H��GԎq��=��sEf+�Db�,X�ՀT7�$/�SM�u���ͅ��<���=�!qܧu���{�p�U��|i<��{�歴�,�Dp`i�����׭ȶ�_���.½�K�x֞���]��O|��UA݂����>�w�ٖ��z�tf�p�Rl47�g�5����P�3P����L��p��]=�bTGF���`�q�0X`�@�lp�쏛v31H%y�hÉ�|Y!G$77����|	aF�1�ycf(sW4�d�,%�i����%`��`�԰�YH+�Q2��}��1a��a]y�`S�(�>��>�a�4;&KYR�S9�h� \,/�;�N{Qd%�`t(�UX�͇�Y���\�nrL�F��I#�	� �?�!]����R߯����:�"�e���Z�#��q��;E ��Q�V9���������vb�����)���h �!�l�F0,�Ҍ�W&��'hGn�����B���3-v�?�������^�
ةf��S����:�nU�G>���~��s���>��A�	v�
��F��2uH)�#�{�p���N��\ɠ���R�:�3�G��z>�2�s�P�[���ۇΨ��;�C$�x��`0?��g�Rb��݉7����v.�7uL�pIg!��8� �3�S�yzA)���"ǔ|��SyW߻�NNON����Uu�1z�`�Q� ������,����s��+�a=�f���y\���pDB���S�h��O��wahf��"�"�C�6ux�\�v����[��l�@��s�m]�?*?��N_,U�;\�3@��� }�����i��Z�$�e��z����V<�ܯQX�6I@��ҕK�hv�j��b��
���z�H_hߥ�8��K�:��m�U�g��~����Y���s���_|��fw|H[X�׋b�zͣm�{�<u��לb%��� �ޡS�jGn`/�g�tu����;6���4@�1�I�,��Mb�1Mev�%Ҁ��� �'���ٽ�fxN�1jsX&���oE%Ǐ��:l�\Q�l�:cd����@bW�ڤ��/�n�q:5V8?�MA��~Y0ف⭪��+���@y뺆��f�������-�bSE!������Ou������&�dH�	�L�Ⱥ{�J'���I�Bn��_��穡��ؤ��	��zЍ���D�j��
'p$ƺh�F-�����\����/�ٟH㳗�-'`�Ѹl�.^��ϱp!w}JU#!zr�A��m��P~"�W��d�Nn����d�(q'=��3�\�#���KQ_��;[[p۹�P]�ʧǐ<�~���� "'$t����Q/�Q�����ި���W��X�=����<�tZ�\��K=Ⱥ��^�E�Q���1u=J=?�	@.v��x�͘�;���\���$�P���0��ҧ�S�Csq��`iт�O�cU��1Vӿ�A'�����b��I3�W��vS��Ss��g�' Z"�#0/`$yEa�F4��!L�����P�P��U#�ՂY����G�J�
:�O�7�`�]�S8�i����9��]��w�,|��_o���@�l�[5쵊�S���_��û~�7�W�;s�Y��o�-��SE��e�TsG�V�cc8��i�M��Si��,eݔyt�%:��*��p�<`!,RTl[�����	y�� �G59��a�ƀb�ɤ�u	���rX/�d�����pxa]:F�x,��nl�k c꓎a�pB1��y����!��uX��i�:
���@Ku�χ,��Q
����
��f���^P��'"}jäR=�pZH�k,V���&��ē:���Q�6����O$���<���s��@n�P~���{�������_���F�YK�#���Mư��Oe�5'�"u�/��4�ҿ�Ҧy��g��U�F�T��M�}�g�����H69�Sӓu+����d\��
�J��I%���R]i�T����u�N٨#"���D��G��%�dC�;t�^4����n���=P���*a
���=o�[��cBh��C�R��8�-S@'�`Ћ���yX;z��h4��<$�������snY5�I�ʈ�ʕ�P�N�u=��;����M���aQ�ӅVE�#�V���A��|���w��m��kB*)Ȣ�EaRF�'��?�g�����M�v v-'�s��6j��vu�*\�r���vy�	q��>y#4O���xk۰s�E��xZ�o���Uw�5b8�����8�`�;�ݒ�N+�)P�o�`�I�J��B:µ�^*���V�O@4"� ��dxk�8d�)3��e���л�a �QP0Ɔâ3̉aA��p��G�ߜ��X�IN��'E���8V@B_5I��g��4ު������
��%|xT��t,�8\�)����� 0�@9�ZH��SH�"���et�Xy8lR���R&�?�z-��x -�2��M(�#U���<��"Ө{��N'L'����밡xX�������gl���NiA���C}�)�����s����U�|�:�AƝ��t:ՙxj��O��oû~�w�Uw�εz��f	O���.?��^��N�i�oy=���jC���Ő�&�-�Ք�,�A%���y
�*��Og���^+��M)Q'�W4�]�3!�#y��������F��D����=�h��y� �(��v��62Hw��M�OGV��ª��������1A&}�\�)�|ٱ;X����vR�һ�9��5�.~Q�����	�����_'A�>�X�1��e�B�6���C�����'U�N��p�c�~P\(���bL�<m���U�סX��^�"����>s�+�?�5Z�̝*�)�j8����`w[~X��,�.A��.^��Ţ�Z{��*��Wŵ,�"��e�<[O����)5�7ֈ��o�mZ����"<�5�t���j����.F�i��:������)J�=L:��ưI��]F�ج{te�fJ�56y.�`Po��q���m�]�9�����)@���c䍒Ѣ��t)���ϩ����8F��ScV�������Fe�\�<8} B
Iڤ�X�xr��ѹ߉��0V%��\:Y_T�Qpl
r�I�	�,o���\!�ry�P������uiZH�^x�ݲ�cٲ��%�#FU<
J#�(`	�JD�����y����8��._��Ta~D~ .�����υ�g�Dǩx���N6?���#�����0�#Px�H� ��ztE�F���� ��"��[*� x���S�L�e:�2RF�W��nXi��W��0��@�b5����u���*uyp��]�|�����w!�;�f�tC�3B�%9��G�L7qq������'p����������"�.F�>21�����SF6i)n�����L擸��T[�D�P���(硟�}"M`K/�˧.V��*"&u���4ϣd�Z5�Zė����[6H�94�M�ϣ�e���i��F�&���� ����(k,m���=���jl9��h<�M���DL\��w�I��r�^�Uܾ4">���
��oh��:E}N����7�|�mj{��He��<�<��r{�Q��U��]*���vF�y��ym��!앴DLq\�|Du�rc1�����?��ɢ_��-Ѵ�c����G6Is ������%EA��i�*5�w��Ako$���q|@;���})�)��pl{��t��NT�{S�A6�X&�ða��t6�B� �&��[)�ה���0r8B9Ca�!;\I���R'���@��ZfP�~��|���3���<���0Ȳli�/���>K�yc��|-�[���@�����u�)�q�9̡�Q�,�	��8@q�U�l�8V䌵�{��aP�e1?�Z܏T����]�Fԅ��U�h�'�����txkp]Ž����R��^�z%\9���L�?��­�4��X�Y�����UU�<��E���O��}�F����j��ޕk,��KU��U��щ�%@Ϫ@��O�8'k�p�o���3�	���Gʾ�L蔤���Hlȝ~�u�K7|]a�~z|�k�Xg�r�ɱ���I;�:�,&��2�J�izƋ�D[GҼZ���_';p�=1R��t4��:y��O�\�%Iw
��C�Kz~����xa�v�)�1A�^yM�-�삲�{~�gC������؝����\��Y���2��C�;�@�>���R=:��d(�'/6/�Fb�'lP!�'F�����$«�(.M��Ut�?��7`�p�M?�d�+����s�hA��O�Ђ�������2���
v�۰���x�K�-���!ka�ĦN�0��Q����D��8=ۆʓYqy�W�*�z@V��ނ�^�ۨ�P<�XC�2Ô�z��;�^ �Ԇ�0ep!����o�2:32oK�c�����k��2�X��$�4�l���$�e"p�hp����U�.���-��r{P��ֹ@EE$�%�G��A��H�������#vO�5x5Ėu�@���D�HC�����9	��9.ހO�?ɓ��W��!"�CB"d��c�FRLf�tP���+�N���Z�
��	��
EhR�g�7⒴N���p��>+A��H�ԃ���qJ�Ђ���N��8�4Mh<��K������� ,�)6H<�����m�C�34�⸥���W)��ͬ���C��j�!�SC֭;��D�F`���id!��\< Ƣ	68.1�~
9�T��6N@��##>p�������R�H�:gB��ɹ�0)Z���4J�,�2�L���Q	ҋ#L�-��<��44ǰ�Jn-HTD�Ӌ[%�0��s��8�j�ꙿ��;v4��W�B�0F�i�U,6�(����h�)/��>�y���L�>5�/�%�w��t�2�卍&�D�`���8���Sem:WA��BG�iˈx��N��#ƈ�wU�Y�uM��Fl`[W�-<ޭ��d�	�R�s�9�q�6�7J�2�tb�2>���-�VX !��`Ƽ?*cX���Ҕ��1y(�cG��'~6V���m�
��/h�@�s���Ϥ,�?����K~7�וT�l#ª����S�Z��1���p�Ǫ�D����]��F!�j��TaQFh����H���֨Ef|���| �:+��q��"l��6x�H��!O�s�I۲�zS�����6��"�k�h(Tr.��f ��Cp��
�b���j�@�m&@�#	�Z�0�m��fJN#�b�H��Dh��D�3R��rktd@:�%]?���S����m�{-�ڭ������<ןL�Noi<��󪂚��ByZa{F�}.� �p��K@�me>x>��`vb[P�8Rl�_K�b�l�����@2�|]�9�8���xFBZ�ZN����������25��pq����*F�6�� t��� �M�L	9焃�AR^��Z�x���pg[�Ox=��n�Aښxڿ�3p}��v�1ǔ]v��'p @K�߻���vz�<V�`,�u�p�F�N�>E�����Aw��p�vjL�
��L,�AK�V�� �V�)��ç�0~:\=�*�7ܟ9���ڊi�z�-Ң��"��R�����F�L�L�}���	c4�at�� �{-�����\D�P��xa�A��Zὼ�F�6w�DnUB��J"H+t$0o��b��R���k��t�L[�;jlIy!���n]����e�.�w�;�Xp�N�+���a��0d02��@���<L��a\��Ib%c;�[@@������m7�s���U%3-��0���@���1,��:k�*�B9�N���P֣f���<�C�c�E��9l,#�*����<ᩓ �;ɨ�i��l#4ި��xqv'}��a!�����)��}l�z�ѡ3.����R�KBO
)]/��5��J�t���b6��z���qT��1�Ht�M�24@��:/S�&96=���JI�g��q�yO����"}1�vzWy�2���4]+�E�Y<5�vޢ�D�R�4�� øСq�5�*u8��n��5����+��T�б@`���6hBg�N֛ҨqYj5�2�	��N��HGv��&mKs�X;Љ^���U��x��)��^�L����)�<o<��!� z=t�Ȇ�VI�0z�IVC ��ꬳ���~&c�b�U�4�l�F�a�P>K{�O$�{ȡ�M�"%YZN�F�!�%�l��ݯ�tJw��;
Ǔ�Vy�O!b��O�J�GL�pa�G��
�7!��tOB6$˶QFH��56�����RL D9����S!;�����8�E.{`F*O�a��Ҍ$�`�>��6��;(`�y����������7D\��N�8�G��d�ݥ�⺒�5l&OY���|�T3xv��1�`�������ǳ֤�o�6�[�i?o<}б!���{��������*�3��*��׭!59o�n���$[�W΋l�D�E�oS�T`��=:�5�hn��_�8l��s�t�k)B�'�MlY�V�X��l�����l��12Lr�0��g�\r�H��ޣ�K���KN��8�`r�4S���<�n��������g
0P`I5.�P���d�\%t �C
��ۦ"Q*"yܓwP4A0R�x�� ��h4��}ބ{�}�*x��7�M�ذyϴ��J�7�Fu�蠂FS��|�w�pf�?K�R$�S���+�.&��$�?��qP!����e�����oi�޲��f4�r��>���l���+ �n�x��-Z8�32�OH�>W�\���H�� ~��Pc�F��d��܈�Q���c��� >\O����ʜ`��}�r�Z�*���s�e�|&��>�W��4.��H�'pd�+p��t���xm�IS�M��렩1aH7];%��@~Ou�L��܇�+�~��!f��(�t�Mb�w��,\y(�;�F�y9�m���eAE�o�p�;�2�<���T|��p2�@EvUmQ���m$�l�&���[�r a?I�]HQW?��B� r�É�L,WIc���J�=d�N�?�G��jћ���1ܼDA�F1�V��r8
�����N��	���
Sd�[�-��ć��N�z�Q�N�Ȑ�\V���Q�J`_Y[�?�LCxQ���z� ��(2	�3i��r��X�>0w(���H±���}k�ġ�х���W�n���;՟7��?E�M�V0��3x��%�V1�#��Du+�o���-7��[O���aW�d㯄c�X� #087�ޜm�#�W�����"Λ�x�ll��=��E��W��ե�Ӹcb{٦R�^4��<zR�Zf�#l'��Uy=�ۚ��i`gy��T��:��s,ik8&{�8-�O�8l&:�ML�
�8�Ӻ��Y��&�����IV���D(��1�)y��i$��zkk+z�4�tV~�����U�fR� `{��y����i�Wg��,7:�`ĜU��t:)�d��!LQ�,?'����(���k�q �l��g�쁻��������XK<߄c��Z���Y?��ִ�/7��|��l�2�����F��V��w�P��6^;��t�ht��!gl�X�pe�i ���P���]��rs������G�΁c��K{.?�{�!�w�t�1]n�
%�5Qc�b�e;�e3i>�	���}���B�[��9�m4X_�-��D�G��N@#�Q�Ɯt�I8��z�t�RCm���i3����|6�;*�X�$nȝ٧Snb'�N7,��R�v[�ޓ�L�%�z�ƚ���Ju)Q��S�NO ���a�G�鴞��/\tg�0���F��������ʅ�g��>cBY�:H��,�ѸhMG��J��g�T��b�Lj>� 2�8eg�t�U�V�[Ǵ�6Z�N�`bX�߈�%��&O���8b`��z��p�0'�$��e���j�.lk'�؆��Kai��Z��)�g\VB�Aw�峓3L�u�W6yͨ���x���"���ů'�b|4�J�B\��'F,ݢ�+����N�7�:ݭ�0�< ��,8�Ƶ�Oզ��ɋW��b����􎈇r:���u�[Μ�;���'�~��	��m�x�b�	��L��.�N�t��c��֋̖�oi�S3��[���"l���=�ki�Yt������e�:�8����B7�\_Q�+R��% ~.�5��(�@&ˌɥB΄���t�A�� �'�����g!y�4�NZ���&�_�M�¡mN�ӯp�ʒ�k�VܒÜp��0�u��i��;�8�	{{{���l(�8��O�h�b�:
����n�����PHe7�2� �c���i��0jk3�>9I<��$)q,'B���B,RN��#=�l��L�����9e�����p�Πu��2����1*�^��@�\�;�DxN߰���7��,<�܅���`���PU�u���{��\Z�y�����N� c�h��H�F%>E�P������,aق�3-�/��ΐ�]�����`�^�
.^�
W�|���&��^z�}��Eݩʇ��PA#���[�]9��2����y�k��\K�\�n��_U���Okd �P6� d�Dẗ́u���x�]�|�&��*+{��0T���g�}S�d	��,��LȎ=ulȃylN��.�kl����\�M*Fc�!=%.uD^g8H9r�*��y6����}fΠ���'�B�Đ�ǰ0�؃�-i�L�	��^�R��h���x�3�Ȁ�V*��,��L�ch��cʥ2!���α��C�%�tոa�Ly�ry�<����V&ƋZV���
v
ҐN��F�G�p�s�1�!.�qt���LO#�,Xa14y���9i�n.��&F��\�q�b?��Cә�/���D���&��^�Qj�RA���k(Q�a�bR]�8��0��q����������\8����r�`99X2~��sL��r6�kն�돴S�%���W��S���P曶un����`��X�eI�^Z����t�,'a3堵�R��pX��0�����!�}�.�	۰St�+����n>񋉅Yȵ��I�M_������9 8��8���Ï���f�S���71]�u����&���N� 
�;�c��eO\��K�`��,bt>������⮻��}�iX��)���
i3�$Y�̩DkEo��6��:�ba��s���ΰ.ܠ�!�m�m��x�ټ;�|���I:��F}�����<�h��0k`:%���-�L�W���!l\��a�93��D�u��k"�a �gyM��"�F��Ar�lS،i�tL��8$�4�gs�j�2�u"So���1�=�,�v�~{{�+�ł޻�:��g491��Ħ�W1m�Z����2&�&�5�~L���L���v�莞�(#{4)���B07�̀�H:E���)}�l'��~>�����G���L+����c�y/L����B�V�{עY����G�x
��f0[[`���*��mі�ʻ��Ϟ�ǟ��b�r�v���ij����V(	�Ȕ�よ#�������m7��{o���=�qLJ�e�/�xz��g��Գ:
��N 8�-�1
g�v��8/�f����IԢi4	6�?A
�u<��j��+ +���}�P;B8�������5p�!8�[�yf��j؄�B:�r����K_2���gW1�&����~�X��̵iĦ���RcW��Ӿ�-������}�1F	I���)���z�}�L�[���߲�г���1%]wLF��YD}6ϗ�ET�J�I�t�ŵtaHŊXb����1�4��X��P'&�0�G� ���K�)*
��yC�-_��&D�m/�q��uIc��$M�6��6W�BR>�y>��mgԇ�M@��G���}��y�I��pH3�����<B��s�I�U*����U��D��ޝ�M������I��f�ac�??�*�Nܴ^o���ҝ�7E�9H�֢���ɻ�Ԑ3F��Q
�q��S��}�O/(�ѧ+��.��r���S��ͦ�Y�7���IN7��ا|�/$$<������K(��hL��J���@H;�k�h�>��'�M㓜MB�$P�(��1`��1��VEm������u�d�m[҃i~��U�:5�6��:�/z�;F���a��c��xʝ��,����,���
�q;^���~�鼂/]�Ͼp	n�>ff�wG�6Y:U������W?p?���D�o���-VD>�Q�b���5&�-�����v���݃W���p��,���,:jHK:F�,��g��=�ӝ X�Bx��}c�P#)����?=��X�O%��!���:H�k)�H�R����JZ\��N�9�nj�.ɧ!;j_�ӂk���д��M1~�xg%�K�?!nq�B-�<�}"�sm"��l6�л���k��ZɁ�bFu��O�a{��2��l2`˥ëT.]�����R ������������΍!FU6!�n��8ߎ)SO�}�-`Q4�����H(�8�4#�Fvb7��,�I�&@� AC<Z�D�;���.�e�7�kS��� ,6,V�a���ҷ�s�0�?{o�l�q�����{� b�8�#D��H)E������/�ˎ#'_T�r*����R�$��I�r�]��-+�hRI�	�&E�E� 	�����}w8���{��{��t���{�ٻ�ի�5��X�q[�3�_k�:^��C�?h��2��������=�_}�v��C�`bf���ϔ0L���Z�_�xvD9m���^��6�:iL�yl�SL[(����7�g�MɁk�wE����(c.:v���i�u4X"�)�-�"�Q]���%Md~��<0Z���E���mYGū�\�V/��<�ϋ.��}Q�-;^���E`�cm=:y�w��9����r���J��i�6��SB�з�M����4O�9]�b�Yu}��5}�U�~�(Sh���u�����@#�ng8_�y����,����g����P�;�p�">9�t��
y%I��J�cvȻkJw�k����Wz��l�{~���7��HHcЉ��.����4�%�鉉=)n��I�d�ϩ�y�L���.{�#�cTP�P2�����Ӌ�9�4V'2z�Z[u�B�;��^t&.{F��f]d�3�/�������R��r%�ڶ�n}<��|�4}����}�W�3s�F_�%�fL�J|EI&:o�%ˋ|�.�kL~=�Pf�L�e�=��@:h����nBi=Y��P�Ý5�h^��1�P�!|�/�kCb��l"�O2n���Ō�n�1��"#�г�웳�d�䃻bd�X.�!q������8Ry��Av��$|g�"|;J���b�
���'�P�U����J�o$��[�z��޽6�N�u�;;I]�z�gfE����mtb�i�2��p�-8�T~?��w�$\a�Q�:5����=��+�L'Ѷ�]���Q�귒&;=\�� g��[�Wu�>m�!Y^"~M����S�ֲ��
���l4K�}e/��p��%�Z�l�Oqpt�>~�>G�K��U���XҁC_O���L��"tXd��i�wtt$� 2�D�&��PK)�����ƽ_F	�
�$���o�� 1��C�=^	��|�+F��l�4JHt�+�|#���vM�Bߴ��ק����E�eN���N­*���s{=�!m��?�,m����-�r�'09<���R��}wzږ�mh�S0��ɩ�ڇ���a��o�5��vS��{� C �������t<?ő�����7�����Z���&��Axֶ���vd��Z8���x#���|��b�[B���=�8	� C��#ǢD���=��%����(
�i��r���_���[���,	��.%K�����s������ӗ������Gx�����W���fVU�^�W�ƿ���2��������?3�����P|�\�nAi�yS'?2Z��
%��#�_2�q-6��Q�9��[���#�\_�`�R�lAˤ�+���BC? ���ajyZ��S�Z6RyK�3ϕ,M�Z�|%9ѓ��>K�ضJ�]y�3�z��{z�d��d�k-�5��o�����[�?��y.;̙B.,��x�1�ʘ2���}e����em3\�us�9k� ��������-��]�7�Q�yu0o�:U`^C�}�R�cL<b�7zϓv;� �!� j.��^����_�ؒ��#DC�
(�Ä�eG ��Ӥ�f���o�ݜ�k&��ܤ2������U�C�/�c�]�(�[��7��ڍ�$����!\OHV��i������g��|���'�����ti#Ru�D�Fu��s'�����=����������x�q���}wt�<������.�v�+a����{�?�
�.G��y=m��,{��$������fD#�B�8�q�<t����/���6�wn�p��v�-�}¿���v� �u��;�.J�8DFs +t�$�NN����A�p'''x����E�((ʖ�Q����96_��e��V�:\*�_/��j4ֱ �2ON)X$�'�.�*y���M����Y�y�?��bM�q褰97r:3<��f�J��Q:�u��Ҽ��B�L�G�дD��"lT�t��	�;��A���$�tԖ��19����o���*Oῒ�Y�D&��h��{�፟�<y�AƊ�%\���"�g"�h�>������㮃}����U"7分�0y�c��b����eX�7�L��0gT�b��4�o5�ew���3�b~��h�*�s��(
�	کoL�qz������x(��
�{�"�p����������l��C�UN��kǘ���x�����E��iiWɻ�!ы�����Nd� �p�[>��*E=�־��A�
����ot�90C*?s~�y�!,�炨h%f�UM�ǘP�`��N����	��%���2���:@o�b���W]�rQ��@�d\��4Jv5<��u�tl;t��&�\)��2��o�����D���t����r� �U�ȼ����C�i�Ծ�ͽ��U��u�����`�����(~���pfP��m�E��X9�Jٷ"��Qd�F�y����K�Y2�lb�N{�l>Z/u���м�پ��;��l:a�t���g�>��y�4��o����d�.1 ��[�EzؙI�՗���{�U�M'�q�4h�<l`4��Kľ���I��zj?���}>��A*�����t���]c�O�W'N�3�a7�]���a�p�.� DG�P�^]ï��ᷟ�������脝�� )��̅�I�4����|�>x��@��/,&�\G��/_�O��2L����)M�{,��@I��:d��1e6C��_��@�4�t��آ����������x��V�ޢ�P}�;�����O�s�XK��Z�r�H͗0��xzH^�;��
���%����M�V���߇��S4dz�����#����d�������+�1&-��C��T�7J��تN�O��o~�i�7 ����d�\�}@���.�}�Ս��3
9��1�Nt�'����H��̋�ɩ�}t��짳��L$kEh~�x�ٽw�	��������c;��P��LNN[Fb��8j����y�2!���vA������4r���h��	f..m�Y�)a����.�����>�h�����<t·Y�9:�p�z\��Ne��7�����C��y�x�I(���m�o��"4-]j8b�qW�pwǒ#C�գj^*Ŗ�T�;��*���饆ҭb���lh�S5�Xn����+��B�2��ʰ4i�N7�8ݐ M��;k�������9�
�u16c�'q�«T�~>�T[�*�H}��*��S��9A�+gz�S�i{��<Ee	�|���w^yCP�cc���;4v�̗yi�ց�PXoJ��o0$�0/	2��~��P��>2?���>X'��({�`�\
�[�����Wr�Z�Z��J�ZGܘ_j�w)�懔"�A�*Y�w̯�^=
̰�ŀ>�*ܳ⤍L�J0*\����y�B���恧J�Iq�j-��F�S8鳸TX^�1�h�M�=��欌�*K���<�^9Vv)�c�3Wxg#pر�Q��&�B��\X�ǭ��sv-Y����3LH۞�����S�GV�7��΀���ez�J�Up�u���{ʝb�g�g�	��w�it�r|^�<y���"rK�96,R_�>�����k����T3/���q|�x�!y�k��c�m��b��t���ﲝM�6F�����̘1���5� �y��)�]���>ȥm'���1��:�Đ,OkZ!��x�~���ϗ~�q��Kffڃ^��"����u�J���p��͓^KOL?�'����{U��;��o~���p�4FԘN����j�����a8l{����	���'�7o¬]kN�
�L*�����YZ��Dw�X��1ZO��x���7�7^��l���)�ګ� �h�W��<ͩ��y�;�r���m0�ӧH �Y�橗^��n��/���WY_�N��Z��#ou���"��I '%}��Ց�T�h����Q��p&L|��b�񪚞����{?o�����e��l�ǈL�����I�^̴��6�	�����)
7�xJ���d3Ԥ�1��B������a�Ax2����]��C՗y+�W�x���ʕ�jC�W3Qf*�ߠr�]��p 7o�M��E�U� ҄���1�Eu 
��<�UC�n���.|��y�XpIHz�\�Ð�P��]\ֆ��_pSw%̲�Y!�?A}�j�2�sP�'�A.-���$�)��Y����`�]m�\���I�k�����q�=�cm!W����,��-��̊g�K�]'�f�)rX���75�B*杢�j�K��~��> �ڣp}6�ׯ�9\i��2}����J)U��1$pU��1|��?w^��Ea��7j`f�i���W���c��)LZ��q^�H%-&�Si�*����� c��$���Sz��\]l�8��fsQ�2�\�S��ٸ���oH$�1�$�s�΅�Y0���R�b۫kNoؤ"�T�V�m��e`��tѼc�]敹��R�e�c����:x��W}um�G�׮\pl���UF�2�9	����3��}6^��CQ滤���J��n��/h�q��}�o͒?�a�\�]�Z����e9-m���au��I�^~*V�d�}�k'#)U�jGy�:�}�L��4�$�te&���H
Ar|	թ4J���jR��`F�זER2��P+�48�Y}�͓�tJ�Q�	����˗������]cΛ_�RU���]G�$���MP�<:����%
ίeϋ>}�T��k�k_9}<�X~XUnS��x�~]�0��3�Ue����'��h�ߞ�in��vގg; 8��xE�6���mK����'�#�F:&s�]s,chkfL	���"yD��2�K��'�h,v3�I49n���N
�� p���}oyc�]X��W�[b�mM�� D�H�:g�*��ж2;�+��NZ�Ј�I�@#?@��1	�<��`>�η�_�
̦Sh�&i*�����S0�6�}L�$.��T�+��-�>�~�(!\F�ոHe�p����O>7*���CtHק��W��>�r`	D���"�gf$���u^9�Ӧ����8���
3r�����%��%�jȞ}V�ۼ4^s����ב�\����M�^�V�Df��z$�^X,�s�v�w�T�L��M����0W��^C��cvz��GxF ����U�}� �6Ԍ����4��\�߹�!���	�����3)5���ʙ������_Q�	%:H=�q3fB�n���8=
�%��VL���,Ŧ�a���F(�F�>/�;���|𠌮�3�8�Ypހ��/,NN�Eg�&)���������CS{j"+�H<<��S���B�a	N-]�j��?U�.W1�$�O,y��U�9��w��[f�v����s�Ԯ
��(�h1͜�M��>�����j��2�ؔ�նN��6�c����4i��(D&@�4��o9���$3�^t���!�446ϲi��Fo=m�STn�\|��b#��@��yInnw���Ι��s����P�S�ҊZ���3C�Q��p��f��~�_���deF%*%���g��6��b�	�����i�x�����ξ7�wvn�1�/
G��(�,~r8D$O�}h�$(<�@�%��(31-�����N���@rG��0R�H�Rd���ZFP�*bj��(�3HK�cs���&A���a�g_�Z�4r�"�J���R�6�6	g��u��&S��{nG(���e(����Y��>��aMݛvؖ��F�����&|5�%k����\���D�N�� /��T�Δ�{��H�{=D%����鐛��;���hCH���3���^r���1���t�^�Nݖs�8�X�̑�Wɑ#d�����{������g.^Q�y�O�!y��\de.m2� ��c��7����7�{-����s��(��*�y����,8j���DI�|��\Wyl�TYen��ī1��E^�v�χW�.#��>���-&�<�`��C��h�Ėu&^+�\�&dç"��YP����"o��<�fĎ<h#�̺hӑ��&�r�h�f~FK%_b��	�aN8�r�����b#(�._���vzrl4F��e�R*C�^�R
�%�8)�}�ּ�������}�b�>�)0�B�5�99J8�0G7@��K�N��Jg�N�a�?�� �Ԏ�+84��Ҿ^���丁Y�EM�v�b�gGTT���zm��c��I�N#|����2�`l@Gh��MB,�A���l�֏<x?��K�)�G�"[h��ƪV�f��g�d�X�Ws<���}/��-oj���G���a����g��~�e�f-���*D.��� �@�}��8�6�2_i7)Cm6^=Te��n�:��3�e3-ǎk�-��5^��%a�5�Cz��ృ[6i �;�5�Nc@R�J����߇�&���2�硶�`g�;���I��g�c���*��5�^k�O��i/|4�I@����?Wbq9ď^V��j��q少X_���RXR7�sk�	L�.�AD�'թ0�9FA�8���Q�çW���t���Hǐp�񋸣C9]�d�T���������A��|�Ǥ�ؙV�>Q��z����W]袻8/1{�J3��t�C�Qǒ-��Ȃj�l��1&*�uzl]k�\��\y}�wQܮ��J�枙rK�Y��!ya�D�dj��YB��w;�8���H'�]��|9�.2�������-�4��[�s���H������j��A!MhD�O��`xm��;$6������I�?�0m�y�d�����f[��8����KB?=��jr�����D��a o�8�G�7��q^z�N�S	�u�m#��#t�`}�>��O�~x
y��W� KA�N���`��~z_�H�pȸQЉ>lS�z"�{�f�F�R�(2��K#-�I��)��|T��$�*��������%}*��g��,���$�Yuɛգt��Fp�(�=��� "�K;-|�+TdBm8��(�)ۢ42���h��S�t�
�x�c`��PGh�&ϸ�p�E�N�*fJ���9�H|�X,:P��z�nh�,��g�
��m�ɩ?;��dc�Vgd�qy9~�{����ㅛ��o�����cx��k��Q!�Fit�P�>����V�+�p�VH�<ӄ�])aEG�qSخ� �MÌ�#M$/Zib��m�?�Л����pR���|pwҕ6l9AF
NF�I��~���˵�m�c�i;���-7���<��_�y��hEzשz��+�K�ɪ��44�C;�s�A��J���NrP��B�$0��hr�V��(�RW��. �*{����vk��?�04v
��5��������e�&��fK��U�8�V�����Uzv;*8�	4��-8������ ��7�#����wY�D�J\u4��=��6쵖_F�����̪(&�]�o�Gzg��M���Q1S�k&��$NEW��� Lם�uG��Ev���̾3,�GL�V�ʇ$�T���?Q棈�s\Vʛ|���E�t�:b-_(�/��{�J�]�p㴟��c��֖Of�S�����.����Iee�Ǭ��T�p�#��&}���`/r��rU�FϿJ5�d�:K^���q��"��+����7�Z�Z?���{F0����ߨ�����ۑ���+���4�V�;���5���MV���m�접ҟ�d`�T�C5�O�}U%�������ptz
W0b*#�+��4%;x���r��4�����b,v��h#����Zǅu��6�`�p�
���{૯>el4���{q��� b��:�$G@�
��re:�{���߳��)�%Z��d|CKU×��<��KP\�V�ȯ׀�-e�ȍ-ȣ��s���D��GǇ��I�wj��s��˘�L�v!�qܧ6m��?_cl?�_�|��Ls<\e4P��[DP)?�F��(8q�$�z��pqp�k��d�3\s�hW�Z`+�nh(�e��=bi��B�2���W���!4�G�(E7)N�bؐ�..��.L{�i�	k�����c�j	eVNm �t�X���UJ{��[�� jG��8:G�'�(�n���E �D'%(�A�����,��c߻�J;����tT�Uh�O��5@�p�g��>��x��%�/Z�9}����(���i�puKp���M�� L�u.��5oP`��.���FQ�'
�iK��������Pǻ�qLg���J����7�	Ͼv�;���rr�u���6�H:��UX�u�N��R��Po�ʭ��dv���0�
m�ˁ4N5x�����f�Lw�%4�t���A�>X~U`����5��)'�R=��/�^g��rϺ���{�[����J��b3U^2&o�ws#@II
��cҏe����<��bS���JG�.�+�Ge����S<TQpwy�x�^I�GT�4uB���I~��."Dx��G�B%}���Ѝ#��ŋ��6�v�f_�XB'o�N���u����&E�IQt�Á���r;�r	-��sȟu��rRǶ�R�!��E��Sd)��`�"�@�44�a�OGL�M�7��iQ�<o��!��ț:Z?=~�����O����u5P� ߗ�[���8+y�B��>kX��Q��Q��='�Ee�E�G�7������ ���ލ���r�yq�%.Q��Bz�A�4����z��b���wg<`�<�Cx��9��D{��գpxz��!���mG�'ɞ��G�
����5^���l0z��f��6�d!{e* �,[�~z o��>8y����1�):���lOB�~�ұ����6���t?<��7�}�:��<��Q�ף�C���	����\n&�̮Ï��CK��8oj���7��X������
��:4h�Y���c����%|�ީ?7��H�I� 狷uw�e�t�e��fִS��Q;��`˯Y$�-O�{a�F{?��a�N�S�<V�BZ��!b�����eo ����D�c5ΠG(�t�2��h'陸)�~��,^UO�ja����&���� Q�W�OA���v�<�cX�����l���WAV�ڰ�&��O;�e
��Oau{�2
$�~<�k9|�)���IO�Y;&O۱�7/����k���)@�JBșju�T�N�ی:�8-q?�c'��PW�P�aqk�������^���l�̆���0��ɧ������+�w�?��=1�W��tN9��~kq��д������^O�N��\|����Q0��ݜh]v�C��z`ڬ�M�sVL��O�ϕ2
ӊ�R�{x3>��Y��:_�ꚫ!���\`irú��E:q�Sn���3�����c�A(o�*S��D��������X1�~����P�*�Ui��6͇��N��21 q�2H�1�)��9H����vp�ڌ���y�Q<r�]R�J�$��C
�c/yR�9�!o��N�K(s
LN�Q>p��؝1��n�l����e��Iu��%��1"����K��;�ę�~/O<��(���]�#�BV7@a���&ΐ�t�����}���s�Q�)�ê5�7��_jF��!x���/;����d�Pҙk�;l��JX˨�Z�oY(9$m$v9cb�76�d��7�4�������O����4m|V��g��3�)��9�y�p���y�x��wc1h��9�@�x�	]�����ɍ�%f�-�t���=c}h!o�h��M�h�~ý���e�'.�F����^�?��,�W�I�|2�7���o��._B�ˌCJǷ��y�Mjx������x
��i��I��RV.EQ��J��՟�X3%�rM�V\ս�<2�!MN*��iP�'Ɉ�'�R��y��2z��ix�P�ÎD7���uWE�)i�V!]<��N��끒@&���~<,����L2�Ch���o�x���,�9`:݋���0;�� I1�/�v�cS�����A�e�ju������|�s��$��K������sR�ɁQ-�Ż�d�~�C�"[�V�)1T��=#Fӷ���ן~^��:ܵwq�b����ri#�a�q��NS��^�:�x3qs�Dbp*��%2���|�޾qp�M��L��\o�ޓ��8�h$�����!��W��?8��'��c�����i�����5�����I��UMdB����xh\,���{���"9�)�i4��H�wm�Kٸ�y���=���5,�Ҋ�^s���O���A�T3���B���`;�aѽ������l�G�%�/M~�����ۢ}�x@�y� '1��B����QJ̬�;4����M�(��F�6H���ncL�Q4g�
cu���<�PI��15*�B��ƼC�hhK��+Qr|J#��tn�a(�(�Y����Q�3R.	�)}��ۋS7��m~���)z���%ѥ)�$ᕸIN"�k&Od=if�g*wV�Rh`3*21���Ff��j^����=�	 ���fU0ֶ��iK�N
�H\���8S�X6}_������\�q�;����x��*�~mn�Mh��^U� �'�+��~&~/ҕ�%JF	�rܰ6}�6���Ϣ(�@��W舑C=���Fs_�����jGt� g���	�Ȕ�0�3�!z��mN���A�+F>��p��`�k�Y��~]��O�U{�V�Q!
�Â텰�Í������o� �g�����#����+O=�z��K���E�%+�q�l��Ɓ�ѝ�%YZѕGJ�3�q ���Jޅ�j�k��ȣg�Ў�L8,}v�U��7�>�\��B�>��1�c:�4��E�Nz`9V�CY��7��<��!�yܓV�T�3/�KF�P�x;�(E�?@VGy�e�n�������Q;QO1���*�;SP6U�����XC=�\���� ��� /�X[桵V��z��.+�|�m@;$��G�%ƣ�0�M�e�uzo��S[�3s�J��Oҡ�*��}R�_�x��W�G�`�D��4�|�,CIa�t3$�����L
;���|��H�9ܖG�n6Fi19�)|��_���c�L�X��Jw���@�Cft@6���ږu2����l���6�lfz4�8��Lk��/|��~�ԉ=F��t�j?ӯ�H���g}z�<Bd��i4]NGn�b��i4��k&�ڒƪ'�(8�FdQ�h����^:�6�)k�0���Љ.s���v����B5gOz
�|Y3���6����^[�u��>�>��GU�>tI9��3��ʑ�e^9����(G�)\_�~����.�@�,?�ertL����@Q'P�S,}����ˤ�d�w(S9v���D���>���1�Y����u�I=��Q�'9��:��灕��y�reT���	L|%�T��4�D�G�B�1ް�J)�HR�0�"�q�Hhن�|5(ֵ(��٭��j����݆@`YH��ͭ^����w�ڵoz������<�2k�|�K�19�9���v:�~��� x[W�S6+� ���k$��'Y�{}�\e'�D�̪|m_Q]*�Y�M[>����YY��&�1hx%O��P ��9bp��>��_�?����'���(����8�ӱ����'�C5\l�a{�z�K�%�i��H�� #}驪?�	�T��� ����d�Hv��"�h�`��~�0����:�eNm�b?������o=�E�\�w�Ҫi��6L�;Ķ�w&I��N���~V���e��J��EG6/��g�5��ؒA���m�c�ɳ�IJW�������^箎��p16^έ%z�;N(+��s,��?h����獮M]M�EX�bw�$���g,�C�j����p�&_vҩ.J��2߮����z|��3����.Eu���f���I!�NB��YZ���A�:e�����i�`	�f�/�Qj�P��2�3���A��2��,��6Y��z'��qՖ?�!`�?�{�`&/�I�l�~~����?�C����߀��.�c2\�4��a�0&�<[E�3���Bg��8UТ���	9����;��&�$~�<�'�������G�&�n���bX
4�y������^�q^x����}ħƲi�a��{�����{䑖�h�x"x�Պqr���?�9��[���Iϕ�wz��	�ŏ���|��:�N/��1}���@�vN�d��_�<�5�
��S���ʙS�֥��)A�aG�,�S�g0�4_zQ����f���2^+z������
ɯ�)���#5�D��}cM���kue�u�5X����q��2�q`�$�yBB��wP���E %�C1jM��'j�5�X�&l�O �}��vRO�`W�~��$��}>���G���Wz�����Y����P��9�	��F�*XC��l��y���|M�l��|�z��|�K
yt�>�S%�F!�a擳�)"؜΢���i�((k�I�f.�u����	���G��ۨc���MQXRMެJ�I�;�h������h=��x�+�<�q7ebg�����U;n)=K>w��Ϻ`s��<'A:Aw*��
xajG���[�/"�{�V$']�r��7m��P=P���ۗ?��`վ\����5�ɤ7ă;���k�8�z�/��[�3�1�����0vJ5P�h�E��jac��{���W����C�f�>�A"*��R�	}��E�"���u�Ĵ*:��'�91V�<��+&�����w����kN:�C8���a���?_��w���%��_�T���1}��w��=���&11$gkPW�;�[{��bHv';�8W�z��0�i_�9����� ���_@s��vmk�	!�m��" �`:q��*<�ʁ��>�9���矃ã�pǥ�-���D0�C����>�����?�W�L�SGqD�RJ�����B��c�o�j�#�W��S[n�~����*R�|�R�T�eu�Ӽ�����'�b/�걆���i��a֙J�
yr:48R��t��>~/�:Z{}����uz�*���C�����"e��Ҹ�zV&Y��4w�h���4��_2L,�����31�H��H8vG�2.+^J�0IfZ��I{�pr2�+���N�s�����0-�Ai2��##'���ơG��+�*pEa�X�f�F));_w�]_����6�n��%�}�w?c�����lԥҭ����aXͪ8vN�~�����o��߁K!��qH��}դ�ʪ}R�����:�
�J�x��]\��!��K���Rt�x�A�4���/�9����7����m��P��ڙ������2[�Bk����K^pմ��o£�~
�v��-)B<�tZ/�{T#~�	\?:���O�ӇG��QM����"�ͣy��*�-{��J��.��zӗ:oh�0�����s�R[�-��~���4����pB8�[��}���N�W��Bh���ǎV�_ԱZRЮ����o�z҅ �V����Qʵ9{�՞�;H�K�c�e,��<�e'}/���2YW�XEÎ��,���C �p��z\�|��V4~��Sx�� >�#����Ax��e�N �������g��\tΐ~ �\���Ӻ�&frʆ�;��e�M�+t�%����;���x���%��姪Ne+�e���Jʡ��A�y`6����z��3�N
�Gi�������l���_�o>�<��u8�� �����҄H�Z�QyXu�eߕ� ���P�kǧW^�/%eB��p1S+eb��2�q�lX�~7I��'��+�6ԗ��h�<��+/��Tb�ܹБm��y��1FG�wr̭��˵�ͯ�"n��l��|�y��e����8V1#0p��F����<�:�� �YA���ZƖ��mc����a��AI�#��K�Q;��Q�	�biӰ>�YK��X$���KG��5�Gw�x�B��]�&�����[�>��w\�kك�9E�:4Ur,��h���^X){�?�f�#�ゔ䋂-ơ�%^�Ã�N�O .�p����w��}N�}C��N�T�h��l�wl0�M&��&�ў3��cϽ �]{�<����d�	���Z���s�\���S���I����	L���AQj� [�Yޗ�N	��:�>�҉�Ñ�G��T���(�<���S��27y�:�w`�����!�q�^Zh���ȑ2�/��U��er��	2u^���.]bX���a��}�K�|�+?K���^U�o滈/�C���fa ��M�A<L<��Hʟ��=؟��v�Z\�N[jT����ܟŌ��X	��˵rs�R냎�em�����^4{�;|���TR���� J$��w�"2����"����cF�J������O��y��Ï�"���B
\ǣB�S���N�,r^���2�.��׏ :�9�2&Nv�~��&5��վ|�|���2/���.�qQ��0	�zKEz��&[`n)���a�2?�k��{�k��?��pG�L�q�\Н{.m@_��7��{n�M� ���>G��R}j���
N]�[��쁞PѝR�"��4���>��ɫE���¸)����44���#�2pm
���gg�����^�mݗn��wc`[��)��2' K�s�Kr�,��`ۃY���x���Ά���=�j5�g:�����sw���ˬ~�s����Z���Ā2�̧S-a���O��A�G�����w��^�̾�����bT3��\��6�r�-��1/=�s`y��K#'i\���X��f�N��������A����_�N��&��8<=�'^x���?�����y�����tU��%	=���vj�1�7L�I��*��@��밑���<eC�M�^u��2��s���d��)^���Y�J�2R��]$���u8Ii�Pi<3+�O���`aHQ�N�L%�I�˩}"ߘ���%`�"��Jz|~�lڎ4����O�ەe�Lkol06���M��(��'G�
��k>�|�9���������_����� 2LE��R��'�)���`t��m1��%���\<����u����Vy���᏾���/��|�0ٛ�(��Z�A9K��y�pJ�0��"Gt����m[�9>�?�����[���/I.	�'p
��'��o\���|2�8�RM�p[=�k��|a\#���=��I]�%��t��QBG�zdK6�u���H��bt��>k=�a���D�_u�#"�@�;N%�Ʒ+�S��L��1����>L�S���s,9m,�f�8�4��Iʊ",���*]G�Bc��.wM�\�+�3x��U�Zh���3O����!�y�U8t��J4$Wi���Ta.<�t�)F,@��`�J�u�dӦ��p^�MZ-���31��{s�b(�NWD��O��ѩ����d�
<���p|�>��7��=�|��o�����p��+0�L=�z�x*��J�4 �3�AҦ��c�<�B��'�G�+]�]�{t|�ׯ�w��ϼ�
<��w��r�%pu������{�g���!\��lxR9rr�`6��KO=��o�;�/��{�����0���c��S߅��?�k�I�6%z|&�F���	����������J�0=b�� u)�E1�s�	�
�ςB	��g�'� Ph)���6�k���9�r<[��4�S�=��S�]	��)�v���m��۸/�0o?�û�]YG���TIڒ<�[tb;�s{CQ&=#Ч>V,	�r��R� �DZ'�%|���!�H�<Dr�R��1��
��\�q��c������w�Ar���N���\�Lk2�U�9�L��0�����B�5�\�SO?��*ԺvP��	�Lρ�CE�>��)���Vj+u
�B��N��K�)��C����߇�����O>�e��,)���I�t��M�G6ȴ0��輼b���t><RٕYט&,�Cg�D]�+����&	��s<pE6k����<���\���aXE�������y¦��m?ృ퀹1Ɨ%]m'��.�����MM�:�1��EN�:ʵ�3d�XrTP��}�ɡ��d�!�O��W��Z��&n+�R<0� }�p�5\��꫗�������~�	��w����py�����/�q5�<��U(��ݧiR�ȗ5�D��h�	�Zy����vx�w�5x��W��O>��@<���ȡ�"G�ߌ&�N֩r0?ٖ�������g?��f�+�0ܵ�Y���N���	��W���/�'�Y�t�V��OqQ�F�4����~)��#��9#|�mz�0���)é<�zn�μ��&ْ"�fx�k��м��븰����{љ-�H��� �JA�]����f�x4�Y�R$����8�\j�xIۻ�*����R�81�tBd\�C,X���d�
�&5�vg�?/��p�G~��;�0��1t���q��z񰣅�d$<��m.�%��-�&�g��V�T�8t�-���o����$��/L����]B��Q��7(�0�������y�U��/�/|�)�^<-�ѧ�4�!��;gbprNN���P��l��ͪ���F�5X!#z�\�I�N��X�t�R\4(�P������Z {c�&*/aoeu'�(!{�7�%u��~���=�E������S?����Ճ}x��k��Ǿ��ӏ���Cp��p�e�x�[�C��,�W�I� kN��,��2tF��a�=�&���p(䓞	�?U�+��S��,s��6���v���T�w����l���㾀��E�g�rr�YU)�p�����14�nUE\���������,���uB�A��7��I�y4�Q�!�C��o/u/��lc�m��XKIP�[�$j5c
T<Z9\�=��0;"d�NT��-�|3�����~������w�;Z�b���}�^�� '9L�
��;p�2��(�]*�ެD!KB�����pZ)�X�L��W�$�%�<I�H9@NC���������~|#�;�����;�;�?c6G�&�BNW�hz������Ҷ�A���rJ&TmYZ��4�z�P����2���R6��>28��������B��t��nn]�BZ"պt�sIڕ֑�m\�X'뤳��e��m��\/�k}5���!��9�� l�ڴ�Ѝ��.�|,kw�Xr��|#p(�XQ��xR�������?k�X��	K�z���-+���{f�ï`_	?f�L ^k��=�]���ς;���I{�i�fy�rTd��y�a��^�<�/���;e䧈}?4�k�[�[|N�x�b����w�~L�Q�U$@9�,�N�v��4������]:����d�y�����}��_|�և>x������+��/}~竏�k�(��?��b�3I�sT,#�#���W�n��`r+�(�)d4�Y.�G���@\h���Y�G�C����Q3��\�ݯֱR־"|ֽ���8=��@���Tr��b�&���m(��	/iO�_�D/�>�{ih�"G��P	+�\QZP��2�aC�')<�i���	���T6:e�:,S���|��o�/�[����'A�ZOڅ�4^=�U
�ĳ���铕$�0 ޯ�wᮓY�r�	�L�9N}�ޛ�֓&%\')�@U�y؇Mw �CO$��3%�\��t�I�F� M�i{��a�qGF��o���n|��qL��|t��!ù���L)�3>o�]D��(j���=s�.�Fs��h^���a��J��L���ĔЦ��5����*�a��[�|�k��;���Oo�������?���\������y��~�� T9�:!S����<���_^1P�8���{��xc��da��̫MA6�����N��d<Le�-=kR��{��A���c�x����%9)�3�{̀�u�*�n�x˙��v�9_(��c��s����(�0�TR-�ws}m&g\�4@��1ۇ�*��eh��wJ�%hAD?�:6���ϼ߶��z��{5�bBG� ��,�,��$C������a ŵ��^�ᵥ�C��h����Я��-������$^^����h�6g� ���ݨ�<9��]�
��?��p����ϖ*j�Rģ+^���)�&Q�#td2���r�HƵ�|4��g,2�|����;���)�*S�aYN�L����W�)|������S��.�{�i�0�jP�:t�F��P_xʊ/Ea�N+��.`��Y�q���ټ(�������i۾w������y��~�Shl䫜���\^��(+D��t�|���=#�ɗ���R���>e8���S��zW�k���u�c��T�h}*�uL�u�C^��<��:�����1�|�8Pj���y�9�e�w�ƾ�r� ���x&�Ϣԧ�$�y9���|VlB��7�\�����_G�Mݭ>����
�Y�������<�}&e����a8]��M��M�o��t����ūC̻�YÑ����P��l�0��bHE�
Ej ��'�0li�6��e�0��'ߕ��T�j�Z�@��U(V��OB(ؚ�������S��W�S�>���wL��Ҵ��_n�	��5�%�圓qB�\����L�=�o��*����`�J��
)�s��$��XV<#8R��ӂ�`2���Jz������oFٵ�M�az��L;��L���+�M3�03%�Mx�N��;NR+�>�L��Ƥ�v������U�,�$�PUјH��u��P��ev��(?s`Q5�u�F��Lj��\����9����r�������/���砹���I� ��jh���A#�Ó,M"831B4�׮���3�jYcۢD)(ER��2A� r��,�*�(�6|�ycە��騐T�|��f3�(d���+_E�ͤ����*��Y�4^a z��W&^m�+�(߄�PE��)���n�W�T�L����S���Nт>��@�X`D9����Q��*)~�':���7۹��q�hO�]�u\�CUdd�y��C%'4�M�l�8͗�!���4��8�����S�ڱ�ƞ�q�hkX�e�20vm�V8e�ߖ���4#ش2{����U�C���e�cl�c�.
ˌ���<ϱ�qȿo��)-�J�{ǿ���z��<�D*[h���u��K�e���Gaԛ�w�v,��߅EL�`�Wߕ��H�h�x����{���w����[��+��� ��i]
�~�����%F�S9�aC���
W����|A��U^�'��>��$G@�9"M(�R�z�T��9R��w��>��4�ZR�[| �[���*�_����1��5
��-�!a-����R�έ꜒I������38冄"��x`�^���W���n�Z���� �c��i�~��?/燱�B��O�&'�ܡu�|����)�`YX��E ���:����G���y��u�s��j����UR?��:�O)��+�y�EuQ����cl�^J1��ĻF���,!��]������bWٴP	��������8'��ԝ,�Q��{�����$Y0T�X��i�Y"0�?�.�ǘc{��|u�n�;fB�Z^����i�|��Sr(�z�V�C'_�F���Q�˱6nb�I��y;u2�t��E�L�ˁ�zfz��K�kkYJgr����x|�U������A�^���_�-9�мt .�j~�����y#�D�g��՟e(�LPߓ�A�G��KE��A,�[h�z�38M�u�p4�P����?��Ž�6����\{�Ix�t���G��ʝJ���eN�M�\�'����5M-�LΠ/�i����0��:i�y8����^�?�b�p�2��1�~'�'�Yte!�ۢ�/m��-���1>M�J%Eψ�Z�N��M�±Gw��6�a��Jw�� ^j�(N�R��"��ǣT�	wQ�Z�o'�.�R^��vb�¡2�^L��\=R͆�9�p���FE�6�js�4g�+c�Q���2��uy&�\ǅ��R.m�;U��Mb�Mu�ӘI������7�l�����\4���XX����l���}@�Yf\����"�ǒrH��$l�8:?��}�a]�qv�C�\��Q#�7A��s�+6 e>Ld)��r`x^�_H�>)� ϊ����@�ǧ �i��̰0�iR�t�M5O��We��[G�K���K�Z��#9��@u�;}���w�Z�#H�"���L.�a�S!-C$�ۛ�1�C�9�r�Yxr��w��Z~�OӘ}�k ����ZFaﭢ��D{-o�[;o���y�5��`o�u�l�}�qw��B������+@��ǔ��)�����Ά��B}�[��#�a���3�E���{K�y:�'2F��W��Fw�H�7}ו�8�w-�d�`�
P��gTe��"q�t�I��Id���ٛN�a�4�����Ti;�O�`ڬ$��7r�*��t��J�2r��:ȓ�p(�9�"qD ^���7M��`���<�)��'Y��H�h0�2ٞ��>�QWx�4�<�:�ǴtM6����A���.>�<"{���"�Y��v��k�����++�tfYL:}Mpޘ����� �jꛮO�2{���8�If^��[ʁ�50�m|qfȔs>�;@9[qM��bJa�qb��?U�W1T����I�O=	���	��c�/]�n���I���j�5�>���1���ܡ�c`�7�:�8�\�
jcֹc�5rV!���H�Ͱ� 34����m��B��l�y���왥���D9W��Y��
d�r��H�vjMz`�E����:�R��c�P1�`ʤw��K^�Z!��v����)?se�+;z���.,�X bH�"tK4#&ۑ1��h�����VEXV4���&?|��1W��q�~y.ʴ#�����Q�K���F�8�D�^a�Y���u���S;]iէ�+A�cf�,7Ʀ�ԉ�e�Cm'����t,N%��c�|� ��8O���*���*�-[��4���`2��������'�,���bk�|绌+tf��"F�l�[�f��3+� q��Z��c/�1L`�!�Y�hP�j8��
s=�Ð�H,����3� �ȞNM#ᨳ�/M*n��-��,� �Y�G�B��4�FsQ./���ؾ�_��˘쥊k'���8���L]�/<�������zDȄ��O5s�9�3Uݜe\���~���0/=�L���+�M���б��۬���)�H?��u:$�7��Bcd��wcu�ֵ,��%���c�>oXt��m�3��#������`M�u����nn�:��}㰕� ���3nR��{��s$l(�(5�g���J'�)��N����N5��E���O*7D� �<{�f�%�ic=��b@�����<Pm#�kr$�T̬�J�V��Nϑ�e/���	�l0(�m�b��3�k�v�3�P����Q�~��:��B}��c�=�W�rԪb���/h���-���F^ٮtW��x\�#l���b�m4�y������v-I���!�dW��7&N_�'_�\�ٺ��[q�-P�b��G	H,��yc�s<�ɞ�Uݏ�Z U����p��S�U��7�G�4�_M��s�������~����>x�q��ov� �g1\P�~6+ĜZ(��6S�0pU�猪�_e"&�'��v�S�)kjp�t�wRN�<"�B�9��������<3?�c�� ɝ�(W���N�rb)��G������q��FZ�2#��Vs\w2\V�����c�s�q��ѴD�GZ`� f�j�6�x���LE����J�*�������ƧI�����7en��g���I��Dڼ0-�V&�.��¤e#���r��W��X�dʺ༕|	��������V
�k��]C�̙֜���a�[v΍Qob^-ƐK��z��7=t=}�XD��kG���2s\�	O����u��`6	�
;J�u����0MeN{E��2*]~j&�+n��ᑬ�F��xٔQ%��c��T/����V�>�M�V����PD��ȋ�<�d5^g��ꩇg_|	��5x�{�a\%!�I�H7�(獄!�����+R�a�/I�f�8��^�%@�J����e���|�ߩWμ�xf��������zO������uK'�0h�]�[}�=*�[���m�@�t�݃�3tH�1�Q�̣(��Q�m���yN���e��R�ͬa�II2H;&*��}K����>I�:w߯�GY��w]�v�Ƀ�@5't�����z�x͋�'�k�<�C��c%��)�)�ֵ�K2A��̓�����Pj�&��k�����<t����L	�*�-�WX�v$-�5�I�Dz�a��w���f�zm0̌�y;��{ֵ@�O}�Z, ��d��p��(��d)��X<�%�;=��j;��Ď�3��\
Q�ڱA�z�Zud���+Z�a�4����<#�J��b$7�}r�<�����o._P4x��<�1n�R]i,-˯� �}�d!��Fr�	ӣX��4��D��������.�s-�5�Zr^>��z�����٫�3P�<��*V���)ՎWOË&���.�tZ�ݏTw�s����(�Y����~?KE���*U�Ber���<�I3�����.-\i��p&E���N�q��.��_�����?�������
�֦9������ z�A\6F_��>���p6l���~����|1Zɑ�m\]B�^Hu��K���A���$�+��7��!���E�x��bM�.��s�;�(�J*zf������PAsD/�2��T88��
��!A�tjW�X�#� {��%%���1�F�~U�V��
'�����ľt>OG�$�������s�~�c�C��#���L@�ui���^(m���:\��!e�������tY#lu��B�%ҭ����U��b,�q�Y�ݼrw�]з'��9[θ�9Ot*q�p���0,]�i̬j�\U���yr�+>5��A���nZ]�-�%1��5Yd|;y�{�_���)x��{;�sT���(5µ�)�G�C�#^���^g��U�����9uZa�:�-�syAsz}����A������\#���I��"�/�z}��09�o�Z�M�}�$O�k2�UY��Lh��r�O�M318�̣�;����b:�ҔR�$�2n�	yt�!� �.>"7�n�/�B!Cr�R�,�Z�R9���Xr\>k�s(X�E�H��s���u�����~8��J{u�L��5x����5����4��Xc�l��1��/:l�>��*�˶Q��9gv
�A΅�2uy��2[���"=&��
������\͗2�N4�wi:���
湝�_l�!g�����8�0o��G���󺢙��m0Na��H�5Wd/��o�K��=Ba�3J�(�K3y����1��YE�/�����%��{	=�u�3g�?���ٛ��_${I��z���H��9����.�q���a�"�����=,���j94�����������3\���.�U�|���1xu"f��ޭx�J!k̛p��%h�)D7�kB����O�>>��{5>�mx����s?p�=���C]�򚦂*0*
�)��ڨlWi8�2Q��t�[�օWg�vN�"oo��D���B�J-K��2٧�����P��7Z����i�E��⩂pe�#��]����gU�*<{\@�͘�8p.�f(렷}�g���0C�YG�LQ����-�
u]ag��]��mX ��.T��܇���Q@���wf���e�P��{�����K�9}���\k�Mij�Q�o�Zw������a���|aۄo���|����-|���S�kf`W���;��m���m;]I��uX������<!p �i~!QJW�o��H_Yy��9��AG�>�忀_����^���LN�B@��*:�$�x�R�J�eo_�t��A�A��$g�Y1�e(f8}k��Ԥ�	|6��mrT>~G�^�C���*{G��)N	�8'�x�M IS��b��<݃^}�������w�����R��$�Q#�>,
,� ��V���e�j1�)/!-�$,�y�"1�6
.�'��e;3���zRz����<x�xB�"cɶk�$�P�+Yw)���y��}����`���~}��9���K@�{Q�&���᯵�����:�4�
*r~������eߵ-�����ҵ�d�IM����s�Z-z���*]%�#|��V6>�톢V�*\e[�UydB��偳d�7� e��J���(�YG�T6�`�DXOUh�r��H�vm8�aյ�84g�l0�^�oz�94�����1(��?��s�&k�C;ςԪ6bm��~�=����R����de�d�ᫀ�{�? ��G�,=B�r�,W�PKF��zJ'�5Ȥ�Y�Jes��މZ=E'�ěP���6I�::�Om�]WQ���i��_����g��g?�x���T�< ����m�ʕ�AŐW�$c� 6�Z���pld�����1z��o���3�󙟃a:[�N������}��K�R82�8��.�_%��8E�&�)h)!O��ݛ�#>ţ��f����R̋&��?�F+�&p���#lzwa��=՚X�(�%UrT����:!��tPO�QN�	��eI�0y��}�Y��(�J��p�ꍈ�9�T����bi��W��n�S����uj;A֨ �1�H3f��L�PbpqP��mB���D�v�)X��=�+Ʈed�!��eSY��0�0�`%8�=e��Dg9#�/D�L��<~WY�}24�S9UҠ|#u%�R U(�x8�N�?~�k��K/�;�z �%��i#�l7,��2���0kj8�5@�׭0K85�$n�j���� �K7k�7��q����d�1)�h-�W�K����.JQ�[����I�޹	��$�̆���QΡ*����٬�����c/� ��S��G��\o�<	I����
��!#ƽ�3s���U�;g�5�J��{չ>� ���>���c�!!�0��N����zf�J��,r0a��#s�YO۶A��O�σ���`g�+�[bvn�Zt��{Ŵn�v�c��l-lm����πD���g�P�i����;�kY��=�ɡ����,�-�-M�����BaB�\^6��A�T�8ã�F�����^{��b���o΅��������7�('�n>��wO�fb�MF��Q�K�&=�`�ӱ���&Y��m��P��ۣ�G ��N�*�l���E!w���(�ت��� ^��k�4U���d
�._����g�?t�>��*_(��tV\l���ë��"F~���f�P�",�k�t��	��*�v�x��ǐ��Ѧ9������$���>
W��%�L(�{6�Kĸ�G�ܨ���*w^�E�ť�y0�:�/�)��_Z/����ZTF����\��\�]�e<��Sk1����NR��E?���V7=�飳�!��'���L)�6e�� �!�D�49a"X�8=���r�n,�{�x�jGϤPP�3s�*G����`�PZ���Q�E��p���@�!#C�h�lv;dKZ��ݶ͛�s�-�EI�k��h
)|E�1��d�y�v�Q�8nJ�豴8o����m:�6���p�'��S���	�b�a�ҠJ��sK�~���M��c������r����sIb7 ��T�uOğ*װ�RD���.E�K�M�����������Ga�1��������rc5�����O~~��'���w\��+p$f�����H^��$cy�b\�:�q��}t�x��[@�s�Y��0�!i?�ЀNۅǱt'��}W�w��MC4fA��`���i�K�F�Dxw:�ptr
���{��/�3/��޸~� ���(�gi�ԨpM�HKQ��Y��ã�J�vة�Y�J���'�,�����j��jY���5b�r��T��4v+t�"�p-�P0^?MAι`bNq�]a]��E�l�p>�v���6�s:�	�[�֍���cn%�[��w��W�E�97�/5�o6_���y�� ażP��P�g�X\�� ��$SAv���덌i_�B�λLx��T?�@q�j�b�W	��v:1xjHF�9@'��rΜ{�e� $
�؀Tt>e�BL�<��RN��bnm0��&"`��sA��
7e��S������t{A���������z��h�';K�C�.D�����|�J�	��uJ���5H���9p��n-�C���%�?�L)�)d�:	�D�Y�S�����+��ͪdt�j��1��O+�r���� ����}��w�K�ܩK�v�}o��4QeӀ�rȚ�P���8�csU�S�t�*9��� HAՖ>�6?�g,��Y,�ڗ�w�H�9O0����UU���68�D�@��g�R���O��i& m�*���'3+���OGF<ddp�w����C���a�_�4�׍oi/N�O�����<�̚��F0c�z�'��v�S�<V�W��g�,BsK3�����	����$;o{�ھ5F�^ �f�A���>ɘh��4l7�FF:C���	y��"c񼔱9���1y�3���ʻ
���/�Ȣΰ������������6�:c�!�hQИ���Q����(�m��g��6����=�uH}l� yr�O��)��祪�ɾ	b}��+�h�ƕ�k%�#�^�
����	~��?��.��b�ɡ�����5��ރ�n����-S5���|. u�|�J��kN'(��8Ƞ��:�18+7Iל\r�����D%Y��5,:2��w����{�x�5���;��]�p�_H�@��ς K�WF�&������fϵ�=�IKې��i[�,�#�@��Y��d�u�FXќ�����v��2��<tz�7;���7�e�z�'���[�X}-ɍ,�x���~�Y6�#$����k�%�c�I:�����dM$�3V�;sO|���0 �9o^�a��94OJr�8�8-;���e}8���V��x�NP�����Mv�@:�ܥ})�tU����״��x^z����,2`�@Fa�zQ�-�� ��9��Ns�s��d���?A��
t��!�w�5�����.
��v�;��>ᷥ(�y�:od�%{�����:hہ}o�Lקȁe��Tv
SO�F24�ݜ�R_�K�V�,��V^^�,��&�Łe<�$�~�y3Pҗ��aK��Ɏ@�P��,?E9�JNޥ�S���a��U�H����\�z��)���#r�M��V&��.���K�Ȫ�,y��b*d�u�6�.F�����3�4�is�2�8�x1t\oz��B�MG��KaY]]C�K�pi����?O���_�(��*�l�N t]!t��<Iuy��F�|r-:�6���*������!�e|��6= )�hQ� ��|/]N�t���.Vz�����^����3���U�8"lZ�Ś��Wu�)ޥ2��Q.�wz��{S�~f���*��åmgT��t~�4C�q�p}	Є��"�̷ύ*!]%C��M�\{�7�.N#9tǲ^�l�����*�Z'̛ԓ�0�4f+�J�� W@��Ki/*l�b��T��@>N/�X���9t�囧]�� ��?k�?�!#�g����m3l���9.�Yp���s�yN�ga���h���4YA����(,�CI��_�� �{}EFJ��CF�45�)�/����/�?��_Ń�l�A"(gM
g���f�����?�~�_���p49l˚F9;��(�7T�v�������JW>DبƻC1��ň���6'���੕�BFO�ȉ:-��{��eէQ.�ٛtuk�� �����K!dAK��Yw\~QwJ���ñ�!,�e�(K	�I�B﷌�
��||e!�i.�U~�eme�6��go�Q�V����/�v���y�d%�G��X�Ue��w��39߿ʞ^�ˆ�[���y�U��[c>C�q�W��ۭ�A\16�S]��P���)Ǭ%��`ޘ�X�/4ݑMə�^�ݢ�'�^���R֮!^U+���d�+s;P.�1�NL����[�<�Ke��"��2Q��b�w�8�rX�&D�N�0 N>��^�� �T�t����%(��$:T`pu�f�k�L�sy_���+RR��L ����p���<�CJ�v$[�d�:[ؖ��$Ǖ��nF��(���A�:���ҵ������e�?�ܾB獠w��ث�6��[?S��8~�@a�+T�Db��e�U؆�`�S����':�B�K�����T�j����W�çn�ɗ���S.����~������O�xӯ~N��r2�MJ����d��^�@ѯ/�;�mٺ-��.A��鉽r=�6E�K>z�?9\�YRN8UX9�0t6H�X��rr���y����wȗJoN��|��F��ݪ;�%s�:��t�@o9��רz�������3��%8]�P�o��#
&}1�/$R88�ҫČ8�X*�[o����:Vm3Hd=%�#%�vB��6�zi|.�xmø�'�)JiVm�"��<<�u�9�<���ҳym=�ua�{���P��rg���y E.��ηVw_x gk���!��5~�+q�w#.� ��NR�Y�׫l��I'�y^�b��J

:��2�C��&.*��
�է>��������5�S:5)�P�
UL�j����a��o=O��R&u+�{�TA�S��Q��CU��7�
��
 
R�F���Y��1��`���xj�4�h����H/Mc	�[ �%⻺�p��ah����N�E-���Z���⻏�	���/�D����A��q��5�����fU����=����n �O5�TJAz+�^�5l����Pr4 (�^����S���l4�g^�*2W_���L1
��$���/Oje�E�u+���N����n��[?tf����{$�W���3��S���E�� �Gr�Q�wq�H:0�F�j�桸�8�^��d�وd��)� >�ѱE����j�V�S��{˃�C�p���In"����u�ʠ%��ޫO��l���{�)���Z�2M%o1lb���>��|�e�O��D;�Y���:��@CnHm¹��?�����gֈ��ˮ���M�a^�v|-Σ-���;qh\�O�Wi�ȝ��	20)s�o�+9��L Uk�9�Q��2��I����aK�f��I��
f ��=/>�p�����wNf3T"��]���'֥R� ��F����P�`�@�m.[���޻ۚ\�a��o�s�}�h$�i��	KBa�B%ฒT�
�T�R)��ߩT�?('�TbʤRTH	�Wb!@�!B/�A�ƚ�F���kf4i���;�q����|�X�k���{{�}����={�����կ���cO4�m4y��Td���ák�wr!<?ߓʼ��.��i�IH�����ڝb"�A%^CZXw+8�w��:�_��)�q>�*ΑM���=�V���&S���5U Т5z����2uy����r�KO_�h,a	��``,��0�1�^�im��C�I��c�<2�y���B3�o��r�X;K���q�쐒b��%��m+��p]���l�i���ڸ�q�Ks��i(��ԩ�_Ş�q���	��~�m0���p�_�B�頋e�,͐s�@�_3V�!$���'B��FT։C������6Q8��K/������������=�0
s���A	�	�>���C���~3��� �ؐ�{���i�;&kt���C�����r�S�'�3�=�u�S���u�C� �ߩ((��Q�ZL���_�y��Ѷ�Y��ŕ����J�)��*�n��>�2
�I��)e-��� �t��K��J�0I�A`Tᵦ��g`�B!�ӂ��NG��JD�al�|�39�.~�|�zu�rL�J3���`J�|�3����u����<R\ݩ�;|��a�Өa�ä`���!�қa�~��/�΂���	��Yr�x� �(X�K�����ADj�s� �P$�(�8��ڪX2MX�C�Qu����2�X	|�2�� 
l���ϓ�*�>�mC;�τ���I7&W"�<�kRGmn����,�=����$!��&T�%�H�	T&�N`C/T�
2�S��u ��y[���B	���	bqU��Lۨv�Օ��i,���0�x ���׏����6���z$ w\c8�^���&TNn$�A�4�{�OVFUJ�@h�wǢ��C�����Bcn�t��2 (�*mN-��ܱk�_/��
.�)_|�1�/^��}����phOU�	,t��������.B9)WL�S��_Փ�A1�UWTT�²-��3|��&��z���=��LZ��P�J$�ѥٯ���W�aa�<,�O�7�0#u�*�{L���� u� t�J�3�G������fn���:pM�F���q������Y��`�C�8P�S���g)[XRb�t�(��=��z�'��	_��!}���a:��	��yc��AO=�������|�
	
c�,�q#��RB��~:�.t��i "�4F��%G�ӂ�cjW�\�Q�����f���*N���vՓp��=�Ή¡�Nْޤ�������r*�v���ۡ�����n3L?4^n��O����I�/���h�-6AV��A���L]cǔ��Ȋ`8o�%� i��GU|�q�
]K�f��Mq>�:T�Jǖ�hjˋ����{�������V~n"ߥQ��`x}wɲU����~�_���)�u=�צT�ꔪ��b�Y`[F��<�Q �0����H�
L����<7S�:A�G\��$�cf���(8��,�~��*�u!�JZO��U(o�H܃ eT]�S6�Q�2�\r���tx:�O��e�|?��_�;R��8������an��A;�����`ZBX�p�jƞ�ƞpwN'����Ը�DIz�&�:-w�$TdΊ�
�.�Y5L�������ǹyP�i�3��s�C@��\{r8�ڑ+�>�£��B�iUcO��}dgM��n/`���Z�yI��5α�=��L�����2W�i!�I��S脋Z\C����o�s9�����*|b�"݃s��w�=(����Ydz]�~G�2�AG^5G��ho�����m��(��:Y�H��L(����R�0���c����	������v�&�����4
�g�1h�q��ήj�l��U�B��_���p�����"�hs��=}�˯H�=��`̎��~��}� �Ӟg|���7	��#�5��
M�q�z�T�^��5#���(w3Fm����K�,�4Ͽ�����ËP��p�]��%h"�RY:ϧR��i�����S������@P� 
�ڇ)-f���lH}�����I/��2�Y0�=:n S�B�z$G�&f.�uJ;��DTs�-�[/�������o����3�=�z�f�G/����M!�rv��<�B�Uԉo���P��zUJ$W�N(H�	� �k�O����fI�N�d�Ut��a��,L�c����7�M�,��jTH��ΆK�C��GeF��B����/:��\����c=�Qr��[�0G�2e�~�
���L��d��X��0��� LCfy⣇����T)���0�H1��>$_2���/��f� ����Z{��NvIq��=PXw\R�;���y��3�$�o���Nva��@y��q~J@����V��_�����3��P�[�rFE.�g"���(�� Gu�g ��ۿo}շ����(s'w�ZA~�-�3x�]s�[��nx�_�zf�7��G�0�0�����v�.�sO���1��95�W�0���$<<���X�捑�I��NPa���|���
A*�m$�:*ԗ��F�hkNBm ݇��ѼZ.>z�M����7d�UӼ�VU���T�#�&+.��iƶ�#}�3Yuk�܇�Y�;qn��4����rB��ـ�xش�\��2>��Y�=l	���q��/6f<���4�[�#s�:��,M	%g3�@@E��&���p�T�S~�\�.������i��1�9��P��l1�s��	�Q�����D	�+p*�Z�Qb
"6t5.ړ�5~n'����tͲ������>��j`n�Q0 ����SW����>���.�ܞ����|��@�]k=��i�	4�2����i���d
���Ҝ��62�k��ƾ�=�^����0Ϛ���]���e���5�ƃ���/>j6�NE���wU����X��p�Ii.�kY��8���A;vaT|�N9��ī4��!� �$�3((O o�⯢�(�B*�QD�n�¼�������=�����jxaQìn�a�Մ95�<<.ƞ�+��&�üv6"p-�J:� Ġ���s�
�]��-8��&Q�w@��(��uxX��&
i(s�ن\~��L�QF#e�dӴ����Y��LG��]8$�s�Z��E�0��m81Qr�K8X,�w_�W��2���x��k�k7��ݸp M��zp(�SA<��H@Qϙ��h&�U�U��	J%���pk�K[����i",�C\3�_fchс���u�O�ώ7}vu昼�܏�09�Ӧ�>�î�<��z)`��D�K�ļDq�x��"$�{C�G4ɿ�\�{憪��Q��xJwN��b����A�Wg)B{�L+��s��#�[�q�/����:qQ6`�d�ۏ�����;���C��up%D4��7�s����^������%h{��x�k��`�<m�a�������0�E�;$[%��u�B`����EU�D!,���"���N$�����}("+|pу69��(� �bA�ЄU��3�B�3-��@�egɦ�=�vi�ܛw5������=�|~�F�����ʱpܾ4�U}�rN6�m�|JQ�X�*H���_PF����c��aAڙR	���v
�E~�`�`Ϻ�_�-u1�	D������I��7�����!k�'6Y0�P�3�^�Y��ǰ������_���p��0�9|�����V}`��t6�HmmDN|H#�:�G�U(�P7"���2wd�P�����W�*�4�g"��ċ�Q����`��\-��&��.��t4W���A�Q.���>oǖ�l�W���ˏ^����$��K�z�:8��v:�->�xm8�n��u�`��֍$����Pn,�
�lȾ�b��|�!y�..MZ��\)2�����e�tU��_��?�Q����N�z9i�W���>*.���D�쿩<�O�F�*�2�!;�f�rS� K���˳����)�0����`�*��]�h�f�r1i��^)��C������.~j���m�cv��+7��5�.��x���=����.�|V�K�
��z~���}�!�z������r���u*5��R�3��IX�{��jX2�P�h�$%�m�%n�TAI��`�t,6F(�q��B(???��爲Z���uC���(TM>m�gy/��t�w��î��7h��	��>9	�*
\R�3��X��UwYG[��F�t�g��4�M��ȅzuSS�������ȕ�����ㄝ�W�T>�����r���������[����j�8��(`,]$��\�rp�� ~������좕��V�PA�G�pW��v����[Ful\t�HI^��y���CHBW�>UP�|A����X��I���*�P�q�W�2�JN��Ě-�%��{��8�=� ���2���BѴ@�O"UPBZp�KJ��p~�.��ع��3�k��w�WL_���gz�a{h{ x%H^d9�Qo����@Ld[��*�T�D^RyD��EP��i]��
u�*c�Q���������cLلY�2Zd��5$�W*��A�#�����X�LA��P/���]�����!x���s+��p��S��������|�]:�c�4�le+�����������d�<��`#!Y�_������{���H4HK�� ����]"#l���j@�`��FB�h�J�L������Fֿt�9��������pbO�r�_��I*����Jȏ2Ÿvlm����*(��W$�PYUښ6m|3�)&�+�dB�e:p�	���'l6�Q���	
Z'����va�ܾ��ԓp�ч����m�J6ċ���3�`b��^�9��ѭ���a]W��R+3P����mt��t�!E x{���B��=��*�$�\��
ȸ�3<�#�k0�Ԫ@������`ۢ-$Q~�bٸq�t��#W�}�@��a�B7� ˣ��d��;�	?������-3���}���_w��w�3��'�~�C��y�Y�q�2����e��}T������CX�y��,˒Ĵ`F<�A�%��̗;�i���ǒ^{Xk�:��K�bo�f�Ƿ՞�ag����C�'�K�B�q�{<-O�7z�l�#�����#ʸ�l��՘+���q�y' ����m¨N�e�X��� �q�X�<~�����]����)8�8�|��Yyٿ3'��o�_x�}��?�C�O~�c�Ҭ
�G#Cq9,��:T��и9t\k(?��'�%M��
�X��Oޅ��a��zB�AF���<}>EdTT�R���!���4R7♦�_�Xc�Tn$���?��f�ѱ1�Q%��P;�(�<�	��U��g�KKg{�~-V��2:�U�;�Iw�E�Gz\um���]��Cq�ra��~u^שuA�?�ﺰS�N���>]���74+� #/A�h�+���rZ��4�c!	k�6�1@�%��O���d[@�Ae�Τ�M1����m0hk���y�����`�=hb��\^�o�t	���������;����:^z�J�+f�ʷ�	�����O>�I��}<^���H����������(=92��{�/fs�i��o�ޮ����J����i����Ջ�G}���Y�W,M QVs��شt�	6z�V�6����7������#�x�I��N`9��D8�j�
�=֡P\fs\��D퉺�Bci�5a�+T��ab�g�LjbxU�%C�����
�-�88v9�W�D�,EX�����!	�nm��ҩD�S9�
���gp�� �y.��r���7��z���	#]�E�K�s�КF��'W���C ����%#?fB2]�&�I`�↗(q2��-&�[��ӅX�����rۂ�,+螰b�Ȕ�̄�.�M����%1?/Jڏ�-:2�,n�����k��JHs�Zsp�b?������?w�ga\�����xr�.f
���7���_����#�=	p���P�*5�BH6sJ���(�J������r��>� ��:3	� i�����uON
�c=��n�.��) 2$����z�J���Cޮ��ȅ�ۺ���ֻ��a{��"�/O����r3�Z�Uǻر��ۃ���J�-�E��h��û��i��54��X`V�v�vJj�(ä ���⽵
��t�JAJ<�V�I�]T
Y�F���n��9<����g�o>�|﷽����1��(`����Q�7��^��~�6,�i������sq����A�B���d�0y��9<�I��@}q��Ԋ����|����R��6˫fcu��A/.i����L��ܙ:�㱖�P�?�Z�"�h��B����b�<���H���C4�p����f�k��<������˖{�v]��r�Y�T�Ky�UʙʉqY�fT�ث�Hc1�{�0�z�뮏�� �_��6����pt�XVi,U;������te�H�c3G��!��8�""=��S�Q�TAƱ��^8�w��Lu<�\

ȺF�g��{����E'�8'��{[�����p������}�|T�c���"%J��Zi�<�Ï|�_���7�?���c�7@�,j5��\�Jɐ
��1W �,^�4R�J'>�RZs���Y�pι��W�/q��4jm.8 ��]>�rr���W�pS휎�� .߼7?�'p�'�`q�vDUse���s�M���5�>��0H��s�m<\3��|��N���Z�G��7�&g�MX��TR~T�DfOzڄ<�T+�WΠg���\Hs��v
�d�D��px�\���p ��m�/�b�l�6��1NW(���W�KfS�&&����}<��t9�$����Tg����|��M��DK"�b:�2)%��M\r-�=)@D1���Sb�D(�#�C[�����hٲ-�P/+���������D�1>�~5�;j��	�����-�����K�����G��ޝe��Lۻ�#��J��c((	�SNY*�i�FR���L�9�����hv���iE;��P�!�����Bn�~�"�L��2���@a���9k�����YGH�7(�����a��`��S���8��K�����)��@�`Y�.:Y�+���+O�ș&�Aed�����o������_�=�2� �����2z����3�}p��|<���o��+Q��^C�mrc�x��U��&����=�N5���)55y�6h�h�QR�h�lh�	���n`�W3�+�����.c:��j��d�*顑(x�t�8$Q�,�G8��')�l8]ؚ<ED>�A4^��{
�B��)`Ch8/2)�=� ?���:a�sW���!��>��m����W�.��7veϓ<)���M��Śr�Ϻ�RP���`�'�ۅm�<z�L�N"��z#�+@!����k�����&�3+��A�ڽ�	\j*���A���z+��[`CI�
��Y��̻�����5���-��P�4��G<�Bv�$����a6*Q��el0���G��6>N�<�PQe�y>�ꠑ`@:GR��i�#7�������^70�*�/K��A}..�����p���p��mh.8���Պܪ���w���ܩp
�;@�Q�χT���%�j8�'^<U�[��;� �Ӽ�x�o~1R�y��6�ؑ�N�Q��& ��^���lX?PLX3Z.��7_�?� �{��`��W@5?�������\X"�5��AC��qr�ц��)�=!�u�\��J_� ��Hs�	���0K��i�M~ln�DHu�`L�����������AS�+��h�a�_%�ke�t6-�x�5�<Y�7\��~������^���<��k�&�L4'&�|���?������`Y�yaaC0�����
Z\Y�c��fjPV�D�OE:dI�
�h��0��R�D"��m�aa*p��'Sop��=�lc<��9�� ��=�����s�8�י�/Xjo4ݟ�;�V|�f}�caCe�a�;�U�8Hg��y*,�(�-o�����|zѾ�|>��?x�!����.�+/ȉ]�f����!�ԭ��w�~���S_�paK���*v�B�)\j��zG~9��T��>^˚����xI�ȣqd�@��1_PE�h4���"�7�_Dtc�:�z��
iJi!����Gl��D�`�r(#wt,F:��jɢ�5��C���~��67�+��Tx�EyA�e�� :�nca��aE�t%�C7�e�1���
L&�Ov�(�+̷�&����g>�<c^���C�B^7Ԓ����(�w�����I;�w�d�XsZ��X���1%p!ݍݥѮ���(5,n�[_s��]o��	���E��� �F���l�������|�鶬�:ik\�����!7����^>C/�{9g����V��`���r�N��(��RY�`����-���p�����N��GE�Z�=��'�NgDե���~�����g����0�Xò����*��4`�'zP��]���qQIK��7���V��"p(܊=a��(U�T0)��Na��^�-C�8�� YB8��o�\��c�6���������ٵ���#�������d	�U�эb��w�4 '��z������PPT�н���!a�����/h�������D�w��^ԫ��"!݋���+������m����7�Ld��m^i_Ű�M�L|��]��z��m����~��aq 
�m�0kӼ�-o������4��s܈���	�0e;%���p�aÕ���AHF���;;�Fá-�;%���uമVXi����RR�sۀ�q�ʘ�1�9�)C���b��� ��_�º}�7wL�Ʈ��۳T�p8�3�lC8�!{OGy
!g�gee�0
,
��0�"EB*�K���9-3*��bC�,
x�0~5���;�[�3����Y+�Ë�%���x�[��]��+���D���������w�_y���~�P�C���-������f�1��Lq宇����V{E`�E�6(3U�y�,�wT`�8��x 9P��Wx_��a*!���afX�|VH�8���cc,ʖљ$v �<A��	#��3�î����|WiփP���y��BY�g��t�G۪�@W��!|^��P:}�LU��񴡏?��u�g���l]}�+��렁��-�V�uo� �[�6$�w��P�0�ϣ��5A~'�/�^�O�UCrciao�k��Ѝ���ĊA9Sn�i�Dv�y��;�Τ�1���w�C�U����6���r�4�~@m'��h���ݳ�������_�z6o˫���~�Ճ8���=Tr�/���P��F�&f8� ����A���I1���U�
�@귧XC9�I�"�"gmM�F6����\:>��ǿ �?�)�ݺpx'jaew�=>*\7�c"����e����
B�&� �o�Sw8��T�@6.���Q�M�.k�Vׇ�#�P����gMH�na��UPm�3CN��-a��/������+�k��q�E)�ai�z��'��G.�h�`�3!���Scj��3�cA'FVrp�J��$���c,�$
�X��y]�,��������wlg��T���BA`j�v����5!�;�,� t�+2��@fW*��68o��+&.����̓va6w[�}�����*hM����{t�y_��W�+�O�t.�8*D�0�\��J~���̤r��NQ�_��8��s������u0�.;|�ڛ��Ss�vą�˅���xZG��v��h޺H'Um�g���5.W�?��9Do����}i���,��S�X�v�o_���_C�R���ͪԠ�q�|�b�*����d�>��!n���q�=� �D��T�HD9 2���]W!rC�^�[�h}�ʑ�	��-��VƗ9aH�B%���	���_.�5~�/M�S��6�=� ���ᑯ=���
��?�Q�cC\mK4��Y�����N�𺻮��X��S�m��+ߚLk/�ig(��xI-d#*�
� ߧH>$�������E=���0wF�Dt1!s~PQ2W��iq���9T)pԙ�v���+a%��+5�㛽��Z2f!��W�t�1�r�ɦ����+77�C��9<DW�	Q!zR�FR�u�:�;<��&���S4��Gۀ?���ǖS��S��⽪Gߘk�r��%��+m��D�u�!,E%Rtɗ��=���8ޚj��i�w��+�����B�ʺm��S������jL�IƵPh��xF�k��#.K��F��"�ex�,��մ�*����f������=��ps1�,M�;Pk~_�/�w��.򠑃,������8[go��[�\P�X���#����`�m���5;q$ ��7��`�pD^��I=�8�1Gڦ����c���g6�������T�66 D��&���RÍ�>'�|f/]��6����q[@E��a;�X�Dސ��ܧf�\�����9ʁ�NlkUlMtB\AT����"]���u!��Ý��0��7�g�~��@���q�P>�y^{��j��2�vn݄�ٯ��aQσ����������Rqj�Oao�Sri��i� t�˹���>�\[!À����b���"|Wi�؆�� D��ޅ�����K��x�*6���FK���cp)e�7>��[�ŋ\>?�\x'6�E�	�d�K[}p /��
T�oے�מyg�qZ�;+@�A����2Z4jII�HC�-�b",G� ���mk�RX��O��Hi��JgGv����EA �����d�\[��r�� ��6�ѻ
%��)�I}C�]r�xӻ�-󬍹��R}��%�e��9r��ṁR�J����o�s����Q��� ��}c���� T��
�`\W�I����RCj�:���FAV)�$��L���I=�ñ�Q8w"���Q�
�FY�~��������������M��VP�B�Α��	��V���nڰ�z^�=�b�W��:::��� ����@)�txI ���:�©!�60�9���X�d�,UK���c���c-�Ń(9��ׄ�!IT�g���Zy��!�J�#��f�Z�`�f�F<���]a��� �;��t$a�H�ݵ�6������|@e�
e����`�@��Љ�䝇�i��m:��z]]y�8#�qF2J|ӵL %�G���uc�v����@�Jx�J�a��ެ�ix�r�~_r��&�Gq�@��Ԑ��q/�j��V"�9_�u>�ɸ�O˧����RQ��l9�܃��kT��� fQOkȐ��^d�\J!)C��Q�9r(4�3���M�F7��I��0�c2�{#��k�gp鮻��9\ke5=C�Ƿ��'���x.��4
zls��"t�/�~G|��:�Ƿ�p �Ѝ>�5ļ�7|N�D���&
L+׽uqb�)8��n�-³�2�fP�0J�.��b/=�i���O����3�[�Z)�M�Dyg_��5��H����"��S�$tR*Y)�ɳ�i%;~{+�L��*I�UlR&(0��Ł�g��FOR���<�[
�mT�M�ڤi'G������]�{��5�j��%u�ư�7j ����] � ,�_�]�g��g�xǈ8\E�P?y�K+�,3�O�oR��Z��5ŀ�#�`�=T`�V�hvd��f�s�/�_�{�x�;� �s�?4p��mx��-8<���،7w�8c�0�y�͛�\�۵|�]𑤭���f�	5��M���9 �:@`X�Xg7U�����%g6qj�N��}�o�+2��QR�V���=m��L�$Da��>QV[݅��6�7��	x<)�E����*�B�9d��-���a�tz佖�ʊ�!�T�LP �$E�T����� 6Ȳ�-_^�H˖�o4<����/����_÷�e4=��:�k�mY|��o��)Pm���X�b\W+'j�y*hcu�u}��rcӉ".��(20����Q�-��H��wlL
Yߣ���A�QIy�(�X-YWs�)���]�d�0�R��c%F�4�e,'��TU���S����(�R��a+��Ǝi姮��u
c�,3�N4��O�v`Z'�^O�kU���<{;PΈj�2�7k����YG�&e���!�τ���5����E/�2��mD���fr81F蒧��c�� �`�r��(�B�Ȋ�MT�c+* o�%6Ϫ7z	�n��̀ּ���_���@��Cõ/��Y���C[�����,1��)��|tЭ��A�W���hRl�v8��87r8E�Ln�D�+��쬰M�3���Ɯ�p���v�1g�M휀�� f�%���n>�i8z�p��M��
������^���T���V��ck�m7XO^�lLs���C�Wߊ:I��e"bJ��F�k�^ӉK��_����;�cM��F�:�
n~��P�Kpᵯ�#��D�m�!�Β���e���9Sv$���Ġ}��'��e��ҌŝǦ�zq3u/�b�D��d3%�6�Z#�%S��I��]Xte�-.�Z��Gj>��>��~�6�5����P�!W�=]qM�vSx����>6�����b��2_�a�~/4���y��'x�,֭S�SPA�,(��d�;7�߼�WU�1��汙�F�~��Ӏ}��;j�.>Ww ��=�uNN�	�ʢJl�N"W���o��kZ9�l���I����T@EQ�JA!��3F�0�Dɴ���R^���Z*;��&Hz����q��Ac~�p|��Ͽ����8�����M����S�n�a\�_��>������J����QGe�W����D�����T"F�!�KD���4�;Ҝ(xu��%�du�&���_Qw�e�bݺ&�\uq �h�^�@$"�(K�nrͥ���i#��Ό�\f�it㰁���Έ{�,�,4�1d�e�MGL�V?��20��3�i��5�0�a�m���FC/���?�㚐�?0��W�<)1��f�eH�Xen����!AJ�]S�=?�QM6�E(��
N:�|r\��"��'�Z�?�i��7�L3)��/�}��j����7�M;7A�H( �?�r�$M�5�����e1�9x(�$E��>By$T��Z��9C֔)��Tk���6B��K9۷��g-�6E�[7��C���=n� �Y�v~��S>r�rc7����r=���M>K	0�n������2Vt���i�(������p&]:�,�N�;o0�-��}�ټ�� �n�]-�hʞ���G����U��tɭ��l��$G�^B9�{�B\MWeDE*P�Dg���U���B�FP]e�f��-,�]2��qE���' ��hE��L�ir��V��S.����g�>��&�LY�f�RO����7���}�Qx�۾�����K���t�%;��Zç��Ux�hաI{��}���1}�ʽ#9;6ʈ)��1h�<��<��|8�� ;A������2��a��+Q���"��NM��U�f.ǘ�/�q;�Pr���J�T$����y�����!G�;a�Xg��{�@0>���*pʲ@��0
rV�w��Fe)��3�\M�����w=��Zs��"*�Oz�{k"S��2zm"���-�o>���?�!xӽ�������q��0o?g3h���S�;�~n9��W����Q;H$M0U�S��$���sj��9Me*I/ݝ���ĳ��F�5�(����8je�O"��z�]%i�5!� y���o�u,��:d�-C��:G$b %Iq��*��㗓��6d�ƈ���w��y��t�0V�2��mA�y�+b��7
S˼}m[�Y�ŷ�g���]���0l{M\�ߧ�j��vE�~�~B�x?�N�/1�,;[�����#O��OK*4���*���1uѨSV#�ǃ��f�Q�#"8�{�q�g,_6K����G>��������]��P�oL_��F�q���/�^iYU��˙�;R.�gDϜ%XJ`iۥN�ՙ�q��*��Jc�*U)
s��F[�ꐋ,�{'�t����l�@݄�<�vM3�9�����7�� �~�/@]� ��cn�DN_`e�
�KW��ӰQ��10�^m\���t�_��P���K��[��3)������8N��:Y�[���*9m��L��hw��:nT�+�����3*Lf���5�`��|�i�O=���f��4
*u���Ǘa����ORg�����0#�k ��@`Lu_نU�M"���Ql 5I2���{�8��A�S�>�>����p�Ӿ�a<:���o���-4��/�M_PV��i�G>�r�W~O�|�h���I�1J�Z66��������?�#����v�[_p٩B��~�h�.��x������0,�3�aV`a	ēo��!��d�M���8!q죠Ze�F���W����BtxA��S���f}�s���90�i�Wa��i�<t��c�-�>$��y�.���(W�p��m$Ы~J��]�k�mCaw�-�)]�M��Ǻ�c�%b�`���f����=�K�������H�Ǉ��~:�5�r&�'�$��ME����9i��_S�@,O�w�秡NMÕ�(�K��('-O�\+w�ܯ��g~�^���_��kƧ���|~�����sX�j��2yE�U����4Od��8���S-'J�H.��"�,I�9����Ѩ�^�A��>)���YYu$M� Wm_x�&�u�d	4��D���,u,��mB�{�|���9!h����XM�:_��^aUF%?=�N�>�MA��.tN�����RXE�J��g~]��~���Aһ��yK�
Sȹ%y�Ҋ�[�k��%~����ܿ��X=4���|1"�Y�1z���ChZ"/����%-�U�54ϣx�hj��L��֚p+A�m0~��폌���i�A-C�f�&��k?�����F���E��l0XM���`̺�t�pOj��z>����u�}T�*�eC;\�Le�X�z8<��~���Cü�˚F��D]�Q��x�9Mi�=��z.K,�` �o� #m0L���-g�Q!Mj�A����C�ϩq��Q��Y)�0����{zV޹�=�	�qc�tc+oZپ�.����_x.��%��}Z9�#A�b�8�5�V�[1�T�Oʟ2^JG�@���'����������� ��KQ�RX q�R!w �֒�����މx�E�*G�  ��IDAT?,�&�k�h]Z.����{�{5�u7-��ȧ1[�i� Ud"Kv/s����#c����� Z��()A�{5�����D�
<Aynld��}ܫ�є2����Y	��
I�����f�Hi� ��u:&]�.�x��{1?�?z�	��?�3��a�̢���M�+��?���?����W_��p־j �{�L��2P�r�L0��ӷa?�t��y��u��AD����������)ok`�ΑY��iEd~W��W�
���u�9��&���	ga��)0������g�
�m�J������1ZX��v'�(	�^q�Y�)��f'*-�rt�6�݀1*�� 9	�}ɂa{u����U��5,�:��n܄��W�O�?���{��V�|� �'�ǟ~������:������k��/@v-��z��C�7��XH����w%z�������4���@w�vl�ftq�/*#�۹[�ωˡ��@�S�t�
ϣ\������c�M�bD�2�] �8n�2J�K�)�T�h����$������w��&h��t�l
��A�u�]%O��d]��x�s�+�Jiς�z*@H��it�"����.��,�9���zE��Z(�,�+�7��Kx`��g��w��Y��D���^��ἁA1�(5}��"�ˣ������`"���k�����.¯��G��}=|��� �D?l��ŞBo"cd�Y>�E��| �/���u�>*;��Q��h��g8-1'i�(�W �D���QNA��p��'�y~�~�1�$�|�A���p�����b���9P�9,�\k���r	��>�}�	8lǕ�����1c���U��/�%�G�Q|ʛBY��3�t`��q�����I-�.Dn��S�)���)ܾ`�&��D��=�cN��j�i'�p_y
.��
���=v=~F�A�C��1���߫ +��x�=[��_�uWf/g���914!�7nʱ�3�ڏ��"��L��{.�Y��4��E�TC��8� ���<�B����Y�	��pO'ҁ&T��.���E�_�7�e�w������U�(�^X9�᠆�n�/|�7�C��<����ye˩+[��
���\빒��w�#~S��s�ǰ�����cu�8G%�.�\��Jsy��^���.�0n�ԝ��p&����.	�w2�g�;������j�w9��Xt�^�0�9�.���9Ug�Vʤ��p��}FYK����b����O$���]�u��|�me���o�/���W��Jx������\_��r~h�Z*�`c�Q��#�/���3�a#k~�Q�7�N:i�$��g��:��;"H"Ux�>�"U܆4(�Q2i�K#�7�|&'ʼ>K��b)�t������œ�P���S�6�&�<�������F*?���9����vV�~���iɉ���N�h��u���z�� _��t�`WǏ���Z�w&������'3��`��Wp�#�FiVt��*�W�*�� ��9�ԧ9&(�1�E��U���޾��*l0��Nr�j�s��]}�%a������?�ڿ���g���U�u<���CQ�ó��<��W���_��oC}x�L���{��M6@��g �!i<�f�M��l����r�E����jBDǷ�/M6�?GN���Ȇ������ҳ6����XϠ~�x��~�9k���CY8�0�ў�����������A �0΁c�oׄ^Rǽ�#�z�2��	-ݠ�Q+T�4�L�ybC���0K���n<�4\��~�.^�im����n�q�Q���B~�a7�eZ�(�ڟ�~��2W�u�� �I����Zp��e�o~��N��&�7
>e�(L7użs8���C��yɩ�`�Fw@4��~~��b���j�D��K�ks�P�,+��_�`�<?�c�W\�jѦ�0]Wp�Ã_����;���_��]���'0�͵+��N�!�P}�����o�rA� OB=���0d!�s/��F�&幧��Ū�4S��;"ú� Ș�M�l�p`���+6�0v�Q���2�EXj�~�o�p^�N����ٿK�/���w�v<��.9M��\�vY��y_��蜔�+�z��g�Yx�j��fD�zXX��<hY��1�I#/��}c�r��/����^�G��"4�f�Y+gϬ,m/�ӕ;����L(7Y��/qޠ�*k5tw �fWOR��e��e�(�������:}�#2
����X�h��&\����r���pHˌYR��sŏR!2��,iK4!��폞5�ÝK��Cd%y�?��wh1�qa��9]�i�m��ۂ.mh[�2;�?��x��l6L�}갫�����#���*rm��%X�SL���lp�rP����=�\�!�w��_$���d����ߝ�'��`6kj��Wʇ{���� ��_����^������}�|�y����K��{��_|\:h%�E+��k#v���[��I��>����cX�a�V>;����vtވ����ߩ-�@Y�=��(h��M����<TM��(��6�ǥ����`� �Ȟ��ܬ��M�0䬟�yf��k��a����Kp�3��Yz^[�iUyF{���ףlkO��<aܡ�h[Y�Q� �Z�p�T�^(O����`�n�a�yBYo3�!,"�RD���`V+�0�Q��j��Ɇ5�\ؘ,��ի0��2�T��6e�"�DU�+z?�N��;p'c���'�&)�0WO�2�T,iR/���( �ź��2����p�%�E4_� 'X0�ջ��%F$C+D���'�h[p��|��d����Y�q�3꺶��E��\]*���= ���>�����UW��R/�����<����7n�hy���y���]e��'�a#m�kc*<��`�2<�P�KP�qx�R��w�{J�G����2��1�i������$�h;��ް��?{4�ѩ���|��]�M(�$�d9���}�vQiA!�$�Z�ȕ'��B'�׿�{]`����a�LQ��h���_����q|1ď��n���T{Fi�|��t�����Y�|r%x%*2:���-�YJ�������wd���*WQVB�	���('�ߪ�3���������놏���nd/���(߰I@�]ʑG9Fҙ�ۜX�M��W�sд�a[���R��KH>4���:��L�Bܘ�QZP��}�k�}���:J��c"K��I�6w�%�r�u�+��/Ln��q��>��r'"��X�@��:�����P�nG�g՘��?��⟅���.����yJ�p[��������ٺ�M�NK���z�ӄ�\B=t��}N�Rv����@@��Ӂ5��V,Ys�F��eK]������79�:��AT%y���a�{��O���{��E饲e$m�v,?�ˈN^��J_RC������C���`Pߍ|E,b'N�7�aUY�ji��i�\�'n݂��?�����V�k>���%|��m�������:\;>�f~s�l�V.S���TEd&SIC��E1����pIT��y�߅��07F����7�/����L~u�7ǻd�w�3�9��#|jHf�ãuK3ځu��	=���_ގ�c�_��0s{������`��_�2�iC���㨒z��0ʁC;k�h��"2A\��Wl�k��\"4�4�3I`L��cڅ2�8�^��g��z�"#�I�H'�N0���YŇ9̺�.�9H �KK�0��.��Y��� 7&��1.q�瘧r�y�-K�FR��\t:�Y�aexR#�u���
�i�'4����<HF�B��	�fi����
>{��쿽�;�D��l������\����2#�`�y�OQ�Q�kP&N4��0hIX�U[�*|Ʉ�/:����2#���z���P�b��Φ��f$9x�!���ª�M�Ya��9�����r���^Qt�!�L�R�}���w%V���8.��i��n�K�C�O�Y�H���	�`��b��,yw��o97]���B�5�3e/W��"�z��|#��M�F�m����"�`�U��ٗ+חsj���U���8B*/u0^+��WYRcTfU��7R�:���2y��򫈝E!�\�����8ITHqT��zzQa^r�Ay�� ?&ӊ�wr6�(�j�+@n��Ac�iNG����FpױJNr�"�$���1A���X������x�s��Y���@�9���T4��{��|�����I���6�IШ��;��=l�Ϡ��)��m;-JǤ��ƒ���.SAw���'�'e1���gp]{����;���i,J9��Я2}���(῰�#��2��R"��'u�������}����>����Ϟy
�����4��l�~����p��5��A<���.�4C�G�� �E�cE��O�k���t��\^R��2��U��3���mvA��Σ��"�r*��Ml4�$�u��o�x�v�1�A+���̗�?�C���p4�aV��u���6v� qT*�S8(C'`�6��&�KI�.����]���i�qW�����kܦP(I�O�D����ߙn ɾ$�UIEB��� G_{�ܾp���y;���mCoaTPoM10�Ծ����������z�F,�Ʉ��j`~�h�e~:~dk�B,�b����aHzH�m�c/F��@��g��Fǫ*��b5󷱦n�fR��aB#7�!1��̍(��f���x�i�ۅ�G�0I�Ek��;,�̉�}g��⏵�"��)��n�=QV��p(�0��*���u �C����М����
�9P"�u� �ȷ��4�x� K{�q؆��t�,=�Ý�fm�pqڼ�&��;ݹ)�9V;��G�)S!��K�O���d�vv�'���Yw��qE�ߋ�vE�$^���n��+��Ә��@?����9
�$�ܻ� D�b�9(t4�9fh^�ĳ:Q��w&U��2������#5�w �X���Dl
Q)R�0s��dJ�M컸硒Y9YZV��2=8N2�|H5���|�ن�v�9m^w�9'!	}8�ֱ��'+���-/;g����𘟼��9�����B��UY�5�\K�����`�k�ɾ�ho�l�|1
@n�%`6�����2��X��!8>�H��]A]5д/fm�����0F��,��G����`��m0��̱�1��Y��Kp�e�'9��Ut,gl0�~��\�E.c���.�H�[
�0�^:7wK�6}�Sȵ��ւ��е�� �v�\~�yx�S���W܍�zg"����Ɣp�5L��'@���uJ(�
5= 2�U��W�@8�r�������i��Mĭ=~�S���<{��Q�.A��<̞�z5-�!�����Sx[ac$�y�o��̳tI����&,�Z.�����'(]�5/s��!^���jq�W�Z���ݩ��Қ\O�O���,k�!��C��#�Qs�S���~��E��~#�`}�� HW�\3�C��$8��Ϩ������%�ܦҵ�n���~	�	oMY��(J���(�N��x�Ұ��H8��v
��c��9�}#����s���S������y��6�q���g���T�,/g*ӞA:��=��q�ٗ�0�gyu���w����݇�~��}X��f�E�D�U�"��C��ʡ�9Q�i�t��f�ͥ�S(ƼRf.��c�$�TB$���)-K�9�e6�)-'u���CQ!�Wߜ$���c9���&A�='f���0����.X�7[�<o�����`O�h�1�r���Aoq�ɝ��/��g�E�,*N��D�?5���y�µ�L�NL5(w��x��ߙk�����>O��hpv���z�X�@nm6!_�q|	N
��k��Z���+o�i`f>�����m&J����/�O��b��`� o�Ѵ}�����L�K�����`�{��P�6�B�e����F� �Uf�!�y\
�c#���>�^�B���?U����_{^�����_���y;fj�&�~E��jqk<AM��ʿI(ٷ�z�h�i/���}1�
��W�L����<��"qa�L'���Iƣ�$!`��E;p�c��ԓ0���p2S���h�x�(i���8bݐ|�Ѕ�<dѐi��u^�4�]Y��1͘�O��f���(JA�M��b��4F��B2��bh�M_����Y!r��*�i@�o���.��h(?LZ�gz��Pa����Y��4`U��T�-�O0�$��i|i[0t��t0� w쀖�����~^"���%w�ʣ=t��n���[�ڰY����~w̖|F ���N?���)�Hɞg_NRC��O
%^���V��N��w.C��	��N�eu ��P��]�;�6rC���z��3�}���'�'��3����e���R	B�Ē
������k&�4M�YEQ��C�F��*[���R.�pw�ƶ)a�A���� �[]����u���<�2�ڭ��k��v��Jؓ?�'x<��閖�73�1������0:�<;�͊U1[@���<'(r`�P�z�p���a1;�CYRYW�N�%(�2SO^��M����$j�62�#����ETXwM�p���u��)� -8;)mI@�)�["Qr]����bJ�K��*�����"E���ޤY���@)�FB����dڽK�4⡒϶��ק.��Gu�k0�͠Q`nN1@�	�C��xI��0V������p��Ы��+T���c=Mp��o]rpPo�
�Q农�P�t���nڶ��V�d�ji�P��v�~�+p���
�=�!^�b�����0n�B�J:zW�F&��t���:o�}����I�҂�^�ŗY�:�	�7C�!�*:Vk��T��W�x#
\��bz��.��N���J�2��O�f��G���L��-i	�F�~5X
���U>�\��uU��T�%ǘ"�]3rs�3)�xJ��il��uR�2- �E�V*�*���&��7���:�F�gvl�2�}��Q���y���&a�m_�ۆ]P<�V�8˃��u���E2T�2}���ۇ��r1��J���kȘq(uA�BI�� #��*EӐĴX@� Ҟѣ�
"�������u�xy��W�E~s�s���g2�`냏�Nr�!i+�s�TL�"��
�FCp���х=�C�F	�΃���s���K:6ƎΒ��� �;l?��Gwǉqr�����������^�\�C#gtX�l��m������];)��뽼����\�ĝ+�bsPy�a���m99��I� 뽼�z����b�bi�Y�z7H]�.)�LB���o����g�(��o���C���D��*إ�6�R���}(�4�V��KzH�|+�`����am#jp���f��}
�:��Tx��	}�wW8�P��0I�wXF:%O���`�XKD<T�+Qk��=�ƴ5��$�ȃ����R� ��)#p�T.2���bX~�L^7��Mq�
��x��\1�t5��]�+k+��kh�W����)(�J�8]�J����\��`Cr�1ҁÆ�`K�pP�s7 (A2h�&�K5��1�*,�"�?o�O��#X\��.v��o	T���t��C�թ���[&q� RA�a�v�Lab��""��Bق&@�B�*XՂ:\떶M�Lq�y�9��e8D��~,�K�'�X֖IwO�{��wb�\��r�Ǎz\����I�l[sϋ7tU��C�2(��l�NDK�Y9Xj/G}� D5I�m�w�����7�wU�v�a[Ħ`WQ���x(	c�^ɘ�C� RA��m�*��)�Wcq�Ҵ�KD�4�2
@���b;��+FR@	T*$Cq.�7 ]�*5����_����"Y(%��Ge	�)+wA:.P\Q:�Ƿ"��{'��bHi�����ص��P�-�'�.�T2�	C��{8�0M��e�=���fj[��Y�Tm���. �U��a�����Cy�@�
���*�t��!������r��H`�w&Ϡ!Jڤ˯��SL0� �W��޲�rf&���HA��T�� ر4ՔGZg�V-	$!O��;䷧Qޔ��{~U�my�X�o�v'�8�lŅ�u��e�hS�w�6���:�7���}t��5x���¥��������w�F�.���N��>3gP�c�h�ҶqW��E\�;p�SlS��<�Ʌt�Ɍ7���v;:�ŵ�a޼
�8`�VC�����w��"�N}�(�Kej�ܩ|Ǽy .𞕕�Ɯ��M�C�Te~�r�I29T�DǱ����as��b%Aq�T(�zR%�"as5�� =�ҔQ����3m�ʼ�)��D&H�q�V��,�����&n�Is& ��:k�vrL�i�R����=lr������L^��_�	w8�"�Ul�d��e��{�D+��>�$;ɔ!��g��W��A�iTe�Ћ��V.{��C� �7��ˢ�(�����Q;9�?.�y�շAa�?��Q֡� ����*֚t�.Z5lN��.Q�S��M):�X�}�a������I��S����	fnÜ���k�	�H���mh����$@L`Ҭ=��9�"]2��m0��̯*�`��#ZT�(��ddzy:�(B�Um0]yzm0k�0P�K��)���������6�m0��D���-3��R##�f���P�U�6&br��吵��sTOe:���N�Ae�~yH4O���1�����sVl�ecB�p�8���x�I�U�Y�ܝb��(/����{��a:���g��/ uJ�3���ĐT�$~n
R�����AG"���B�"J\�2`�xh������Q�Iͭ���nAd�n�u�eO�6��%��b�G���-�opF���K`�����8��0X�I!(�� ��u�tH^��j��L���a�EE�}6XW*�+0r:Z7 �*䊌H䒞6�j�)�{��=>_Y
-A(7C�8C�P%��!`��%�2o�R�P[�n�����8���K����]dr��%�jÁG��./˝7�ڠC��N:��S����]^ѱ����/�U+�5��V��ZRf#C�o��rcS3%[T�V��Q���2�~�x�iT==|V�J|�zJE�M��3�O��F�zt	��$EQW�fR����?ݒ�J��O��SU��b@��B虈�h|'$.����Q�?��:!P��֦�=u8�����sD��j(�R�S�gE�2f�u��Ω��)Kg,	���%��������Z�L�T�e��|��s L5\/���n�K�"SKu���~G�wdd�Hm04#-;����It����*v�!i$��[���?�<�������]��R�/M�'v�)G�H��Ғ����.9�u�{��W�#m0�I��G; #�R�Y:C4_Oț1;3ѓMYԵ=�WQ���ڷ+�1�j���£p�n��ڷ��W�h��v�(?��s�� c�ˍ��@�,���������#Ƕu���ӒDl���
�(�`�=[�*�.$�W��EQ��}"���������7oB�4�)�䠲}&g�
�߶,�a�bJ�xY2�*|�����P��!#��2#AN�T`bC�OsŪcZT�)�s����핟�4 ��!@�k�]8o<%c�k|�X��j��ZSf��!7b�3�r�� ٮs�wBQ� �_�ۢhI���k�O,@���������v �5�+���X)u���!�U{��iǟ��\�����aҐs¹cݲs
%%�*��2���6�L�����ֿ�г�Z4���d���$JIWP�x��,#����AyCVi�3S�3��@�ա��"�b���~�"yVB5�����GJ�$r�B�Yr"T��5!�	<~L�
=/39E[�Ӏ��*nŢh����9�c?KE�`��r�x���̇
�d�*w�9�NY�i ��(��gN�����9B���Ǒ�9؅=tW@�z]%�U:H=��� ����2�~�'(2���D��)��赪]�4�xPT7�:�	�x����a��v��ҟ9~`\�%��3*�HFr�&F�ǚy�>������Fj��l��mm۶<���	⫢$�@����s��&����^\Chٲ�.��`(0��4��J�)>��;4@�9(�x���5�W;"�$�K��uc���o���V�B�l�}���ie���n�z�p�li3Ӱ4;f T�M�ҽ�NN�`��_5����T_t�[��j�a��V�S��ѷl��(�}ĩ�I�(tt�Y��U���lA�mqU��Ԧ��f�n�lـ���Q��ٙ���6ڙ15Mc��� ��0Ȳ��A���1�Ǒ(�F[���/A\��I'6A%F�D:�I4�0���������Q�K��t����<�qz�X6Y�/���ǆ��w�Nrc�$Ú��]��)e�h�}l�$��i���x�ε)�@�FV��
��u�f���#�k8�����l�z������M��cD�Ek��qwa��Jȵ-��*͋!��7����d�g���<��m+Ay��Cp];z�'��v�-�;$}VmI�a�_��%
���~����k�b���v��GtwǗ����/Ɉ���ڕDht:��Wz
+����A��<���X�My�5�}��(;%��`���Uu��4Z���Js9=���%ڻ���#�fg�@/"��.ĔT����O��9=����N\����M6���)��U����L���h��0�;�����o�1�ȧ��~Ig�;t�:R>�v�d(o�
�;�>"�a�U�l�u�����v�S�/KA?6��9֍]>߃���[��uW�5u���#UUyt��8��l����
7�-c|�0�se<G�o�2�=e`�k�y�ZAs��[B�AƜ���u\wx�B>aԼ]����ـ̚L��e�1@�s�<�x@,O�_�{�2I��8#�T�Eb����t}��E�+�sK݌�H���Fu����"�:5�[UW5=���ˆ��+s���}���Z4�}��	�Am�Is���Fߨڍ�'j��P��)�Y5��N&��� �������t��_���m3�(��J'��T�B�p�s:��	�;%SeB-����`V�0�7S��M6�r
۰!z�����l3nda��U��H:� ��0a~2
���l����mO���C���J�4�B�C�r��<���PF��f��0:���E�ÎoCF@Ǩ@�?��9	��S�:Y���$�*�� ��<���M�KI#�Ed�Б%�L��Y�_��퀣�~j�����/M���0�٫woN����(o�;	�(��^��_�uƠ�x"�}��s} ��~^��!�r�t��j�S�ēv&��V"�v��ra) �'�]��36�ˎ� �i'H��t,�En�4^�D9��_�Z��){MK���K=��4(�d����gW�,ڇq�4P$ :���\�8�� AłB�_����RÕQ��v�ul���|[7�jg|3���;��W�,,J9��vNF��Վ�0�I�<�Yw�/�����S���
���vc�hU�b��p�{����@�������S,%zN Z4C1���������݃2��2��*]���������E��ض����Y2�	�;m \��K��ĈF	 A�+M�$1��X�C�=�a��L��H	eP(?I�^	�i���A[�Oc��U�A��Z8�+�6
�E�Z������Ï��SԬ�תT�+����x�~��[��'86���V��p'B?�/{Y�E��*����T�.��:3���-Z+ddnO��_��\.����|��w���;�D�b1}0��7.�~b�a`
(��l��!\�,
7��@�I����VCvGV-�$	��b(�Yb�ܗ)S�K�l�RQSd�RT�&��m,��}�㔦ES�\J,F7����[�۴5YO��)Q�^2�>��k��?���L�����)�z*�,�bK���a����0Λ�ngt����A*�$lbs�%�A���,����9V�3!~��֑@����N�k�S�5)4܇�}$J�F�=s⸠�LŞ1�C������h@ju�{��4�LG	�����<Q��O�#&(Z1��c0E(���h�+�)=b֞e>�<o�mt[?ä�sr�Z�Z=�4:��B�m��Y_�.%lW��j�u5��.�9����,��'�}�����`�!�)i9�,�I�8�"g5����}����Q��!��kbPpz}<KGUT?,����U��	y�nɣO�S��
y��g���`�%��q dˉF(�PR��4��4/�U޾���h���!��Ȇ�<4@aw$�U�/�'��Qt���JK"ETBv%�	��Ry?;��8��"��b,��ݖ��{eC��'`v�&�C�H��o�����`S;�_P��]�*Ń#��b���^����i����
����]j�nCs�f�자�.@}�T���צ 'ᘉ�Ӑg+a֯�	QH!t���Xj�Wd�������*E�ق���ȼ]B�8����"0@>s�k�z�m�t�Wq�-�;�{��o�9��:��z����"&�I�o�AX �	m�f�ZGOʂ�+�h��"9��p_0�B�1��S�V���w��n�%�mws�3�^���.l�{�>���6W��.3����=v����|�*�M�[�_F�/����8�~:Kp֙�cgҦ�QXPV�T3�S�IH.�HYfF/���� >�յ�酸bS;�e�#�)�����5�{Xt���K�y��Q��?T��ЀEx%�+�V+�C���3�W��*&i��g�q*;R��Y�M8o��'��6��M�ޑA��{:&V��z�05~��w7|�+�=F{ ��{����Q����%;�����9�QPԫ��������Ҽ��h<=.$Qx�]6��!�j� �_��m%�hK�2g �{Bh/�b�6�IThi�	vi���!9f�DK�o�L�VP����'v8){�R��|pf�R8��,M�5��M囈�t�`)"�:ǃS����k���S�8�v]8>��_x.�E���F� ��$����H������Ĝs2��/���"pd6�O��Ua�cD��7������a���M��pV�Dߨa�X�6NI���6��ՙ(|�W��]c���E��p��_ym�A��:�7��OAJ6�&��P_��R�v7�Yp��ؤU�</�>-�7�7�HGg+#y�'Nc1W��`< �������\5R�$�7F�0���\f�4)Az:�*��X#Ɵ�2�)��	�[�y���t�N���B7��_P�������$�u_ͭ������O���ǡo�n��S`�����. #��F�m����]��X:�%%�������VͿ���80�ڀm��3~;�T��f���Ry�OG����J��o������h��)���,�Y�ϳ��.��){�HZ^o��W�|�.���)�7 �����&#��,��p���j'HH�p� Bw���T��9u,��dLTˈ��yN�)���	~���*P�6=�Fi��k#`���g��Xc�ܓv�H�]��j)��So��ل��sw�6��5b���j�ݔ(y��<���_��6
�m�ow�� ��oFg\���|*�5�w���2�H�K)��8��������8��5Ż@G�{�ٚ��j�L�h���'v�����4�����H�4�7V�i��W�K�߂QA���Q�����32�JcB�P����^�1�9�AA����H��>i.�����з\�HW.B{������>����BE�#$_:�XZ(��ح`��̮����e�l?�,��/����n�űi�a����9~�
u���t통�߈��u�7v�8�Vs�B�N�d
M�FvzL
�@�����
ߧ@�:�w���
�0j�[�Ҝ���F�����q����z��3H<���R�nJa�Qqר�}�u��7�ʽh�2*�𯏾a�w�������-����|r�(}�������g"U�C^���FZ���q�pl�P��[�����F7�KǍ����2m�؛���;�T<��i�5yLd(#%G:gl4�K_�#0����I���p���g�]�mۮ��>����ss�"��H��� �`T�Z�h�U*UeY�Y����ժ������W�~bS�UM��DEA�Њ	y%$ᆼ�ͽ瞳����x�޿�ǘs͵��{�������֚��ǘc���&8�"��d���-��]���FW����c��"�e�Pu%s��k���n+j^5�m�C^p݊��K[
�­9z�L�s�;Nw�B{c�!;�c m�`�3�N�1���u`�d��N��9V��n�[)e��^�"�y�L��z `����I&$� ��Rќs�&B���!l}p8Dnǐv�V�'ڋ�C�u�r �-���d�c����:�.�-"R���Z��_�u��)X0v%tm�&y��Te~���|��;����������`о�~��B ���g�l0�+���^i�b��hx�6�i�D��>u�6���`�){�3�!o��W�{?�S���^��y8E]�]y���=��X�Ջ;5QF�Ӻ>��F�uŕ�����ĭ�5�o3C�ImW�}�Гw'7���f}k�_Vt�A��M����V�+
�J�wҜJs�t'Bc�[0.F�\ Z�߂��亾 �'��_#�Ʊ�����l�Ӌ[��.ҫ����U.{��"���S��lYa���,�]��z�e�E>(��ʐ���,���E�3��Z�av�����oF��4��ȧq����=�ca��`��Zϳ�B�0kl`%Jj٨��H��Վ��_��s,<��'؁0���2���#�0���Ϛ��掋�Z\ 6�QkWh�� �渺;��'��d8v��C���l�����?5��9� =)N�;�<X,�Y�ga��i�2,|�z��㠅���X�$��Ә2K�`7�ez)�lXy�Y݈�.��v�3nŷ�ΣA���W��5�cp��N�:��	�F��GŌ��#��x����s��k��iy�|��Ef]
OJ?��x ���Pm��s.�9��s4$:�1�� ����%���k[E܃+30P�������i�^�j��I>:s�D��c��!�m����#�Bs�Ȭ�ťEM�5M}*N���F��{_L��x�ǰF��ʙ>��=k�+�~�|"�7��Uؼ{��u}0<t=��_�M���sVG]D��`|030�q�A���6���<l���i�&7w<�<���C:����ӫ�֛w����I:J�42p`ت�W��VZ$&����������v8�if�ٞU�aA�;^c.�5u�|�J!C��g�M�)3�0����py<cƭ	j��%<:�oBp�]p����ğ`�bƬy�I�gі�n_<�e�HN5���:�c��Z�%Fo[��>��v�f�D>&C?i��Ӡ�FZ��23_���K���,8�U���OH��j>D����#�H:n�Q�Z���o�q$?A�ގ9[�((+���x�&��RT�V�eZ�H/��s��1d~ԁaAda�\6TN�{��;�0�a�(��Έ�p�q���mǬ�vh<�*�E^g�<v���A��p��g�H�9:Pc��ȱ̭�ҩ��9�U?�r��d&2�g;���s��⴬դ��/)l�
�]
�m�9�@6�` л$<������ylZe����T��ݪ�/뎎�o��~�@8��0}˥������ҧ�.����y"
B��DWԹ~�[�����3���z�o�A�� �5����C�w��2�}�^�TM�۠s�pS�υh�f���ڸ��w����Q�)^�	O�[�*�ڕj������ZmL�F$+C!�o�A�|$>���6���`=��0�jL�j�a,�i�hTOi�g�'�l��BZ Ӽ��>�OED�m8�a �G�}&��P���U-�m��H�{u� �����b|�|{#��64��G��t}02V�;v�=IP�������hZ��=�ڟɛЦ׳q���kd�dMI�<�k��n���!��g����W!��A��*s-kIwr��깭qHI�þ��,~�q���*��n��3���C?+��{�yX�᫽��ƨOh��#� �4T(Ɔ2��%�6	�u��Q�5��h���6�������>�{��y��
me(8\&�i�P�3�e.RE]�x,�X#E���b%�����E.U�K>�(�Wq�< ��kb����dVS1�ۉ���M2a���z+k���4xU�i��yQ�C�Ց��";�^��$愕�JLB>�K�p�sN�`g	c�~~�:'�l�)��sھ��f�-�vP�Mt�T;�K*�h}`����?`$�M��bh� ����c�m��`,�$���v�fXY:?/�ԇCL�&�Q�������yu'�=9��D��{_��k\i�*�Cڍ���TV*k\D��N`]�h���h�g0����9Y��Eu�)�V7S��Nk��:;���Ɋ�Lߚ��M}"x�h�\��ס���a�U5괽C�
��*FYU�;�vF�-���Spq���y��6TAu�UoΘ�|��(�^[h�ʔ�I��a{����E�"�iH��zTq�dO8�vԋs
n;�v�-�d�L�i�^%t��.������"}�*�5�W��6z�1�h���Z�Y8��x����������c�ـ�С��� ��c �����	��d��e�j��5�x�*CL��$�jL�g	�Unun�#���F[����J=��0�U)e\F!������C����M�HO�����%?�������-��b�72�4>ԣʇ�>���1X?R��xqb���X2�U��������f�Izz5��u��Ķ�
�������!�y�;�ؑOo�1����o_�f�܅���تІ�:6T]������*����A���>E6�)&hV�Ai���ՙCY-0o�H�	r*�cس�
$x���F|A��ж���1e�`#�N꫓�\`�����*�>����x
��da¹���8&�v���g��)���)9t�NxBG>���}ʩ��g���;�'��������.28z���N�Qf5O�7QNhzg�S��t�t*g��AX�@�7s!E*n���2p�㪌)�1_�KRڐ��bF�B& ����L9�\+c=j�z�U���'�^�1��YK���(A)�.�3��Q��Q�m�����w�i�\>�+�q��D)�A5bv���XMV��+ؠc�b����)s�v7W��ڙr�=gRhg
��%}��=�pT԰=p� �� Ǭ�6:�8Gv�����j�U�;��L8���=�yY�\�s�K��ء7�L��2�|�`d��.�C6 m|R��.��$�yC����"}
�������=��,�����E&J�r�}s����*�h�T�-w)	��'�m���öڣ��5������S��Ic�+�MY��|y1<����`ZlҦߊ�I�P��Kdd�[X��=�$H�hI��vF�?�}�zĶ
��E�eCLՕ���@O���U�]�='�E���$1S���a�ͻ���ˇC˨l?a{��&w���O�玽���n�CZ�����}U �� ���\#q�n��.X� co*���o��Ͷ���1t�9xڏ:s,J��̴��qЍ���=�n��X��HT}L���	 ~�|�SՕ�ȩ��1ȸ7|0X���1���Ǳs�S�����qL9�B��&e��_��2P�t:B ��e��Ϡ��W	���ԕ�=�[(�O�ڡ������K/L�I��O6�JcS�����r]�����:>P�����^�J�6j>�b_z�9
���r	�)<����bҚI@0S�~(h����Al.�"���C|:ғ]���	)P<�|HSw�t��h��9Z}�ٿ��dH�����W�U�kŷL��>�9��(���>�ͤ��s��:�c{1���q�1=Ib4�ּP��`�+T6�İ�g�;�p��[���y��^l�)̲޹uv�yf�k,X��Л��],�O��!���],�!� ���P�H�qFE	��U�C�XX���C��S��5���0�� Ncaۙ�'f	�f�U8eF͂�y�����{�g+��Q#3��c�ǣf!a h1���#��萅�Uƅ�"&3xJN��؂g�u=*,���!�Ր��ڈ-�:3�t�V8�0�M���pR���1t��2L]ߗt��o�y-��r((�Ёԋ�C����U���>@�0�`�C����F�5j��n,�µ��e�g��)ܔ�~M��3;��H��q������>��W=޶k��ܒ�����)H�d��k��:�.A^�>�|��ꢹ�J�Wz��n�����Ϥ��h��\���ؘg݇�E�n���
�3��R$v�*������h�9[͛?�yUF��=1=��-��>h���
\�h���Y�oWW"K��)��0��N���Ɇ�p�lwpP����q R���3�� �=�"�"�c�Jk���M�Է��rB�.��j�PK��O
�%E��/�H�=�,���U?��'����@�ME)H!>>��I��ᄆ|�H����7�>����*��$>>�����)�a�7����r�[as���0=�N��৑���&شx��wT��9��,��7��^��8T�a]����Z����-�}0�y�f��i2Ľ�\f��n�ɑ`��u�t^ng�4�F#�sNmA��F2��q^��U�"\;z2^&��{(y�mZ��;��H�?��f�4����,��}��?�)��򇲹(oLO�
RwKw"�q���J�C�e*pq0ewx� 5������9�cg����'�/^A�����a
g�X����Ȁ|���ܮ�C��a���]�¶��0'@�q��߸�+�htBd@a#�1�s�zTW�7m^�ZK�/�_��W�_�E���_B/{�Af�9ТFh&��n
�H4U7�����e	��}T�u��PE�8�DHө��W�Ą�l�Z���|�����V1r�zS窌��jTNK�jZBep��M�F�Iu�c�B��u���%"v#4�o��>O�g�Ǐ�ه��/<zD��}��������g��E"��9YN�H�K�	���ob����y��,���=jn�I�̷5�:B����D�9�pC������E|o	�^�w`�(���Z�1G0*�n.<y�?IC�brv�1d��\D� #����"�K*@	�[[-��]�	�[�x
%�팼��S�����o�Oa4'2�>	�Z2���v:46J?޵�.Xi��n $��}w�n	em�d�V��S1�[�̘�ʎ���ti��x�_�X�$��Uں4�^gf/�~����;��#����`�wsd+l��W��6�Hͼ�F� [v�;"ԑp�9�֛��;ەX�,�ޗ�cP�~�J�ȅ��X�i�c	�x��W�z�k����/�W?�4=��>��+a�y5�S.W���'_L>y�
�r=�X}1�n��Sr�Ȱ���a�EN[���wA�^)u%�O�?L_L
Y�j��l�M~��Rn���U(�Y�$�x�if�}%9^e��^���~~v�����y�Ϝo�����m�=���Ǐ�s�Ϗ|�Yz�ه�g�����7�ge�n,'Y����� �+:B��6����97]�c�C�"H�����a�|K����|�쪫�t.6���'���i���s�|y��4�>~�,��V����c6:���� 	~=�`��������^�Y.M7�mC�S�"{pl:�h~hG��`/8Bۺ�v�2��s�8�c�O�s8i�s׶�\�	y���'%��ée�}#�D+����!נ�Ij#��=�0��������r��7��&�߾���_��w�+^zJ�t�<�I-���n����6�T�:�C
�0J�����<�#��@f������&j�T��Fh��C����a\pps�ԟ��N�=�̂�?7u��|�����1}���������Ч�ߧ�����j�+��P��o�7��vg� B��(,XeD2ߍ>��`	���9)xj>�b����,��$P����N�$��X�w��w���W�6��k�nn�^84m�'pL�ϻ����*O��]o�P=��J;�<3J�Nu����M�
�3�n��g���M=@[�n�C�94�a{k5��Z�m���8D'��iĭҘA�Xَ���T;��p 5�l��o�X�˜*��*XEuƺ,�m�\p�W=��;Ԯ�� �������g���܆~�>\%=�^�o�<��e�x�-`$"aǇ��7߮j-��Y�8Zq{�7��^&�����{+�g�Cqup�G���������+_����O�{�����Sɷ0=N�u�u�]p��`���6��!�� �
$���l�u|#�>���]*Q�>����������\�[j�U�w����i}��R�G�H���q����O��?�Yz�i{u2f'>Q=��^𪨲>7���)��8�T>Se�	���������>����C(|�����l������éNV:�O��|���u�����z:��z8ͅ��sD5�cצ�|yjS�����?Ta�ݭ'-9(�ss�����N���h�_I�w��u�4Qo	[F�g��nw+V��N���'VB��Ė���t1��܇�t�DX��9�Y��z���ʑn��T8�+��(D��E�e�~q*z����m�]Z�v^@�a�p�f���4���Q�9�"$S�䘮LYo��g����������+����93�:�3�96�ҩ&� �ű�0j�1�V�A�V��Ce@�AQw�U^>:)�� ��8��>o\�����3�{1$��M
����N�+_�{����/����W������~7���j]�c����X�af����(DГr��֍1)��BY�"�A���OS�<�f�w�H��JD���ͺr��z�s���n�`w��w4�1�-���/e���G�n+�w3L�S��Q�\a�ؿ]��C=aj�|�E8�j���~㳩��}��ȇ˞{8���޶�_���|��!� k8wЇ��p��y������P����fFjB�+�4t�������-Lڢ�E��Y��=M��^�ˎ��a�� ���)�:�Q��\~#��P�U�����|9Tr��T��`l�m2Ed�ym5S�&�G��D>�X�<��G��F�ɓ\#��Ξr� �,{-��up����%w��������F�<�צ�9��Ȼ�;m��l��ұ����2b������t�pGOl�$R?�A4'�������WK�i��*ˡ����o������h�nB�.؟�Vu#��oQ�/�Nh���^���Mo|3����Vz�k_�����3|�ElЍy�o�~��� $cʘ����YOm�����D%x�^բ��c������?*�Rrֲ/����R��K5�%�ѣ�饧�|�[髾�5������~����uʘ�tH#P����$��dX��ތ��]m��C��`��n��t���h��t%7A�]`�d���{�{�<�x,�)m�H��k�����+��M��q�������f�l(�n��e~�j#�9�)_�H��������q3��"K���V3�F���{'��k����v��1.GKOf���Q����Z'��^���=�;�{pp�g#�H_:	eDC��Xo��ϑ���mD;쇨�����)��]4�az���S!�c~��Y[�7o��3z�SO����}�[�l�GϪ�0���W�3�5&>�	�9���
9-����@\4h�!6sT�t.?��{x1
���s�*a������=�?��wЇ?�;�w�����U	�J�!�W����ܬöYK���* ���:�6x�E�A�ƭ%��D�Hq��^�N�mώ������a��t,p,Q��y��;�)S�S4b��]�·{�w���m􌡻����M�J0���@۷�Ea�,���U�n3�싛�O��4WpQ͋��� ;�g��ҭ�>kh�ΘI����A��c��w6�4��|�9s���-bsc�҂>׀Q
̸Ī����(*F�`�k�ǋ�B#�i���A��WT>}��6u���N�V!w��h�'��� g�4}�;�.0��5�Es2�1�� �%��6��gs�7؁an�����]B�`�ta�qv[�|Q�Q����]�^�Z[�t�2������F_G���ݚi���T�Hsѧu X,�T�>�(�"��):���G>�o|���{��w��^��MB���꛰�z��KCW��~��]����U>��	����$}@Ч"2w�6y_�`x̪&�_��e�H�I�r�qʛ����z�K����������t�C�^�)!�<��ux_�fЉ���d�S�rF��8=}0���B.���f�,�i����+��M>�ž�T��n��r��˘�ْ��i\�@��Q��'�`�@��E*G�$����5`;l���×��{�\�LS���ڷD��.��{��:���b����C��(�?��e��"\s~"!���"��(��YX���>��ш�� ��))_�gT�C�O��OU	㣾�iY�_\?������7�7���W�T ��O�!a�t7���W���Q\�DAF���=3A^�!f����J��L��&L$1�|1�@
(]�z�[�B�������A�
���+�`jB�o���� �G�	���<��&�^�q��\ňw��Lrq��H��{����.�F�rG�����]R����<7z���2�]��p�w8qL�3�!lý�S�~�0���{W�1g��7��i�����m)�U+o}�V+�M�9�P?�>�sZvh���i�s���m0
�Z�O{�
Q;�����b�E��b5O�"�F1s��v>=����mAZBhu�_����Gň[a�C���|V�?^.t1 ղ��h�AmsW����CT��Z�&z<h[��M�%��>��m�C�2ܖy���1�.d�[��}�e�e��� �@���b��QGjE��󵀭z�7ٖ��#�N�y�z�c%����	�Q������#��O?M��w'���/�׀䍠a������-�#Y(.mɩ��j���O���=�څ�(i�-��z��XN�D���K�)4�����z������Z�ɏ|�V'�����Zղ��	�q�����53ԾJ��>�f�8��J��J�(+��+��rU�XTh_PjwY����<����/X�Pｔs+�������(>~�O�ө\&��|��i�ܡ'm6(�S}�߻�q'�۪�M�T�$�nK�R8�v�h� G�m�ǳU�W�/c��u8�{�3�O���ar�D��٥�����ʓ��Wz$�Y@4 q�E"vaE�����~���aA|�P��4俱��F6�Ee�L�F;W(���z.�*@@AP�-��?����	����f�؎8j|�
ь����R��7c��^�*z����F�2pmu��ɯ'��? g�B
F�ʔP�Y"[cc�P���~j����P�,����vB�q�Ńw��UOW��
��26����w���ʳ/~��)���Bt�r�7af1�
�tM�l��f�jAI��6�3�92Hw��DMWaT�I�ڵ���w���*���n)�n;Ʊ� ʲQ�s�#\M�������S��5<�G��u""=��S��Ie|�z�NX$�8[�j:S����Œ�#�/c=˂���£A}���V
���A��:BێԎk^?����=�!؝x7j��t�l�������՟(萚�ԛ��7D�`��ĸn�q$���`~/���A�C̀%u5����� c�����.�����`ZO�X�������VDT��9�����3��-җ{6��s&3L�|D2��E<l�1%]-�d���4+:�?���ӛ^��z$G�Rd���:X�7��A�{=�#��6M�(�R�>k�pW	��l3)f��X�o�i)PZ�G�s����s/�z{+�s��H�!�f�=7K]����5���0�G'����ձU�`.�4��e$�Ӽ�_��%��ʴr��|mɗ�i��Rt7M=�q�Z�ʀ�)N7/M�=��~����!��3
��:��z_,fxk�B����M�� Xv��8"�p}����3�4y��}�S�A��Tʩ
	�����)X����tH��7;�ֿu��T���j���qSh�2u�G}iQ�Pe�0��R������b�����]53���
'���:��i5:u�7�:U��$Y����h�x�%�R"s����Wv��Z8�8z��Nl�ȣ�r��R&v:���?�x�AZ�y+hD�=�F(@�|�^�p_�џ�o��A���T��"c{��x�n��t�.�)���h���𹌱ۛ�C���8��1e�s����6���F�VG���@�R�N�f�rq�#{#m������#�U�����B٩l;K��]��l��^80���$��C�[�[���A^�L�NJm���9���Gw``�I,��y@����9���ü�@A|�a��!���;�Tv���	uh�8`�w��+"�~��G��n�F�), �Lo�7E+a]�����gL!������+������ϼ�d����|����+��Q�I�ߑ˧;ӕj��=y��~'�#�Q����M�^p�U:���Ǯ�m�/8Z����ҏH���^����E�4�!E���A�ۓ�7_�����_��il[]�&��O���dЍ:A}�6/�7�,)/�M��w��f)�uIU8����i�N�gW�yc�^:�ڦ�������[j����a	���Jy�'�a�"�W�8M�����6���?�S��Nш��`���2�	eB���j�(���Զ9��oqiӪ|ܑ�~,�`�@�ٿ�t������������x^�+�/Ѓa�S5UO+i���8C`�=���zmMQ"�A����j��xHk��u��	����������7�a��?�(����
f(,k����,3%k�d߫d�XqO~̗��8���&�QB%7Aq�A�'C�,������=J%�6N@�zzR�ߟ�H.v�ʑF����v��lwq�C�0���=[#�!
 h�S�t�)�F�-��
!lv�%����㊞;��D����iǌ	�����}=���Fӄs�X��� �(������	U[䘽0a�Rڷ� �s.09�9��ϟ���H�a�y|B+�/.����ҁ� �-���QU���lɁICF#���c0��)v�+�x���ג(�c�ۺ�P��P�-��W��9�P�/2��*�2�ݯ�iy`��+��K�b��POY3G@�:B�@{ꂒԭ�q�@���"ߓ긙�L
R�����>i�ϟ#����gA��:C�{)�dݠy��ZF���u���U^�x�?���������F�#H��}�жrK��S�#�ߩ���X�=b�9�F�c�d��:�w����]�A��,�ݚ�k�ϙ'�I���Kξ�w U,�o��@ӝ��s��{�}[X�� ��-R۱�k}V*�+�ӕܳF��=�WX�ԩ"�ԥ���`�͆{����Ӣ�M�F��m�h�baU��^[�1P��7�1��&��1����9c�u��kdwr&uλ����(��3��Q3�U~G��sjϡ��Pq�$TLP�����8
��}]�mpfT��Kj�e緰c�Ay��G�m��.��K�O<��d�2�o!�uio����Xŵ�Ki=禬�c�<�<?4|<o��1�6ٞ�_T��B��`C1v���iF�kC��m���;��XYщ�<,�&"�O|0�������ɑN�x�~L���cZ�Z�8����,��'�֮�Aw�+�La�[��Wg���Uj����+��~�|e�������������4��Ł>��1��X�<ٰ���W!�����$ҹ��p�����2�<t^Lt�S<2!�nl�;�=S���y~O��H��.,�8�k}؞��c�(�^�4����/<$*o�Bv����<�A�����H��=�5eD����%{�ԡߌ�����m.5�C�9�HB8����A'�
������*\�$���ᐄB�{�1�3M8xog�.�L�N�h
��!���`0%/V��Y|iu/��>G��ߥ7��K�E�H��E�<���F��*`� ��M��h
�G�2��,�"�\y¸��h� G���C5�AN�$į�Ky�1�@9A��iIz+�{'��O}����3:9=�����x	c�:�{k`B�0�͈B�7���D>@h�!�v�<h�����p��'~���f��`�&�]I#б>�w�n㻜YF v�=�=�u@���V��I��=1���=gbS��Hd7578b��Aq�[���C��\p��)}Hyw�`�}���@;�,����:d�;P�*z�O���O}2���Պ:R|n�3�r�MT�G�����ԍ�=z�~/mB;g����Ӵ5�M��)�K�%W=�*2d��ؖ���z׶V�z&;����v
�s<r���-�����)彋>*��|b�}i��[z2����zz�;u�%.�;�� �0��i3[��M���s�F%(�׵@��@�mNSd�w���B����2�c,h�ۣ�n� �p�D�yO�O��g\"H�Q�u	Nu��Bi�*T�45�EVѯAQ�ZN2���9B�NP�k�nc1�⧈"#[	]���s��^��|�S��/<O�|ً)��yϴ^����ש��z5w�3d�{�h�+�T�'(λ�dӦ��u"�
a�I�뤿E�D����O�!֥~!H�q�4\|ÊhuB���G���m�r�Z�]���H�M���t )z��,@�N� xc����d�6��0�pXD7�1�:	�d��+]��D0��V�usv����}҅<|���	8�u��Uf���TY	�S�~i-�K��`��T3��8��tO4B�D��D�Q�<y�����!w \���yI,'�iĆ"Z����$et\3���D:���	-�I�I�� �1�����c���~���;�Z#��Q/ͥ�&��Q��g"�I���Q���8���Ŝ��<�;�����ΛQq���I�O;�Al�Y����q��RwV�o�_��ߠGiL�$T��}��rc���P�P��>�4UY�/P�PA��E4���Sf6��A�wD]�nnvlw;��T��U�]�W�G�o��(�� ��>*��O��c�s;ݑ.�B�����*m��-�m| yY�g�q���:�+�a��@������M��@wp,p����c'��1�{rm�\��,4�8c�l@R���}�F&��8�;l�=�b�ت�[�!.n���G3:y��;DXm��#�X�N��*��(zmt��m�=5ʧ_$�oYC-��(P������¯E����y�h���ywwp;���g]���n}ԡ�N��ҕ	w��-�W�R�t��\ӸlӉ&�rl�2d�d�)��'L���2�����AWc>e��qnj�`*�ކ����>$5u�4^i/�b(W�o��5�	��Q�-��R��C�O<�Y��3�w��M� H����儗\Q�7���K^��m��CR�'�L'�-=%����w�!H����$>�2��+�T��=�����>A'��m�j��S�m�6�T[��vkB�01��d~F/�x��n�E;Y41����1�����˾\q�У?\�+���b�=V�9��=��[�r��L�k����~�����ܺ��]��NlKn
0M���{�&Y�Iڷ1�p����`����أ��c���.�����iͳ&����Ǚ5��W+���:=��=��0���|����!=5ʑ��!f6�)�1��\�u ʝS5�����+W�� \R�G��(L�82NzB0C��+4y=�E帚8!���S�+.�?}O\Q�F���G�W?�����А���l<�TUR��eIGD2��MCϤiN��n�fj�_��%�3�N��g=�g;/��(Df�>�rj���QP[>3�<�l4x=���8�n�V��Վ�݃~,�x���Q ��V�<*�-c`�g������Q�'�Y�2�����\",ݱwY�&��s����gǺ��d��B���`_<h�<-�q�ũ��-5�-���@5��T��c>�H�S���`J	�`��G����+�'�Ъr���2�!o�y���wo�g��v��$�kN�ៈw��1Èݪ�3��w����`i!Y%G1�	��S�r	���7�6�t�ȍz��Z���I�a4E)�y��[�^�X%�7X����9Y�<�<X��`IL�N�5��=�#ߠ���u�c\j}7��`f+Cg�Co�}�?>��>ҟ��־�5�m�<��G��{�N����Ο���Ȫ���L��<B�-���׬��i�|��%A�S]�dȨ��s�̉�},qÊ>��!��/�*}��?�b
�H~�!k ��ʻ�a?B��g�sY�Zo��zz�����F�����B����Ր{Ed�JӅ�נ	S2����*}��<��3�d���ʧ���������џ�~��ϡ��Y�`{\_���`����J��po����@]��<��M������Q�<.��%��pЀT����i��G�����,��\�VG� >#�4풿D`���F�1{p�E9���
`��Q�]=y��Jl��U�;z�D�IXP�Z�H���8����d��B��h\W'n�0VB���a|n���Dȝ�:�
�϶���yl��\�b'�s7��>��q�iI(%�c}�}������~��I�.�p��*͞�P����BچtRս��{Y���s]�����n��+)�EH)�T��N�|ʳ�
C��ˍ�jT�n*-����T�R]鸭�F�FE�
�����.G�U�OJ{eŬ�s�=O?���{����7�d�ԽM���[3�Q!*'|ׅ����"ܙ8D٫s����ϕ��j�TaVd�E�2JKݴ!�[G������������q����a��v�PsQ�d��֍|2�uN�k'</TTj��6��(m�4n��C��=�9�p��JV��Cm���<�O3j���-t��e}���F~���Q��]F�(�bt��?�\��`��"��2��c����A����Y��/��zx<d&Ep��lT5U��*}����$I^2�K�0(�vi���s���.]�l��0ֻ�jK�Ox�v1���U����ց7�u�����Ò��B��8�)��Ʌ5��ޑCj��9hZO�P�\/�#�Y�i̧5Gπؼ_�_
�=��k��߷� �:���/>B:g��"E��k��d�ھ�^�J�n#R�I��<+ba�8�����|"O����t	�`�Cֽd�:���\�`�k��wq,�<�+H1�Exfe?���99������9�#{j7���*�bT����*�Y�%��Dc��8ȷ������Q�B�����l2VM���t0hǠ�A~3=+����Sq�B��B��ڥ(�&�p�:f����J7s��V�f��0�ݱ�;;9'�'�}�:5��^��W����f��(�� PG~����V,s2�cb���2������
�p�z}]^�l�q�:�jTN��h�R�{fCM� ����N3��"0�<aӑ�{������W���W�1�_$�WB:J=�	��=�K�kO6��&�u)�^���|K�Nq���X�#R�H*��i���7��e�Sa�r��~J>����4���d��#~]~�-�(�l��M���}���K��#������=Y��P���\n��'7���/z�t�g���ϩ��xɯo-�ȯ�W�С�2��%�7V���\����+~L�kȾ8���p}N��\X��_���'~��ǡ�(0���l�	��|��k`�2��8Z�|}��P��W_g�*��3���� ?LX���w��U
�k���z;'�Wt��4[����r'�DӶ2�?���d�������#=s��~�}�w��M� ݭ���9�R:RF��O�Km���>�����*����S��^���� ����S�a�0R�f��R�C|�U������*cʱvP�*�P$�HS��1�%�qL�����3�~� �q\"��o������3��}쳟��S�;�=��i�7�YB`X�|O���(}̰D�qS��+5:����c�E���l&�#*jA�HUħtHM�K=9�T�}~�w��UA6\#��{����3�~ʚB�Wn��8�W,5m�ӌx٦��+�֝��)s���x�HקVT�ʍZ�(���UP�����L�8MP�1�lA����4�։i*�A���8�8��,��z��a��Y�wԛ��Z��0(PF�]@w"��~"a��8nx+�ǁ���6S'�+�#֥��������"9,_�S}[��u���.�Ox])����v7�/���ꉧM���,ܡX�KP�܇�N��>��R���-�Ś�dW����[i�hr�gZ3�
|}(AX��э�f�r̳E��\�w�撚Q��CZ�ZW��5-@pp�� 幚���O�� -w���
�-0��#�y3�{������4��ؙ�zG�k�
�6�������k=:=x]���)ʝ(G�n4���BI�!���'". ϢN@+����1@;��"�Jt�>��d2���F�v:��F/ �˽�A�rz y���mq��_���1�c���+�����$����0�>�ޗI3/b��@t,�c��E ��}��o���-�Ҭ=��dS�Y���uc��&��[��='�	d��z�H��~Gyͯ�]p��g��D��� �矱�@��X�#_�Oh�Ǵ^��g>M?��ѷ��k�$���O�(�c�4bP
�_�z�����3�3��t��)=�`E/{pJ�r��HC�r�Fڐ�>��3�
����Ӕa�Y��\G��-�`��u�4-�2r�a�~�X�[�,�k��`�ש�1��)��<���s���/��?���g?K��3���<^��N��P7����c�F���v����}�Q�������q6���e���7��{	P��=m�Wo���<�)TaE�L�-��<�����tة�M��Ξ��T��/;�a����a7�`�oV6).j�R8�xɃ�;\�q�c/C�i�V�L��(�-�a�]�������`��G�Xva6=�f���'D����	l#@~�`5�*_{�ߣ��_���͟��|�k�f���qD�3=;N�Ax�~�_�,��3���~z��t�I߈to�>�Qa�5J5�p���h(G˭S0E�锘��U�i�_��r�n���Q��y/3����qc|3v�մtTYjg����k h�W���7R ;���$!*�9�,�7��i���:��J/�8�Ĉ�Bi�*�]C��'�6�Ge�[�"33��^P�|8�P�U��8�=g���k5H�F7��r%�T:����h�W�	Nh���
���l�z�Un�Aw�(��|
�U�+�(�r���/���m�4|�i�Iá�M��0�a7�vK���`�:~�f��a�6����C�
�u&1�����O���E���y����gx2��p������l
l�?�dGϛL��8^e��/U~�{�����ɳ����.��w�X��8�,��IԾC�&X��b����S[%���5�UYŊU:���][�ZMK�c�?h{,�q�vB�*7s�Mv8D�����A`�W�������K��{����*���a�N��#���*B -�UJXDP�(�]|lP��Jz�a_��r�^����-.�OM⾫�~8�7�v�q��+,�}��mi�<����\����!^�~T^�����ӫ/08(w�V��q�N���bѪ�����a��F�\#���Ϳ�t~�����,��7����@P8�"d�D.�2i:�b����@��8}d#U�;M�o�tJ�w���C9��d���lʥ��a����S:�U,a��)�I�Iv��=q)o�mOwd9 ȩ!$*C�J�� �f���u��	�n��-<��v�f������q�6�S7N�����+k�9]6"���G����R�)�\ �70/P��y��5禲?������j�N�4��Cj����@9V}�w�O�C�n\�g�U��Y�7��q}���:~&h�@8�n@��Kฃ� Đ�l�<��	�LC�F�2
%1_D��w���u�b� D��c鵧G�V��iؐ�0���"}��G��������?K/Y�jѡ^�C��g��*�1�^��ӟ��7�{?�����Y
)�1�6Ę�z2l�j(��BTˑ^!�UO��O�x�����>U�^N��:m�9D4_-�%��¯sZ��/����Q&A:�,��W��4֓<X H}��B4�<߫@C�6��h,gg�-��z����A�G�|����E��Y�	cX�h�-�a���z�@J�
��Wh�,�P!;R��`����P_!X�qJ��&��������H��.�����+F֯�{�+g��`�N��m���rS8�6��E������D�����b�ֹ-�x��(vdL�ƾ�`��-9I!}=�Tw'DQآ��w�pێ��͛]��4�r�W����f3��AZR ��{���T�u�w�vz��I ��ٚ��$�>��[�Ȅ�o!�(dpi��V�1�`U��������3*�F(��(� �IR0/	�5�q9� �������Jm���8���yT���ݐ��~��x�����)�	t4��7��`)�2*�u�e�h�r��l�y��T�#�j�7Tڬ�b[Pz�8E��6�ȿS2k'�&��ʿ�8��4´0�hYڥ�7�0��]����bN��K�6.a�����P��!�Ar�M�zKy�q[[({�Q3�L��ԟr-ϖ����2b(��UH�~4ܻG��k����_��z��Sx��i�,Z|�\:����@��5�����w�k�{?�	zax���^�ϳf��&�!���U(���h�!D�o�$d_�*�+JF���G0�|UIv���F:,$��3F�Eu��ʖ|K����S(gX���u$8ɃX�;�/TJ���Uo4��4��|%tc����L=�5�����q�����FI+�!p��A�>�`�G��	����eh�Ӿ�[�f���^�w<�sb�7�3j	T��Qumn�>
�N�4Q'\R���n�y���] ǡaf��mlƃ�܎ɝ��%�K��gL���0a	�r�LJ�Q/�o�t��v�J�%�I�/��Gt��ǫ$Hl��;����C�mo�?��� :�/��5YV�Xp����?D��G>F��#�^�<�@B>Yc���\����>T.Vݡ�6I��f�� V�2���+��h͘�	qE�����+Hw�<�Ic|S+)(&�/�6u�Q9>���"��C"�81�RR�9ZA��2'J��ϡ8d4���j�+7�@�;B=���B��]�;���~n 4�ݗd��׋T���p�����bCL�����|z$/��E�gZ�������<�B&˘�e���ޢ�-gbL|>rl�a��}�%ia:�����$�.�{wl�Y��.�-c;;/��U#F��y�g��8QQO��.�s߶��cS�j�j(��@.�e���zL7��ܖ �{��RY͈{��M$sS1�evt���	m��Ocr����:�o5GK���_��)\{0Q������8e��Yl�`s�F���:\�*/�:��a�wa&,41�8�V��
�0@Z��W����e-� �:z��� 1������� 1��_��1���Xq���ˆ^p���N��L(� \Kmv�;"+�L�>p>������AQ'��P�!�9D�d�禓c�d�Y�}��$���	2�=�'�{���3���ߒ�N;����/�_����Iؽ���8��G�?Q�x��9� d�[�<M]��������@%�<���x����|� ����N!�_�T2$��ac9��< �@�/l����������^���fY�{��a�'��J*���O��E�_ۻ����g�i�'��q6��K��<u�'a�����oB:.�Ҝ(Q}8"�I����II[)�	8p��#���jU��딃?}�ݕ��a7��Q�>a�u�! E� �L(/�<uA�':���R޶^#�!j>�7^ѥsP�p�@d!s~�WB�H�}��V�v����q*��5��w�-���,�E/���rO��Ss��ϒkM�,�k�o}@(������=8v�L�@�i��R�+ �!=%�����`UR�|đ,>�)�?X(��gf�DB��%�����ģ���&��ɱA�Mv�bV�"
��`�X���
B�C9�+)�)�,�|
�sO���'��׿����Kk9Ē̩�Ij��˾(�_yכ�W>�Qz>�D����t�[�q�
|�F��P�eY�Y���L��̌��2<��0��H~�2z�XPNFnl=ʸ�
Ӭ8U�T� '~�8��^��wք��(׏ P�c�m��� Ք좜� �����a�t�
��T008`.�[�~����<~ߣ�/z�@���u����}	�No��Ȯ�O�ȅ��ς�p|�|+h	�e����0�m1��x!�z�����ą�zd����:��4�J#�l��Eq�+����<�{\�v	��~q!~t��k5��&��%�r�h�������\_�j�bNVe��/hHP�l�� \���y��|�ϩz���W6e�o$ ���U�\����+�'�l���])�µ� R>@>��-uS�;1���1��2OFO�����υo@�"G�Sz��5�k,�ựu��35���eg��I�!�S���3��2�b�m[Q'q]�����=�DS}=6}e_�50�E} #������S��8�wTi�MN�Ղ�*h�W���\��c���V�S�2�p?�3��C��(:�`�
�>2R��U��H6v���
��zѵ�������N]�;m/��k��8M�L �c��aFF��lFs���{�����г�y� 6��G�3<����fI������>Q�۴-�Ŕ%���s�<�7�/}��w~�G�{��?OO�Sm0�C�Y;���'U���_F�k�H���qH�����㐯L�h)��7�t������W9�Cy4��L��yP�BC��KRY�5���j�⬗���_�M葝@��T_���c�>D�,�F���#}eӈDvatć,z��'p �0v����<����A�;�����1(����y�B�Y0�_�	#:���㪜��H���10��U6@447���w��+;��F+���A^��ڇfR^�xL@�����1��Fu�g��	��]���Ҡ�ċb���,�B�*�&c�+�u�Z�1����S�~����s?G�=�L�Y��DT.�.���6N�8�ӷ|�[������iu?���a����/	*�p�	c��l`�0h?lOJ�e����I��+cI$'M]\<H5*|h�Ş��%� ���HE{��V�����&G�RG����@>P��z�d��ԝW��PL格� ��b#4�����A8Bڮ˱v9����'��p��[�$��v��i�VfX��šǐע^��P�?��z[�m�VR�P���i��\h�v�D9���4��q��o+�8\w[A�=q?������m�}����<�N����� ��8�BԜV�H?q�#��[���ve��aL�]ׂ'FT� _Rpk͂Y�m8��%8 D�rS%��~�h4#�kx�5���
v�IX3��c�N7z�{�����Ǌ۶�~�)�����ql��d� ��	6Ƭ���#�d�a'|�#hąZH����UZgj>��ͻ�!�` C6#1�����D����<y���
�|�ю;XK�����h�X��U�4ޭ�^P�����ϧ���u��\j�ޅ�{�C6�.(���*��vA��:��t��W2�([�:�'��p��m���[~#�|o��Á�]�q�v�9tL�z���mr6��h9d��8Z���!_����]y�EO�����O���׾�u��P�t��9�3c��)�ԃ�����>�[���>Kt������k�d�|ƃ����<��������G�U�f�<��u;.E�"�P��z� ��ߑf+yB͟���r��z�6�i�3�>"�8��%�J(�L���<�m"��Y�Cׇ��I��o�Yj��LXrb��!y>ȶ��9��:���.v��LF���;ʯiܖBwx����+T��N�xu�߄�&s�	nD
>Y�N*�m�1:J��Y�e>\f{2�N� ��1�:	����̓�ߧ���?�U�7~��j���� I��:���K�Z�_�����g�6I����� GW���dX�(l��
O
��;6�Z�.��@���*QK�!�1a0�\U9���/ �3��x7��R�Hap���OY4��Y��(@�JHrl�ļ�2
��f��5@Q#���oPE��U�F��m5�*�UJ�$W{GQ�Q�7��w ](G��

�0��ޫ�X驈�Q.�'��Xӭ���5V5k�>.�N��D�<m�Y+�����Б���UQ�9
���r��\��fqwi9��]��~������ڙ�=L�5c{ �B�����5���u�m-z��;�|��S0E��v�|~ĘTc��zt#{o�;u���lf��=��~#�N���2Lzy&��/���w�9�E+�x�YxM`t��nk��M��h	Ak�A��� cT�2q��Q>�zT�e��4ϑ�ڳU�>�o)�@��B�[��Uc�j�c�\hz���szz����m��3'ۀq��Vg��$2�[e�!P�� ���|�k��u\��KP�9�Ґ"��$�����V��O�O@��GiozQP�:�����I�3=�}jhPG�-uCZ3\�l��$ �������s�;�9�wD��^�0�ݙϸrsz��3�A]��N�oï�6�i�, m�4ѯ��EO}R��XG��%�;��h���G��"3�d
����Lp͞�1����9Z�J�ӷ|z�l��I8�m<:����k�;?���e�����'�'�hs$�F?O����}��_x�����g?Eg�X�|�}����tjG�L>�ć�	����9��]�ט��`�V�]*�X'g�J弌Z���o�9��m���o�A���� ��̈́�֗�<w?B�&�䦣Mӎ:���5 PJOAW9�� � /���ْ�o=ϩ�mZ��G���"O;�����z�1� ����� 7sW�l����{TV����Ey�K�����H��c�w+Hb��>����He�E R/�I������������i>Q�ÿ�;�������������"2i�o�W����_�:��w������"�����R��8��Rd�°Y���7��A��C6�~壞��U�\�V�SY�9���h�PۤwbeF�`�CJ�-,`��b9]dp�Y��*e;���0���5�a�
4xU�0������T侎l��
,��ЫR
�A�[U`}Q���=9��{%�����o���w����";�z��mY"�uG�ci��S��x}CD�q��`)>u6"A�����o�tϳHS��퐦
ꖴ�>_tl��p,�M��p9����؆�~MA��qd�2�ϫt��
׋��Ǔ =C��)S=�t�s%��I[F����}!`�ש:��8Y�AH<AS-v�a炙��,�3OT����&RD�!���Zm[1�rB�#��٘�k 3��2P�Y��%�X���F?��['i"�p��F�\o��� H�E�Q�ͲZ	I]Z1�b��?�;,���U�Vҫ��s��[���AA�H��&_�����>s�Ɇ���.�tP^�J��ɡ�tDppS\x�;ٔ��A��P�S�Ea�ה#���O��*�]��t����I��o�Js28���c�r=t��}:u^��1)�{h�Y�:���h�gp��G�m�S���^*U��m�{@�,���Y�/�L"�֤�w�҅I��{2:�`���j��^��tcx�	_��|1}*�KW�Ǹ��pB������{��v��o�:
�cil}Nf�g�x�rw�s�_���齿�����|f�;�`T#)'p$�b%t)�M���Ѝ��wP���S��� J�����ށ�F*^�@�������|0�UqM���Pi��= �R�r�L�ٴڃ��JrI���5��������OQ.���fQi��r
��`���ˆ������P���⼱g�Q����W�M�a�dm�����q,��,��A��L�}IUc-+r� ��� �<_�<�{�M�A8`�:b82��)
$�i��fҔ�P�8�+�7�<)�[Qe�Y;A):�����F8��~���?�������Ja�D�#��^���T�b���pB�����������6so�/#T��}��E,�����	C���0���@~Ń�X�C��v�jA' �z�j��%�|PF�(a������`^�Ȍ���E��t��;��H�M�D�q��2�lm��9�ӢC���p�Q��_5��]��9���;�o��nq��L�D�膩t�4�Ӝ�c%h�E�{G��쐴u���9��Q�����EW�u"G'�dF�l��Қv�����-M�Ϻ��� w7���.~��˅��ŝfp����e�Z".��3��O���b�:$�92���Qhd�P�PE@I�zpH�d]��<Ns'��*�v����o��߄"���4Eq�FuęwY�T�Ǳ�ZтKt�y��Lz�ڒ_� }�����k�Uk_B1șC�R�Q�:�O���7f}o�'8�|��7y�Fz�fZ���S���{��g��ϟ�����h�7�i\�ɸ*�;�儆�.7���Dk����ب�6� <�ie���
�tRx��@�C���>��.W���P�h4:'������7��iIYP�˸S�@��2��mxޘ uNF�/;2�=����l�:*�o�ȸ�-������8�+O�y�gN'���%��w ��;��-�ݧ͍{��0�v!��L�(x}&�ry�b��{��e@�C�5,�nt��?M��ͳ�_`�5΋�3`�7^��=�:F�9���n��{���'����;��:7��fE?|���?��7��^���L��Š�++W� ��H_��/���O��>��|?=��E,D.�U�^�"8W�9�!�S�G�k��:���:T_�`�/A�.���� m�GP�&7&�9{,+�1�+�c�I�ބ�!S�q��MX�y�8`=�i��\��,J���;�}��`aL�B/z���y�v,�w�=�Yd�w#K��!���ӱc �a̝�:���
qbQ�SO��u��<�j\�J��-�yh�j��X��3��j��ؓ::F(V_JA���o�K0@Ta��m��xi<	�:�0�ͪ���H�G����/���<�N�R|���e�u����������{���?��c��b+��(�G~&�j�a��ź��[,W���I�B������Ȏ�FxS��#n��E��6�'�
$5�$����Y/Q�q���)&B�ez��Y�7���2��-�/���+/�s�2{(��&�8��E%�JV���
�P��@@��2�'�WYD��j]�ZT!����j�D'����%�R��m�C���T�PR�"i	���i-��44��4C0\;���4�-�U2�I�v.w������3�	����wq�P�&�Ý|Z�c|��yu(/�_�x��l��<9���Ǎ\V�����,8��mt����/u����W~[����Y�����%9XV�� bh�U������:�G#v҉,���'�O�N0Φ�XA�I�y'�JM�� ��)c,������|M����}z�k~����f��7���/����>��3�s������֛v�X���q#�e�����D7:�'��2X������#��"���wN�ZVzh�n��;��]h���t9�;�)�1�_�Fw��S\G���CAy·�g��YQ��k��Ө�e���T������DE�����F��ͻ���EKd������.�{��p?�N7��ܸO�p��u��|´��\��8x��!��Q5�eq�+�M/�n�6�rñ�
�/1�J�k	Z6����?��\���z'#��ڃ��gB���A�y�(�N��C>����	���I������������u��2�ڤ�r�ţ���w��������}�����d�t�w��p�Sq-�$�z"G�HSa��J9�3�at��0���G*����PH�=B;Qi�llY���kVЙ*8�HB$xr�<(~#AA�'%���s�9x�ҿm>'��Op��t�K����4l��@ău5�wNfԱ�����ǹ��.�Դ�؃� ��������{�P=7~�o6����GD����i��U94��^��9�<̂�Ʌ� ���H)=Gh�3�6�xz����I��~�������z��Wn�7�g�ǿ�k����!����4�夎�UU�Ge�\E��av���f3Jf<�oe��'
;Uf�=�'��7b ��5��&�j���"c2c�;-C�/ׯ<���O·��
�V�5FF�6�DS��8���8�cw��v�w����$s �~�bOD`��+l��`��S0M�N�8iJ[V�� �e<9 |�]nB�R��æ3����F�Jf.-��#��%^�7�j�}�q�i$F����O�3���?�߮�O��%i8�d��yli>�������W�Ig�i�޼h����0������@�����M�f�D �K��"H��±�&��1u�NuPYz\ڬkU!�:�S��fʨ�'Eֆ]܀oǺ����F������S�.c>3����,��Qƀe��Yv��PԨ'm$�J�F9�9ه���qN�����4_��G��-��oz��?8�a]?�I_���o}}×����?�A����zu?�u٨9T��.!�an��A~���D?�s�^[���G��6��(�A�\�mS�VY^C؃��v��n�:�2pdY �l��i"��7:z�~M�u�+�C�R�-�m�D"b��}�~���袃4�h��:Ve��ȿ���e�=�"��~q��>�wtt��pߢ3L/�u&�I��z���=��P�Àl��y���r�1`/���1�gK]x��+�]�Z���Y��:;���f�rzw��0���(UU'�כ�7i����'����w���З�����Y;�D8���w�7ӿ�w�A��X�P���6���LވJ�;�u5�9	GV}0Q�����K�_��V�){G�0��~~8n�G�F[.C���X��.��l�	YU��&H��l+:�f!�D~����y՛��6��1��q��9���yx} ��b4�4�e5W��;�嶂#��pb�ƛ���|�k�&�qѶ�&n�w�b��|�P*"h$ʎ�a=�P90����x����*�g7y��?�1���z+�⩧)�+ب޳��D���������;��C�=���P�28�"0����	��d�BF��2C˴U�Q�R;M|F�G.݃��2J!��������`�Fh�f:����#;�{��3G�h*�A60�ڕ���A��񶁎y$v��X_�S��(��7��H����vJ��J�;(V���R2��p�΢ǵm�["�<B�i�zܚ��^d�Cv0m�N_�D~�^]��td9�4�k��~!�Kp����m/���^�B�~�Oƌ�5lw�5�2E�Ei��$�$�ʸX�����D:Y�l��|4Wd�����p���o]�.��>�gN7�d��؈�v�e6�/������ʕ"Ļ&��t�?&K;)�/+F�Ff�A� ���w���DEv�ҟ��z$c���p��ϯ)>:��6����_B��u_E��u_I��_E��	��tM�c��s�@�Dk��	}�[�B�3}�?�C��Ͻ@�!��Z��|4����I�=)��P��-�:�җ8�7��:Ss�Su�* y��Oͽ�p�[D��2k�Y5t�Y[�1����e^GV��n��id��#�љ.�Xi�-OZ���h�E�C��S��<�l�e'�XL�Z�u� '�l��1?�2'�S�wnV��1���}�n�$����b�)̔�4j�����2�3��flC��7BY
�����.�"8z��#
K[�}�����%.Y���f���[�K� �T
s>V�+���O~���?�Q�����{�g���}0���3�������ӷ}�[�o��/�9=���堇��������mo0�M1/��/���O���Vp�|�E@�7P�3A�saP�B|�����A��v�nO�P�!Vz�w��y�)�� Y�ϝT�Տ�����>�������C9"�˦�r(~��n4�&���RӷP��8�i9�����B4�����dgw �x'�;�&�-�[�3�mq[��R���t��B��V{ؐ0�V��4�+��~E#�VF�N�������R���{�O�6��{����	Z�4�|D�L�6��ZS8{����7�7����ӿ�iZ߿���T�2��i0�<ƃ
ю��U�]��Tw��dƮ����i��`GPqn ��1�|�
>�-�g�W�� ��҂�a����69��ʬ���CGF/��Fa�#��� �@Jk�r��H�}�Q��𴗫k���ϾV�vţ�^׸f�=Q�.l��#g� `ED�s��������ݎ�)Y��W�B���k�M��ra�\��P���Is���Á�ҥ~\.�������a�h����^Z�i�4Q��utqu�w^H�������Ӄ�<9�Sd��ީ-��a�w,�K�wpx^ӫk:��=�x��s7���{-X؞0m6A���`�.)���m�H�@�5$eCӡe���r�C�b,3�,�L�T%�J[�`�)`*?�#��j�M'k��(��� ���#z�����u�������m���|1�h8��ʟ�K ]j({�Y竻��xMt�����/�?�����������@��A�
�x�]}I�.ˬZ��6������&{����xd��N���7:TP����Z~�`��q�u#�QEM����t�k�å��jRP?���|�v
��]�֭�l<�w����	�I�G6AeB-nډ`���3�d7�Τ|NmZ�#,L���}9�S��m�nҺ�`��{��9�g���?��:���7�s}��*���O�f}B�1'(k��ć���K_�e�e�._}:�è���K��&B�}-��u�w�&k������c���NOO)�?�����~�_�w��?H��o(�G��̣�s:9#��?��� ��s�|xG�1���"�V�DH�
�B�G���*�e�:��ex�O�U��m�e{�7�=��u��4Y,���&L�`�ϲ���N�7��W ��va�C�B�}0:6>Ȥ��x�8#k��݂�F�Ѣ���f�A��݉5�$�ǧC-��Ҹ��0�'�G�ԡt�iA��&�p��'o�2|Hɾ�x�wݚ�]^V����?{okkr�U}���޼�!��*�I���47IQ$K����a'Hl'?�Ȃ @~%�0�'A~1l��A�8q"�ڠ͂�h%ER$%.�}�ې��w��:������s�=w�[3�s�ު��k鮯zx�&�p�1\c�	gR¢��FUQz�Z����{|�)4$�ŷ9qq���g�F���6��[��YH�=�Q�]avWǰ>]��k�G����7�^��g����琤||���>�7௿����O�<�o��W�w1w,�;Ho��y�XuR�_bc,)],�ܙ��,ܥ F�'L���P�WKy��WBb�z�pDt.��B_=$FeV^�������U��-HŁ@�u���Kb>�nH�4�s;B��Q��d=T���".x���]*^N����n�p_&z	h���;u,�A5�iUF�*��J�ĉ�!k�h���6��T��
�e9�}��&Z�%���v�p�Lk���o*�p��Z�.(נ��i;���a)�g�W"o�F��L���⹹5\�	L�$�C�_��YZ��� hϭŸ4�����}͝����zI���=�r�_���.�Bc1�9�w`D2V�(�Iy4�[�m���t�+���-E}9�
�7=#~�(}�/%~_�y��a}�>��cxӋ�?��W�;_�x�K^O�u�~c�N'9���P���&�O��佁p�I~�����?� <�.xb��ʃ�	��&q0�Z���|����Oe~�Yu�*�L�����t uZ�-+�%�5LC-��hF7H�"[#��q{n�T(�:�q�"�`Ʈ�i�:͊���>����Ȍ x�Xѹ+����J�xy�:E�-��Mӥw���l/�M����0�=	���WU�Q'�}�[��`�r/����}��i	��]�<���9w��F��	B�&7vV'�r�{���8�L%z�Z��b,��jL��S�	���c8Y�1F��W��+�'��?����O�7 {r�&X�F���fS�e�z��/�O�����i�u�|��x�B��t#����U��!�|P����C�e۾,�>2?��L�̛�CU�o�� �����>o������-Т�q�o��㝙X*=�zN>7+|�O�(�Jqi�G�2۔��/rݏ���+�,{:��)�_�-����J&Ho�_vn_h�vR�T�9p\~R f�'�	�K�T4����-��Yޟ�)Wa���l���5�nkB�\5��)9,H�8(�acPP�j�~]�c���������/��������!.n���� D�tO[�H�.��yρW|w��/�-bC�F��GN:0�x'��M���_}��E�kбWz|ة��\+r�Izf�9{���4Z�c@ºV�wbCCW��s��|�����-��`4}�j��X��k���B��9&�=�o�^l�UO��U��8���q��%i��!Կ��/(T��'p-�Z�+X��D)�A���R6�hɺ�vj�pX��[X>�i���Jkg۴}�7��?8<~�p�{�N���� �~�d��{Eu���T&���()�0�"g/�������*���n��Q�z��?��E����]� �5ɻ��SZ��j�ꭌvm5nu�V��@?�잍"�!g�>?�}���C����lX�ic�u��yz�I�q�>�졇��oz#����?��#ތ�6���F;�wk�.w���+�JC'��C8�1<���ptc�n_	�QCɑ �.�Y�,��!���!ȹ��B{�h��PҊ��f|�O�he��1�.��.zS���0 �� �5W�9�����0��-�Nm[ߩҾ�������'�,�#�~I�)b��D�e;�_��K�wN�F;[���.�m1�߶�,��>�m���N*���	��u9���	��Q~����a����߹�L{�K�5;*c��V�d]on�²�m��z�O�D:�\�*�,�.����hW���m��g=~��_y߇��{��R��|�B�u�}F��p����xZLZ�9�G�a��3G��$ۋ�F�~$$�̏�K���K˱�C4̣Y��S�E�
e:�y�x���2f�Q��Hg0�]��&|tP���+l�([A�)��Ԋ�t;�vd	Ҟ�[�h�k����g�p:iupo7�$�P��M�Fd�*�g!���Qv�ao8�	�=O��nS�XA�h�x�(�M��1zQ�
)�W�wѡc���o���/�����_}���kMBv��7l��(/CG���5��J����
B��u�t�\ƫ\{�P�J8��C(p�j:j�,7�x�f����H�P@kN8� �h'Z�4Շv��\4� �#�Q:J�����S���J�$�Yk4�qG�ı%�ګ���@�mt�D���|>X���Ji�\��e��1A���	ym�7�r���)C��)U�Q\��IwH����1�N��+7����:=z�r��ʶ3�״�����W��&����͋��g	��4�ZJO�2��`��S .�[����h/낝c�Io�b�����N`�!�қE��9�^,"�5�$.�=G����`���#����qu�(��^�|٣3pȕ����m��~y�k�'П�����GVG�C�z��;�o�����v��kO�`���'���ܧ7�"_���"^i���!fEF������:������!+C3�g;��Q��Ǭ
��N�49zb4 m6+'7�FK�2�kDy�;����VMBY�*�� �����5s�g�C�]���~'�ӪR:$�7>A9YX�R\X�'��.ב:��PO*�f��G�;R�Ǩ
������o������fR���3�4�.���ྕ��m)m�FKmA��=�@���'��{a�>pM��$߼���-�g��8�I�����K}��W��i��ֳG��0�O��3���X�%����U�ѵW��U�k�w|?����ŗ�^��go�^�e�`мcT���nt�Jzx��1���Q�B$��.���>S��yL��n^T���s类����&�S��n��6k;��`� q���k�<���- �,�}�N�R�r�O��6�=���K~��4����d������;�<ċE�]@:�@�����؁e<˳�?. ��/����֚\���s���g0�ST������lRk��b�������6�58ql�����O;���?o��W�K~�p��&�D��C��窇�.�/}�cpwu��Z��1��>�JR�-�+��$�.��hmn>X��?��ׅ4����ܠl��y\�Yԣ�b�T$���
^s�F�C�^y�IDi~�D�j��|�6�%8��."O���>�����q�c� w���`ט*%lqi���hM�v$�WoR@�C�b�J�� ִC�*m��Ik���W�x���vF�\uNiA%�&hU�mಘ�3�8�LP�=}fl|a?ʾϿԡ�G��.jp�=<E� �:�U��5�,ˌ�������W$e�4aH7/hu�8��W�	�'�Zp��z%c��N7�"'� .5�ř#�cA�lP���QH���l��۟�D���6���E/�}��ox��yφW�m@�&u��1\������m��M8���7��Ͷ䈭)����~��;<���G�r�P�f3�ԡ&6����6+�ɥX�8��xh�V ڧ-�|�Z$T@;7p�d�폷�"����������e����Z#��y~��W�p@��P�=P)�mm3����6ԊM��g#���%���b�*�!?������
)7�[X��=��}6s�ԶvG�_Kh;U�c�혴����e�3?8���_%5���5�g5p�aY�U�Vm�Y��í���`��� !H�(�dG�PP0�1c�Y�mt��Yw����ϟx��������3x`x�v�����p��t�xs��o޹���>p+a���z�_<���Xl�L�ϖr_���5$5ɕ]�=oއ��r��23��./mR�}�S�K:uH��,i��U%"_e��e?B�6PW��kA��>X�!�k�C;M|���/�.%�b��bn;��A��2r�9��w� �A9�M�|X��+�2Y]�����o���]e��ɥ60��VK� �xy鹴NkkW����T�p[�QVGGp�Q�F'�����/�
����o�j�Hv�EbE��Qz��w>�~x�~No< �M�x�mv��5��$/P�Iʔ.H�GSc��Sy$U�s��U^�����K�\����6��$d�*��1R�P���1|972MIq�C�Ca�HyUd�e�H���S��wp��p�@��rO����rW$\YX*�mR���x�	�a`D��e@�OJs��V��i��g[A~���y��&�8T��NS�n�f*���rέ�I�ͫϹku�_s��ai;K뜃K�c2�����&~9H�u�]`���P�:]\�o0ߝE�6[R�.�.04����}ȹC��mڵ���Uwnm�K�6jr��r�IW,�4����I,����U>t��O��α���h�7+w�����6�V�ADr�裻|Hw� �Q}�I���]Xݿ/}�Ax���~�o�w������
pS֧)r"��>g��'��6�$eS\�1�F���<Sau���~�#���}����Ֆq�1���񡲁\�oh]���8��(s)m>�/��k\�V�Y�K��l;}��,x���Up�Ezq���s�D���Z��&��h��O;Jv� �rp)R���r����G�Wʡf'��r�m*���{h'�W�	o�iM�}������h��ӬC�ϋ�v�I`fZ8���1i�Yr����~��;f!I._�n���^l�Pd�Mr��1�U4�R%/4�����@�ɳ��c��|G��e�TA�QN�}�AnSno,\ŋ�o�ٛ�'�~㓟�_��ÿ���d�~��0���?E�"n܀���_��|�Q�n�Q��M��6J���F�K�cLj�c3d�)�8ϫ�"u�n(cP"o�������� ������ӻرܰ(t��AM=��GT�)A:99E*�6Zic�#���~��j���<�3��W�XY��&Ku�Q��ߙ}<�*c�I�*o:#��y�����c9�����s����q]'�T�pB޴k)�q��8�[>��7=O(�JI-x�#E<b�:8
�&���
������7�O��pt�J!wO7y��xw[8>��|�Q��_�M��0Aot����v���2&��!�B<.Y�Kg�5��6�����8�E���:%�k�P9[�e�	+����I�9`zMʅ�m�<��l��ҥ�:�U6�4������*��^��g��.2�SЬ,
u�̗�9e�2���d�|�YB�W�H�	>���}K���fqy�|V9�}���y�4p~�rܷ�Aw�Y��Y��l�w���4��~0M�)=p��v�_�MP!÷�nmd�J<���z|S#H��*���x��[w�Cb_k��[�����Z��r��������������&V��[�K�����X�E���H��>�sFt��W������v�lO�k8��}���#GG��}9�;?���׾�������j�t�����	�echot��6��6�u�sr��腟7"q�.{��W�<z�I��?���nê�o�e���3�	;�xS)7KX��q|Hu;N"b.y5oT<x�ќ�O\x~�9���~2��?6[໩�h%��ɓ�zM¨B�3�"���,�+RR�Z���J�P�P�r`��S
Z�r<�{!E�,�Ѽ������!ڋ��('� �Y�F����F��k��M���/�N��e��� ��?�)5-;�˷�B�m����|�T+,�F�a(��pYZͭ��z��O�3��-P|����V�/N� �t��?��7��χ�?���>;m��a��F?:�?��������𝛷!���@�
#�i�X΃��0��9Lm�J:�TQdIp&���R�2%��R+��^��B7+����kk��p�L_TZ�a��P�+�2���A��oidD��/J�K�����F�0�40D�����E(���$�)�۰F$���<yD�/:T滝�q_`�j?������}�`l������J�������/)��3i�r>kA�����2�>�Twߜ��Ɂp��;ܧ��͗���?�������u��?��7�;�����o���&�<�0[�љ���! l��E#CB�*]Zys\��U������w]�X)�؜V"pՃ(��.�q����Jq��_����j-`iC��Gy!�P��@:w�g�y�@F3
 �oدQ?�H�y}_C�)C���k'��]�`lU>͂ �YHQMuU�[�bh#F�U����yviԯ�r8�&�u8��gۖ�4m��tb]xk�*���N��!��u�ƴ)Ć9\� V�������r#��e�Վ���Tv���! ���0^�
��A�N�Z埥!d��8o��q�A.�>;�(�C������#7��=1�3Gt��V���z���tOރݾ�~ë�'����u/�x�3�۫#�*�tp�@X�=��^��C�z�e2m�&]�����at���
���;^������3��{�S�zVǷ6�N!Es4�J8U5Jz^0u�
#�T饦Zע2%_��v�@����8a�Q�9?P����UZ��Y�I�`���W�_9��Z���GZ�ô4���q�]"��<�X�D@o�'++<��2��bqժ ��_.����{��4<���Q��]��+mn�}���u�*�����y�Gva+��^� �C��	ۺ��@ir:���]u#�,:��3k�H/V�G
��C���˽�<3�i��;�����w�.���� >RX���§�*����"|��?>��/+��C��2�{Օ��_�uh��9A{`�Ț�]9:�68c��ͅt�W�*U����[�֮�We[���SRYRvL� ��.��3�_n�R/�_z,<�5�m/o
a1yQ��e���E��)6�ِ�Z{����"�5��U<ㅋ�/�J���pfg3�.��_�h�o����e�ё@膷�����[E�ϯ�������o|�/�_}�[��o�z����8��/��ڇ>
'<=Gcd������S�a!�Dcš�(��P%�uk��|��Z��̳V��r�]y�+p9�r�0ժ�SSC�ூ�@o�Z��<>�0Y�)�����y�
_�� ](r�A)�{p ���
�_ Kǂ�%��y�9҆׆�?�����P^�|x��<o�����_j�:���'���O챊���c�|&�:zi���B�y媶E9l��,7��<���F��_E[�Qյ~��c8X#f�=����u`x�Ah$YZ��ܷ�t�5�N >|����y�7˷�V3�OjJ���E0]��#�j�)�ji�(�SHԢe�l;T�4?�׏����Q�#��$}�e��]��l������u����!4�8=9�����]��"��׿���7��^�\�u����7v���a�����z>LM�ݓb������0��c{-� ��@!�ӛM�m�w<q�|��_���	������n���඿��+��K�$�qё �1���]���e%�]3������W��%�r��s���e
�@6����e��8f��#�m��]+��; �uI{�T>U��e���<\��/J$f�C�iG�'bE��S�\���Y�Ӎ�`[L�A��Y����Ý�ƶ���0�\�G�mE[�r�e�K�-��H��W�_���v�Y�Q$��7cPَB7Q�6�*���8�����O�;�̘?+MV:�d�b�1&�����-M�v��d�*���ˑG�C���#����7�������-x˫^7�:8ݔ��O��{>��oB��P��0$w,�4�kһ[�6�UY{Ce$�[����4l<o�G%�3AcB��ZE,3��Ӳ��_(����O��Bյ��I����J�(#VR�[�^�܋ t5�:���$M�v���H�Q9��-�_qYѳ��E����xe>� ���a"�X]õ��il�aQ�6)S8Ь����F��^>gy���+��	�w���I�!��1[����F��	_[������
�����������>��G����]���BJ�?��D�&	�"Z�aV���ĪG �Q�1�{JQ�<A�yy����{�d���������Fb��e�ӭln��~95(�Ր��m!jJY���j��<T��W�
�k(����2h���<���Y�c����n�;�dMU�ϠB�9ZP���&ר2B�4���M#��z�Θ�6��+8o��1:8��Ҩh?�6~�Ӹcw���#B���j^8�*x:2HL��k[��l�J짾�>����8$�q�8�~W~_�א�Т��q���V9,����ѯ���6�4���N��I<@?s���a����]�)|0�2��AU:xLq.��^��}V�ӕ(}v� �ͶЧ��n��S�{'�����<���co���w�^��g��ѐ���*:w`?T�E|��UB�%�-(ZP7�;��(^�G�cӿ!}��im�c89�_��c���|���?���?�ow���[7����q8�3б�CCHy��{�N�2��I��J f��OÝ~ �F9SJ�LS��[�(���s��^z�A�Mú�����׫c�i-P���D�Z� H�߳W�u *�*�}��6Sj�\�J;�`��3eC�
��A���}�&Q�Y�#u�T;0b�8����w�}����<�Z��ؼ�/����m&�����>���rPv�!��+�!�P�]]p�f�=0|�T��g,�t/����Jt5o�\yb��\��[�լ�����3^��ZJ��嚊.������,c·�?��c�_���^����_�����?��c��'���nm����tC�1o�c��a	H��)�Ƚ�i�g0�.�w��]U�I��1#j�疤@0����JCN+sU�ʥ�T������K�"�/&" ч��>Sp!�P�?y�Z}@��q�y^U��4�i�^%h��F�؁$4�<���e�����A�v�e[2b*v��fO�\��t�~�we���.8�(Qz��1U�<=�,.[ixV����R|yb��C����r�.%O�a�r�P<z��Ǿ�����R\[��m��
b��̀�ݖ��	-�6E��@%ƌEV*:���쁥Ip��`�Ρ�	���l]�^ά����'66�켐��"�<أ���¡!Pf9_dOHp�r�f�r+�7oa�A`n��SN���/��a-����p9o-OC��ym�`ź6*����Y@�Y���B��M��K�M�Lò�y���|Iw�����i���""M����]�r8�����&�D~f�N�(�-D��8�8�6�d�+��3*#��g��p��J�P=��i�=��5{��x.���sm�'85T��
D���Œ���|�c�����ڻA�ib_un�î#��(QL|��Y�����B]���~Mn*�@'t���ҕ'B��'�)��!��i�D��ɾ�{�Hæ�Pv���k�pocO�ܽboz��'~��#oz���χ��=�C��' ����j��t1
��.}ƃqɽ+�`��8����t����W�����<ÿo~�q���}~��>��W�w�;7n�znl���
8�D���q��~k«�q�͑��N���C�z��rBW��B[v����!繤RH�s�JB��e����s��B���������޷s�)�n���\!Y��q-G� �~��[(��^s!��J�v�.,�H;@4���oD���[i-ۢқ�ʶ�v�f�v�Lk���ݗ��m͠_e�M�mk�U�UPu��c2F[�����o,�Ͻ.�{�Ħo+.�<�9NГ1���8��ħ��՜JS�5��.�w�/�#g�������I!�\�.���8s�2��Y��[a��3�:�9ΨW�(2rе�
���.9u�ͣnc;lL�M���߅/|� ���Ɔ8�7oB�Z��Wb�бM�D�/r���ј�=�U*:��@���O̵�.V���o�����lSRzV�����P{l�7d;�h�蜇_�J�g��6R��z�lDRD�qx�qs�e�lq� }3�K��o�
-^4��ho��;y4Π'q�*>ǞI
v:ɸ�I��D���x��0[L�k0L�@�ߊ;.R�ָBU��i�*�}�t6�BT]T�zLC�Ӛ>�"<��\5�N��btݴ�ץˏ�ᔙo�2P�T�+B�7fY���T&J���^���+�9x�t���>�r��S��%�-�`���3f�]	,��F$�G*Vq�B��o��'�PʫzJ��0��t>$H-� ��|��������v�Ha7ˤ�,w
�_Z�t�@Yh��&��O�
it $9	ڊ�ȴj#OvJ�V���>iG� ?������4=d���m�~�Fp��
/�&�������t���E.�,��(��jo<�~m����ԍ�FQd?�SfC��e�9K�/R#�jC�
��M�Ԧ��A�W�L���L0�E��;���"��>�ً":V�^#l$W�0O9�q����������y��]o�~��^�x��-��Yn��)�����U+=�&b`��HƁ�,��q�U��ڔ:�<Zif��S����ǟ����c��8��G>	��oÝ�N6��ꡇ��QDp(�J>���&��[����X�w���"Z�R>�.��^=g*�E�/���g,���\\�x.<�����٢�w_��p��x�0�����ɪ�v���v�j�kOՔ�xo�l&�̈́ ��j6�t(���*�1��<���.5uw�&?�۪�y�\��
�)�v�;�l#����-��0wphݩ:�O<&ͦL�]�it�R����s�iW��ȃ�<B9aO�R%ڄ�����"B�b��^b��P�4�9�N��k}p[@�;�'\���6U�|R����e�W���~z��a��Hy��6z����qDh=�`ǽ�.��:�%�7��p�3(�]�o,�!����;�i�ݣ������d���S.�n����Q��K$&/�����9�}��K W 5!!�zi +s ���ՠ^��A���ycV[�S��t�2S$��I��Ά$��ӹ�R�vฆKr�{�n�U�Db0�J�V6&��2�����re�>��:|����э��q��BG����k�I�I���7���oͳ] ��V��v�U�(���㧵x��T�u�h3�44���rJ�I��ʦƃ��5�E�)����̙�|z���q���5,gUf͸e�Ut;L�.�����l�� �ZnP�s٬j�aSU�Ԉ�*��F��(Dh����k�K�@��8l�]������[�'q��v�����,R���ď �4m��Əq�pM�&�LUN��̣DS�`�ެ�ڴ��\&]�傭Tk˨�JA��r� �qk�R���4!���2���M!�m)��(���٧����8S��:E�ؔ��?���]o|5����m�{5<r�&���8M���&h��s��un���P7d�k?�x?p��qSO��҃�}��ړU�'�8�O}�Qx�g>����G�<vr
G7nl�^��Cu�b����������F��S��h��B_BY����46ڱ?�.xp%���*�Ѹ������2r����3 �pU�p>�^���Sg�C�f<�TJ��e��o^̢L�����L��[^���J���ԍ�R�V�e���+S��g�D-�G���t���6Se[��|�~�^?���K��/��Ľ�ؘ݁�[�q�2�-�FΣj��cW�]���h�y� �G{�(2ֱ��Uh�|[~V{yMXKay=�T���`)������<|�Y/���/�Z>���fнWѦXe�D�|tp#�T"����
n�DߔͤÒ#��,euL�P��a�w+���2Lk&�3��^���SjΤ�Vr�r#�rC��ع�����a��d'�3����̕�gר�-Yv��߂f%ߓ�I��K���>G��%�k�k���8g��q�%NB'���U7����Gi�R'>�oA���I�X�7���R���F���-��Ԑ�8�^���ZuN�¸�Gh�l(c&�ČBs,�s����y�Hd�M�5+b��a��H+�ؐ媄mS|v<췃C��sQh� ���Յ {JO�8j�.�綼<����nZٝ"kC�q�U����xV,�ci*M�U=�$]DS�u^Pi����x��L�jC��f��Ciw�kpo�϶c������į؉�c�� �?������Dy,m!\�~�^����*|���(�]C�C��6�H��R��v;ēɟҦ #�n�L�n�zX$�H���n�u������Y��u�ï���]Bv�13���kO܇ۡ����U�7���W�
y�6��U� �NbY��5Nb}=d���Hף��k7:���!���C��.��Goل�����m�[up����o|~�C���O��?�5���{ ܂ӣ�'l�6�w�\O��� �q��,"�#�Bgic(�@�Y[~(�A-C������4���_<I�do�6(��|%�����e t�H7��I��%���Mn�c¶Df��'�wY'))T�&��	��E:rQy���<��s�W�&��
��m�z����2�"���_�Ұ-@��6̘�>�6��a�?U�C�I���o�X��8��8�C�1���p����}�~��SFo2n|��%'\���X�E�C;q�v�R�4ک�*궉�#bG�$*Z�����'G��@��tYW���V�Z��F)�G
�
\�sA�R��o�����,�Y\?�$wH��ǘ�
%���~�5�r"�hH�I�kƅXQ�>N(����n#{�3�R8/}�LO�ǜ����K��%��7�	΁�+�K�K`��>:Ŀk��J;����+c�6��Ό�.U�I�YҤ�������:)��Ӕ�ea&�G��#�2���'W��nE��a��96>�{ea;��o)|�!l�bٜWUݕ��D����2��XW��L�r�R�!&���bS'>D]�ZB1P��9x�F�>���|P�wc�����kl�����K��
� �
�H�d)g!���@�{��'�5$�0�!�O(��m���H�*m?��`mY>i���lZX�D��Q��!��y�d�c�S]8���'�v����V�bK�����sq ����=�fmܤ� �!��I1���Q�\3~�;�����3w#�:�.�C�Ǖ��X%��JN���='���"��A�B��>���E4�*��v�M�.�e��K|�3G�
�}����#�7�����<�Mx�t�}�s�'��N��^��g��7�owO����๡�ؐ� �_�/�?3�:BE�ec�>��=|�O����������|��O��Uݍ#8z��ё��u�G��G�
c����^�C��N��Y�-��*R�6�nS��Tm���5h>�{��t&Y���>���59��]�7U-09�\���� ���%�^�V�MP�H�vȮ�҅"�ț�K���o����}�t�&{d�i��/�^�C�4�31]m��El�`)�����=Ce�L�$w��]�FҶ�}v�;��d��>gm3��Z�$~�%H_��@�)| EzR�}P�8��:.��|î]m,���X�@���?���E���©ɱ��f�*F=����k�y^w4ѣ~^��3�lnR�{I���n�g��z�Z�����|�y�z����ߡ.^��{I�Q�+�ՕjCU��A9�F�7\e�ʤ��}��r.+{\�a�����az��E3��r�3���)ЧJ�&�A"pT^�p�!��CEސ8������5�a,�^Z*�vvɹ�F�R��Fi)4pܰ���bS����h�ܣ\�1�e��,^�[�|��d$+A�I:s����m`#?KӤ �1�75�����w>�v�ƨ�R^�H�X�-�P(�\��DRHK�WdS3�:��rX�6�xԅy,����s��kĽ��Y�y��%�>8hk���A�7󘢤�Bo�ݖ�B�[d���Ui�&X*�uɼn�)'�0�l�'p��)��~��<���/�lܫr�0 hҽ���f�n��45&P���l�aN���OئN��B&�L�j/9�Z�I��%db�;0WH�o��g���Ћ�=��$(bX��/��l#t���/��R�V�P��R:�g�j��+ȿ����L8��E \�a}r
��]8���܇n�;��f��7����WË��0��]��M�M��p�	�0���#G+��:M�KX\�!�ݤ�[kH��7��Xl������c�;��4|����Q�no����OBo��VG)��e�K��j�19�۝ ��ə��t���gϽRo���%�1��S�E1_����)s��E�bzj���)��^��E7��a�y_X�{XEj�'�������:�+��E���A:Z��(��P�#�6�:��P�z�$�\��ѩ�n\���ƕm����U9i�vF���f"*��!j���c�I�g[���	܉e��Z�? p7��, ���>���B�	�@����_�2)d��}XRR7?$�M�V�����>h�{��F�L�VdD҂��3r#�߲� Pv
�P^�g0�5J2�̥3�339�A�}�K�c0IV�ZyA���8P�p��|��@(�:_��C�6v2�R�|��E���ތ�*)k�#��</��EZ�2�w�t&مQrxq��pu鱩�'a Ą+#9Z'&��W��hn��mZTe��<{���(:t�[�4|���"��g�O%��)C{�co���|�̰��=W���~ÆcȟQ�5N�(�流�K���%ҡ�G����O�rr����O�>�O��P�J��S�F\�>��"#����$�S�r�x�R��������h���E����Hn����Є����٨�4_U�4��&�!_��D�g�����X�'�?E;Q��4]x�n�ͫ9i�/߰���$.�v�rn;[��� f,K���xu��O�����I����.�d]^;Rv��䆍6�o�t�:I<�r�ؾ��-�Wٿ�W�����61��ުQ����ߒ(Pf�t.��@*k~�8��F�KZ�I
eC�Y�l��K(w�B���E9�)��ɽ��?y���o�+���;�o|-<�ᇠ�G�D
�$F�a7zH�{ژ���=5 :�w���}��^a���g\��RX^����ؤ�}�	����_ÿx���< 7��t��w7�\6�Ǔh��r]���Ec������e�ʝڴ�F�(x�xbrц]��������%��,
}�TGt�q)קx�E�#��������E^���$c8?����6p���|�-�?��ڹ/�^x�q��!T� �T�{T��f؛�l��Jo�'6�����̷L��E�)�w���O���N[���j3�ꚣ�O�5K�1ܕ]������~Opuѳ $;��OC�;݊�l�[��x�=�K�;�DYl���6�l�jI�:'=�d��i���PG��09k�q�����YÄ��<L���w���神?�#o�q��ȓrClN䱍6H��g0��? �x��،��`��!��P�{9��8��@v�� <��uQ��5#`�O�]�{�u�z�X����F���µ|@��lv��"���nTQ����Z���� 6��;�Z�r:�ً�%ځ6�Z�L���,�$�2�F�DA�i%�C�sK��(5�Rx��+�� ���6)��đ����a�"p@Q���'ǵ���X�q�	���urzQ�"���)����.�Ҵ1���ٌm-���
CB0�h�+�m�d~�L;j�̦5�ýjG���uAi2�d���8�{�\�I�)d�j��@?=ܱN����-�}1gT��<k����sfn��]�/z]=�AN������0�s��R⁧�΂����:4��22���P��^�BUX�rJN�|uJ�{���1�`��71a�po��'��������O��;�G��:xŋ^ 7�Vbw����!�z;�w�����t�D��H��C��I�5_G�=;X���.u~�f��ic�08�?x�n>|�Ϳ��ݯS8Z�j���u]ߧOL��{��m�Lk�&\�x	��ٛ38���|���EuD�ʁ v���ޔ�R�-a,��(��[��ֻ�.>�m��O��
P��kz]mIqV:A"{Y���[Jٮb(&>]g���X/k�~�b�yC��l&���S��kF��-�A�0l�H��걞Nmٙԟ�Iz6�4(i���͎^_
�8T�U��L�����}���c��p@?�*'�8T��~A��1���F�_{���(}� F1˧��}pG��$J���U/1T��%�g��l�i
Z:ܾ��G�n�#˹�	��͌:�i�Y��n�ѵ�,!ϖ���^�5ߦF���(H��,1˗:��:�+[����=�шX���T�nRr�几J5�"p��#�̷�E>�e<i����/?�����xЌ�8�C����t��6<̡`R��$��:D_,������W������9K����-#M~	s~�ڡ��7o6�;�#�広f�<�)���S}�y(��z�7�H����ONK����H`�a�ޫ$�4/=.����`ߠ��PE��oS�$������A�m�?"ΧK�ͼ��[lyg'�WX� ��hT[�c��h��<,�\] b���XG��L6FJZq6�z�3'��ڦ.�;i���6���.�@�&Vx"�u5�*���me#��$I�-7��yt7iv�Ф��w,����t�қ�a&Ө];� �c�Е@�)2�=Z#�̛�[�#��}����50`�۴��<+������V]�~�څ��5�h���4���)ly�,i6}Bnt�Y��Z"mi=��(��B|���>��?YCw��V���<���������� �����_��6�֛��t��0�N�Փ
��P��;3D�Hs��1݁�Q�t���#]��@z'�V���=�N����Q7��ףώV��R���?��(�C� �6*��1��@�"g��B9�ۍܺ�7
e(�<�r��x[A�g��X*GZ��������$��C�M����aE�����C���L�/��z�λ]����1��-clg�����|x(�(�%�\�b�D 0$K����ť��鱠�Ԥma�����LU]�<n�
hҌ���pK��l&k���FZ�g�׭sF��@r)��U&=��}�N���3.+� �%�ہ�3�_������g;��d3�e��s`���UQg/RQ�vM��?����Q�iG��E�����9��Ɩ�h�����1���He�� u�VPº�Ƙ���>҉J$�Ғu�P�I~���g0t� ���rS㒂��,�z��(guJIN܁��kFe�gq�J�k�`S�Zv�Jl�\��fq���Ǜ��n�S��)`��G��)8϶���l��}@(��`�)\��vJJ���YX>j��Z��j/^٥���M�Z������4��Ŕ$-��F�Il�
\X�����'��D��Iꏦ���x��9���<���`��*�1����(��6=��Z��]8��ϟc&چaoj��|R�%b'��NsƊ��x�ذ	Z�� �JF��<��Y�dײ�r��K#����=Z0�U��y����`Қ�r�k�V�#
=hi0U�[���+Yb*��ٱ�䙗&xK�����1�F�2��i���ur[�,'��:�v-(g�!�7 g�<���lrȷ�K���e�L�����Ct�'�d8�t�jd��g��?�#���&1�t�R��[�.�i~�)�F��d����!Z�g�j��6:89]��;O��Sx��O�{�����+_�|�}�ᕕa��0����;�}���j#ݐ�1�C��� ��_t�`�1\u��W��Y�b�}CHF�ҙ���i���[+8:B8£��u�5HףW�@�2����	�>��V>r7KMh�G8�y���1���������ZVh+#�ș����R�:L/����!��E",���� @������E �}�'<r�7��a��h�ѿ�^�����S�߲���%Y���U��;�=�tǞ`����G�u����S�@���H[�LKo���;£C�����3�׏�E�ųs��a�k��ۘ��[N~
ܧ�>7�5l�]��O��q���j9Lo�o-�jöS�Ú�{�IYE�}���������o5N�Ev�hd�-�%0;3��3`� �`P�@ys�ø���$����vZe��0�̔W<]�Ӓ��!$��e}�C*��VئXl��+S}+G���]��ȣ�+ ��8T���q�2g,�f%"�+�~t�j�	@�"_�"��~b�b�v�Rǜ6�8t�y%�h�3��3�Eq%d�Wh��t}���1�T�J~g�򘄶&��~���\!�� ;^��75�ª��%�g[`�tzmkuo��@Z�V� ��P,���S��Z-a�h,i�� 3�T�#���\�\kVSe��
W��C��9�A��Zt�7�7G� �)=h-!%�T��hRe�J>P;o��C;�C~D��օz]:���ă��yx(���y�^[clږ�x��1�'pa>iqh�o�����u�qF�엇_�~nZ�rU�ׯ�h��_�cN�pJ�\C����F��CBu�J�54!h[)(e*�yr�8CgV�4�ڶ����.��6�o���RZOM`�	:�T�5oT���Q1�)y#�C�(Yw������~�S�{���g?����巾^���#>�"m�� l��Ãa�)_���&����
	1���@�Q���=���b�}u�&/j<�������<�ps�Aw�G=$]��i�a��q�F��!�Ѧ�n�����u!�w���Ft� �D}� ����C1��QG!F6�6L�'K�)gy�7�t�ЖQf/W3P������R�C�?J����<`���2�k�Ȗ3�ȑlt�v�ќ�Qnud�W����j����ڮ!��nqx��eΔ�"R��r��uC��v8K^������B�4���-d���Weߘ������jUa.'��~�-df���>�a����G36-���/���y12N�.���됼��2�=��;����C�{�7^�u����L4�2�ǜ�dm4�h*��E#=G��hn����RΛ3����E�-���	{DZ�����0�3i֏��Ui�F�3;��{i/kO�#Z�~�"qA�THW,���w����ΚKz?VϜ���^8@T�� �ۂ�װgh�E[ֆӳ��Z�\�z�T�Ŕ�ǅ���(�s��)�1,�vѨ��`�0ŭ~4G���x����8~^��%	4"l�J+�R�9�Xy� o���騠B;7���	�Q>XS�`:��iDx!�/2�+T������޷a�ק�j&"��@u~.�IZ���@�\֩=�%����f���^е|J�/ۑV��,8i�4�i��޹�uq�p��q~��_w�i�^������D�UZ]���=,Y��M��4���\K�x �(Y�8/�]�\@:D? ��Z{N)�~�E��2hx��:����Z�E`G�mc��^Ǩ��<�|�wN����k����~�����׾����۷`�ʜ!g������vP�r>d�$[��G`���D�N"=��j��ώMm�!<y�.|�����>�e���|	>��/�#�������g��ԑ�H�]9�vJV�kS�7�-M���(�y#_����Z�ԟ0��yÑ��� ��k�E�q��9곭��4��rg�WK��hd�����������tM�}��$��ò�K�T����Qq��ʚش�8�8�y�����(���lr��4yEEY%d	�	������C,�Ȟ�k,��)�Q�t9�F���F�Y�'��	�[H�i#vǨ]��k&m�ڣ�\\d�x���"�V���'\vyq0@�#�r4�I�AM���h6����﹝�s��u���9��:�n��v�������>M�-h�bΘ��"�B����-� i7&�Z�ƞm.�����
RH�*?��Y��u���K�&Ujl+E��Mtř<p�Z�R�MZ՗�3&y�+o㥶�ܢ��>G�`RM���s�U&�Č��  ��IDAT��h�����,g	4��!��9�3.E��g�x=��p� �p8�S�\�\�2�W�(,��0��If�c?���94�T�#�s�)>z0�(���{�4���E&]���K��銰M袞����,�K�����"�v�B�Z�yb�V���#;�4�O)�L\���
9F�!�Uw(^B8K�aߔ�g���,&eW*ڔ�* ��!�4[w��eLycI�O��ɛVr[�^��?���癰�f�IC��0Ƹ��{���aK`�;�1��/�m�$~�7���h�6�k�Y�� l�j^�w����`�7|�7\'����,����߁����k�\���gE':۹2ڸ %��l�N���,�6��ꋓ�ѦQekݞ7�J��7|�q#~�h��o������=x䁛���}��[��y�k�=����w��s(.ҺAZ?�`��Nj[�F�<�:�J�u��G#�k%0ջZEǉ'O��W��ux�'>���������{�����p�
��&�w78޺�P��E+��}B{�C�6�����G�̎C���Dq\�@X�����l+�Rb�e�$�׬'g09PM�"s?��d��%jl�o�O�|D/����Md:�Y!G��z�?S�Q�4�&K`7Ǿ)�f#p�r�C��@���R�T�����r�����r=�z��Rڡ���8Jg�tc+[:�}#i�� ���H��F�z��7���pm�:��E^�&�8(���$Tפ=:Aw���C�V��n-.9,�Lt)��&J��xg���M~�3���0�fr(�|�*4UY���m�P�3	y
�3����N��I��g2��gh��[�v&H2�
+��3�@D|�?��[�a���u	z�Ҡ
�bZv���'�j*�3a\�>�,���C!��k�ѡ��6BF���n�׸}]ҔXnے��W�3"=��^�WXw���j�B:p����I�Ip~pX@!�4S%<��ڔ�����޲��|��E��:)�(�;[
���%HY�R,?��X��em�-Q�+�j�u(�^e��M+�SZC�7b%�Yg�c-��)��jS��{x���_Q����߼����=�'������
�;���&�(��D��X����BFe��b�r�ޔ1kH�e�i�9���Jy�@���@�Q��� x'1�:0i�6Q�~y<H�����]r\�U;#��h��~���X;�4S�MS8xuz�ɩm���^��H����1e�ꍦJ&���[v�G8�v��_
=�@O�d�Ĥ�^,��<��7�e�g2j0��ց��
7����������r΃���Jn��q9��HQ����q#$K�ÿ'���| �Ə�(����^��g�Q�Ke��Nֹ�p���Ȅ��q�ё=;��ӿ�o��{�fխ���Jb��p�ɰ�2����dS��}��S��_����~�K���Noނ�۷��m��Mɛ7�N)'���7����~����5�w?��]�G�3�ŕ�@o|+OO��mM�r�NT���D���g-UҧhN�[V�.�9��!���	���z㼢��-D�yo�.�Y�w/G�$\�x��*'�<c}�
�7'9�w8���h2Q�EynAc�L�*�u���ޅh��U�ts�6���P8P��:Op��)�������ʎ��I&t~ٌ-�����#z}��6��,���{��H�e~��)�'��0Nw������c u��ȸ)-�\q.@��d���!�C�@� ��C;o�F��[�m3�噃�_�q�J�4�K�ԅ���j�U`l=t�W ����d�Rh��������������j,)޹��AJ��� �J(b�:F��~�N�编(�Phk�ڲ��ZQy�YTy�z�iM-n��:���!��g!�����z�(4��t}�v��t�Ȱ�;g��fKw]%�b9�ˋ4,Y�0��m��'���T}��t�g�HJ�JB����\&j��ꠟy��ۂ�	Xf��a��6��y�y֦=(�j�CSdMuH����-�ѵX������C���ԬCxy�`�^d#�F��J��pHoTƣ�����	L�n_�9.�X��rŖx�����j�T~��b�C�)IUћg�m7�:�Q����VZ��~�PN=c�R\�Z"�Q]��,O�-9��L]�4�I#i�8���q�%M�A��A��4�{��c�?�*�� #i�E3m[)[��4�A�oG�� �l���)�.�܄� 3.yQ_
̻.�,}�o�(f�?{�S�[/�ʶP&13���ʵR$'�<�I>R�����}��b�{rr�~��������?�����P�ic�'.�S�4�GW�
�A�"ِ,�0au��:������b$<�6-!|髏���G����g�C_�"|�~�'7yV������p�IXupcS���7�FH���(�/˱L$F8��烠.E� �ɛ�a�z�<i��"4�
b���1���<��"g�m��c���#Ղj��� �7s�@u�z�w.�=��ϸ\�.G���85���t�M9\r���l��̍��M�.����I��z��a��gPկ֦���|Sw��ۭW��mGǝ�;�� �W���^o�k�M���vǘ]4��Ϫ1����T�E;U�����Ss���>��}�����f/�G�@�X=B��%�9֦<��mS�Y�w:�Q�L.ԸYA��i%�}�N�uJ��2{��A��5�{��U1����O'�=�)Fj������P3P�ž�o�z1rҾ��%��UT�g�hP�"��cz�yȚ�m�??��#��Y^���#�G˔m�d�W�޳��̃�/�LQ�gM�@���ȾJ�w	\h��]H���k84TƗ�Y�L`f�Q�0�`�O
���挟Gl��`���Kk<�*��66��z��.,}��֠8�
٢Po��ᖰ��U��&oʂ(����[*�����{nJ�@,��O�[Ǘň=��^i4��i�\(+�L��i+�j��>+�YyHk�#�P	�j�4JSY�M닗�X���V+h-�g74i�
J���P�U�0&4�D�%b��x��V;�4UN��y#��FS��4I?�����	�W���_�o�����@p�����PՑ���q�+Od��A|g��ﶋ὿9Wm\�W��U�h���J|�)N�i����?�@�Aa8H�m��8���x:�G?����|�8ڔ���֢㙑e59�t�Cyk��\(i�.V��}9�+^Z�Mǿu�|�㟁_~������|�wໃSǍ���5D�Xo�\���H�t�9��������*544A�YD�L�����@�xӲ�}���ۃ���:���@@+o�����FK��������Oc����(�n7թj���\��|�m��Y�m�k������o���<Ý303"�h*�L`�ζ�Y�Y8۫q}�U�q�y�yJn��b�z:������#���%9����a��muZK�wu��4�{eOɲ#��\�n	���t�3=Sy�ŘMbqGQWeA�%�b��	��3a���g}��5��:z��ږ��<z��7Fr,�n�Vތ�V�`0�=��\�o��4]g��|��+
E��AT+�`����E���r��l?P��c��K�'�]�7��� 	%��凢�z�rM�aR�}��ρ�d��
�}u[�~�v�/���g��J�^vyc�8���rװX2�[2l���;,T�� ��/�a�JEX �l�,ce�|�-1B���$��e۝�G��S��S�g^�E�`� �3=xc��*��*h��m1��uH��Ay�i�k,�J����e��a�k�gߐ~� ���KD��A�X�3N��՚HNWr-QŴ�9��(_��J��j����Z.̧�5<yi_�+vkҙ�C�EXz�M�a)~dyx.�]��Jh��~a;m1~�)a[��^�vO'�ߕ���w�ͥ�W2A��m�viW���dʛ�"p@.]�,�!=�g�ڠ��p��=�f� ���2&�igP��\e;���h6���S�*w`����HW�=������o���NO NB� ���0{ ��� Bv=�+($]o8<��:6� ^�1�5��S��޽{��o}~�}����?�?���pz���Bw�8�g�>�z�m����|#��l�8D�8��=�5�-�c�:��G�卫��Ǎ�Nn؅�y��H��Q����%ozΥ%m�ơ�hRBс+,��h]?�~m���E��Y���*C��:9��g�-Pv	6�j+@Qߘ�uN����8��#Ɉ;c���1���J�JĿ�h���^�����xP9PD�d�bCi�4�O�9�VJ���c⮥���ǫS��l�~���7��,o�x1~�^t������<�ϡm3���#c��5��3`��8fB�����e:���3��v,/��-�1~��&ͲmZ�O=k����2q�&N�F��q�79�{��#�3�j�`St4����^n����>bV���{tZg�zU�'�c�U!���S�,���QЅ��$k���峬���w�M)_�K��p� ��l��2ہ�Bҧ�/%�B����c��&��6�T��Y�����Z������P"�>!�G��,�C�2�L�CY��T(��l��8a}UGfZ�;%l9tc��D'��CD\��d�o�W�ޖd����o�d}15U��H5��X|gd��fE��B�rE�г+�0�g���i�{�|X74ɯQ9<��L&� �o:zkL���:E��� P�P�O�s��f�����j���@a! .�gҖɆ
�!���Ri�*�4f](�@���獈�+xi�_�a;��o��M��s���m]���ݯ1�pw��fH�E ��Nw��׶z-]ѨB-.�8��`�U}�� ���w��s�Er�<���w��U?b�I�e��y���\��=ٞ�h݀�k�������ơ��_:X��������)�_����/8=M|e��.0�J1vޠu�����q;��B��@����z��ՠ��d��K��6�������'��>�U�ʓ����1��c8�V���F��d����'p�h�w��;���.��r7D�=�!� �����S����cI1;��e,.3o݌M�J�o3U����Oy��(5�ጃ&��(�,���4h�߱g�����R<e�΅1��Zݱ�r͗�y��L�'[��9�y����[ʉ����x�1��4�)/F�KB{�	E����C�� ySN�s+��'�9y$�!f^F�%���k�l%�M��+{�������t�9i
�M��/t�)g�d��=�R�y�%�Ҷ�}&i4�_��k����>F�"H��ϱo��V��+��H-Q��a
4�g���p��(m��N�|ͩ�Fҵ�-��h�!���¢��o��v�a�w����9�*"��(�S9�rɡ��*����?��6����,��/�]6&7%���(�/W��������;��-I����/���߷$Ǣ+T�#oV�vB܌��n:mt�Z��,�&�p�2o�F} ��=M��i'Gu���-.P*,�0�a�
/�6B�ΏN�W�\�"�!��q�ް�J]u[i6�eIp���cU�#[�}������Ms����Tw�Z�j��l���r]ML��A(�!$�|+k]TP)@z�� ��66k</7=K\i�Y�qڎ����k���m7J���ߖ%����e�="-�� n�c�Z�T
UF��Be������[�V��EbCTo�M�k�	G�d]�4O,�ϱ4OSx:���O�ߜ�[�g�����n��ߜ�15�d�f�������EIY![���r�X�(�u�����ɥmR&��̃�|��쵇_����س�m�s4���><�e�rc朳�S=v-�����#�֨}��ꉆK*���� ����R���B�B%�a�����/��^ݐ��.H��~�� �K�
:Aҽ8q��4D���;9��k�~>��/�|�����2|�[_��n�߯�`���M�a�qZ��aNtL�U��V��5���䁃�G�TԈ`�1_@�1JH�5�X� �1~��>2
����:�w �y��`)Ct��� ՚֟.+iQL2!�"Vk�s¢59W���f1]c�� ���h�>D���2��]�݄��$�GF�H�XE~)�#�p��!���>��dW�����,�J��sZ�!5�';]s)(�����E��X�L���:ho$�'��e�p~i�	9&���'�f����$��<�z��s��(7���N��:�cF��9c"�Kk�3I��؋eX�K�M��=�k'��z� �W�����J��&���\<�|n�r�T&Y�b�#,|.;�����%AX�W�֦F�/���Fg_P�C
��7�?��מ}J9/��6��¬�[u$�&�ܪ���\�nU���JW�#����1s��*B ydA���Qr<���-sG�R�ɲ�[��,e�ݧ#����X���
��#�_�(l�*Y�;��X�M,�b:�)3������H�q�5���E��$:��x� �-l�:�����vO�-.�Rs�n	�Q���\3b[��4����\5V����($n������8�J	� ��B��P��+>\q���fQJ�ң��q���7"d�BZ�@*�Al�B/Ѳ�L�mx��-�\o��z[��Z��0��QK9\q&qo3ԫ�� �|�F͐y�����Y�����g:�}�~��X�S<���%/�@���_P9S�BF�,o�T���������r�i�����@���)GI8B?t���+g��� ���Ϙ�ݧ��9mUy��Cʈ�EEx3��k��ɵ����Ul9�}��Я"C�>T�$dك�M� �ZHR��<����`uk���0��}���D�dzƣ��_k������q~���_����G��8|#܇���p����k�G�5��(���a��Q���\��D��c���I}�e�8,VJ����IQ���ٍ+>�J"�����Gqe�r����[�L��菢R+Nh^zzа(����y�ه��A�]��;uj1s63dvo�������c�@�p������dtG�M�u$�)��g,'ˣΓ��#p��rA����]q^�\{��7ϵI�6$V��4Q�-9�^��r��}��v*,�����-�v�mP�b�kԾYJ���C��H���{������}���0������%ϡ{	x%(Z@��A�;s ����"���Z�b������[��>%��e��n��Ic�m6�֓Ss5.�B�W�(��c(��&\��(�5bS
�Ӊ ��t��ţBa@r<EsA��Ń�thda�>H�2���*dg[5'�A��Ԃ��A��rq.����  �v]���E����D���:G���4�w����0�9�=K��J;p��k����П���BS��-������w,�(ܥ6�P���6%���7Z��&v���y�|~�v�B�k��/���.E���	��Nzq��@.^� �q�W���f2^Ȃ���N<R�V;�\���������6b�5w.�ws�a.�f������(��L-�T�ҁ��P#���*��e�W��:�9�ul:�8���4�1��]�.iǦ�Is�n��f�ې����F:��g��k�ޠ��&��_���DI�T�WS���-H/�9r�bˈC�3�0��4��
z�F71��z�1I��T�*&�x��:L72T�O�F`\��|�e2����O�ރЭ �J2��=�ÆpV�L�$;K~�a
v����>����?��?��ß���y!��nn�;޴��S�.tG]�p����`�m��AdO8���$�-o��C���5�`#� ����a��ځC�n~F𪰡���A�o�_�*͒�ݖ�|��Jv*=MD�p{pN{H�G����m�U]���*���.��솵��2^[��U
��vA��T]~!D���W���fy,���P��G*��ET�EYm�)M��c6I�N�tl�>^�HX��Ew�z��i���-{�}cq���t�/�ۖ�5�U��w8�ȁW���]'�ԍ��s_����s���u�KbD��I��P���; �{�0s�`�˶��G1f��>hU��G�p�)'5�(�Q�s��M��[
����<��o�Xd�Tɤ��F�A�%}-�h��X���,{�P�*ukڥbl���3Eיn��ǜR4�8�����u�k����sHlaW�SU�d�X�SBі�ZiU �_tʢ���-Z��]U�}��\�V�d���,|��K������u�����2�pQ�3�:�*���:�Y>sѠ��JD�H�;>��O�LuU;�b7�z�*�e�c��xA�W�:�"�P�O������׽ل�l���x�#4��7hњ$e���r�%]ʵ	V$QЛ�ԎLo��:e]6M�@���284Eق4�=L���{�.�2aH�؍ѯ��G?�`�#��h;I������E�4>���,ᣇ��k(u�h�k\�ʹ!� ��sO]P�o�	��)��C��j.��>��\�h챚,/��������o��wN��!]� �Z�rm�@��$G�:,�fC���^��G�o����_�g�[_�2<v�d�zV�I�.e8�<��Iw�pp��r��?�G˲�l2���(]��g����c�Զ�V�	8���lw�5�lL��nJs�L�P6V}�'��TȵyPe▥n�cvE����RPOԒmX����22y6��@HK�``��$=� �6�����'}�P�%
Z�����(�xQ�3	N�e-�ŨN=���4��8���f�6f)��<�cW�}N���O�����g~�賞N�FҠ�{�/Y���=Xz��SB�y���=Kh�Q6�i_�E�����ܵ׶l����`�>��sĮn϶�Z��Z��ugC+��־x^Jyr|�����85iDBt$�}l�J������1�J�h��Q֕�#����ځ�\�(�)u�}[ց�l�=�J��&Q�X\�ĵ�<V�x��A�.�n�b`�����?��Q�d݄�j�9��#p\����8��&��hcG�4&ڕ�3[q�߭�*�>KÉ�≠I]j9�����t��2���
||SR��xṴ�FJ����0Uw�y�`��BZR�"�K2.�w;�4�U���sO�'�1����QQz��[��sZ�5���f���<SH�s��Ap��E{q�EF��\�4o��� Msǣ�׋�&��!��T�3�/�v��b�w���.C�ݐ��I���{�'ێ�N,���~� � H,$+��M$(i<��<Ҍ��G�?`��8���O�pL�=���%4K(b䅳��IJ���

)�;$����)�SUY�ˬ�sν}���C����S[VVU.Uy�<&�j�4]���<�F��v����3�����N}���h�];��a?eP
`�h[���7�t���J�@M�@���V�m�೽:��͆m���-�Ue\�tYn��z���s����J ,p��Τ��|W`8���sm7�ޙ�ټ�����}G�z�Y��׿I�}�r}������Sv�v]n�c��V����[�Я��c�޷?J�����<��_~������֭�ا�R�v���c{Q��بKk;��z�{���0���ļ;�}ͧa(��q�Gf�������ؘi�z���I�l�ƾ��p���x��!�S���l���u<}B�N���Qe�p2}��eV�*0��c��2Z�wZ�R.-d�~3}�B�RQeȡ���������$iu)e��]��佐�)�<y�D-/�u�\����i����E�JC=��r���L��Q�v�½�wU���]��J��/+��;��n�t�a�c:c����h@�<�[�4�d>[r~ߕ�l�ҙ��u�LĤQߖ��m��K�V��} ����zf�k|Ω 9���g-\�r�F�˺�VLV+��E�,����s�uE�u�is(\��T���Gc�C�N)���걋<�W��˴��!-Xv$��z�s����E�_/֚���.��ii�q���;Tr0+����U��uⅨ� g�����7<LE��������MÙ:p�P�;"D/���#���؛
�-�u[{��n�(��T�'�x�5�eԭ�n��C�����W���1u��ƶ 4ncW�p��d�b�J)� ΃��j�M�T���U`'�/�G�'/�(��s>�2���.̧�I�1�)8� �@O��sS�����Ǯ��`,\��Yp� (��Fټ|�ǩp�J��c-�ԩa�Ø#�m�66�D����c�:8�Ns#iV9�w�<V]ciڬ�|لZ�w�G^-��I�4b��Lk�'����des(�'��g���n[��t9kCW��ָd����Z�Lz'87֙�c����V�$�	�R�LR$d�5�RZy�K�8��s������
H�9q/ه�B��S�ۣ�\}�>�G��=r/]r�K#�.���L�\������Մh���`�a�z�t�ѯ>r7��^K���������I��s/�_.�p������,�U{G��#Z��~������9�ϣ�O#�;Q䗔u�ˣ�J�^�VQH���9vb�'���^�E1�)�G55��0�-���{���y�	�t2J���8�Ε�zrmeO)�k�׶���e�J����0/�%�c�_MP�mѢ�w^��+�7�s;>Vhy��dؙ��y���J5�I<�z���Qxx(�u�:�@�`�ۤ�B�eǑ"<�W�f|�f�z�nLF��M�E��/p`�8�I�װ}��I��R��`̶���E�u����Uy7#����6Fl��c� Ȝ��O,������=d�K;/(��4�iK8{�d������ 9�<��&��vj���>'̂"�fg��[��j����2�g�K��Y5�
}��"��T���(=m��2�o�!��z�y��u���񣄈S�!Ѳ���,��=�A��\�'�_��T�G~)'�n*�e)Иʸ�y�I�� ?(��+�uOK���EghS㐯T��g�mo�=v��\(Qd�:'��3u����w����h]Um"��1��,�QKȜ��-�gP��f��iyS�X�43��%�9ɋ����^���x"���s���f���H��h*��t�]�)kك�\ј�|ܼ�ծH�"̜���/�(+`�j�+)�L�i/(�4̭�:����\�������@�oaĵ֘v~�C�l��!�ŋ+�ר���P}���<L���B�*/e7���30r7 3��k*Ω�g>]��4qи�5��q�4r�~᧙�t��G@����e���ܽJ���L܁�cҰ�����r ˷c�*'gJ�〴�Vj�X±�v�7�Ne�YL0w�̘��}�s���%G6q�ϋ�:8h����;�p��=�9z��@��ēD�}D����'}��)�����m��);����~p������We^{�f�{oy�ңo�O}�k�����ҷ_�F?[5r��A��1Կ�wYl���5�m�}�����dr+zW&%�><>ӆ��o��$Ա !���2$�4I��)����B3}zWʔB�	�爃T��84`#z�r�6��X�����6��͉�Y�˅s��٨����4ó��Äӣ�i��M�֏4S0Vԍ��	�xCa�/�5�)���<�����zP�c��8��v��+<�bC����7l���H;���Q�5��iDu���Ɲ���:4j�g�Lc�蔝8J[?Ɲl�[������wL�p�aܢ���ݥ�s|}��J+�΀Ԩ�i�~�� ���s�[<~�!���V��Q�J|��R?�;��u�u�8����?f��K}͉�U�\֩�`|N-k�DI*9�&3m})�T9�F�_X%
�������eJ�z�q�y,!\��]���^^����
嫾�b��,̦'�>tּJCR��f����|^e�#:.��D�z�~K�y�e�[���<���
w2����LI.й���z�1j�?Z`-ޱFfż��,ǔ����C�ZȎ����Q)F�����Mݏ��jO�ZhQO�x�o|ڵ��Y3���m���՞����J*\�U����s�Z���<�h��UTƐ��ޒ�>�{�h9����wȝ��ਬ�낮�	����jrE9g���8C�������'nxf�iP�A�q9ą��I�kr��,7�Ҝ̏`ա��r��8�N�4j�5pi
�9�ъ٠���a~�i��)g�ޢ�5/F�S�v�,���ַ֯KZJ��F���e)��.���']հm���6�7r)�N�-n��-+)k�y֢	��2�̎�ԥ�I��h�ӏ./�����^q���{�#��]a�NF�`�ɽ�7#���Q���VP�i1\��yZ$9=8Q����o��Qz���7��	���D����'�����=�/]�no��p=
E�p��_~�_�N%�*��b/:uds��d-4�����x���-�q~��Р�5�Du��"vԣ,�t�O~�T;��:���x�ٞJ����~�|C�'޴@�9�Z'x!�uY.��"�@�a��D����=�̰+Q��7�bx�v������8��+�(������b��ꉕ��0��@=�S��P���c�N=7��6V��k���~Y�,�b���Ҍ>[��l�F�a����Q��/�}�\��V��ի��i>�o�
�m8_����S;Y��K���ќ�k��sz��6nˌ�8c^i�/�Ou� ƕK\@�X���k�>�r��ѻ�6^Y�9�ҳM�됵�E�`}��1������CW�]��`�A
͙�Sɔ�Q!2�+�&����(X髷��,�`@�ӊ�$��B��{��'Ά�<�uו�u
��O����.u,�mP�c����>��F���#��$�M�0���l'�(�|2�D�1�����LS�W�E+�2�tH���H�O]�(��zCd�
��S�؄p�_T3̵0ڟV��A��z�����y�en�����p�/D䭙��_.�<���-�����㛭j'�1U����rn�F��IL���$�(C7��b6�`��R�]+��&V(ϥ�Rmf!�Ґk?;n8������Kn��F����LsDR���:�����UuZ}��ܙE1��иd�f�#�C;��c97^�j��m��K�K�P���@[��9c)���Ե����E���
�[�M'��ބ�e��:�UC٤@�vMx���Cy��4�Ԝ����п�"�ك��Z���9��US��l%iҳ4oA�E=�D߰d�ü�s��	�O6�\*�]�%}��?����#��~�ߧ_x�^�n|X�Eg%^>��h��1��s9"Ft(�xp����a1D�~��$��2���*��-/�������6��O����㟦������?K?;\տ�Bi�ם,�Qp���6�p�9�+l�t{Y_o��H�`Ox��>m"�!}���y�19����<9_��ǆRmRŧd�x.8�Y�窚�-��� ڞys��&ڑ��D�����,,��-T��\�&�>��'����
ֺ+�����=n��m�	mf�$kUHY��?�=�@��A���~�+jB���q��OL)��@=B�VJ��:�g����g�7���#i&4���!���Oթ�8K�YB�޴s�.Xv�k�.�s��ϲs��8�񢺯��`Ar�H�'wG��͡�q�1|aeE�8E��1*��z��@�8ׅ��ݬ���ά]3��3�|f+��%���%ݍ�M矢q�}��Π�$��/��Ӝ�1GW��8���9�©*��#�ɫ8�8@�N���UDTvT�Y/"8�v5%<�7��Ufk�] �43Q�t:���f��z�;�ON�3賑G���c���A+DYx�Ҧ�}]OW>�zN.G�7�>��Wk�f^�$�[s��O���8� ���L��t��ƻ��M�R��/g�eq�-�,UY��)~�-�1��LV�>�VZ��$�UT����ej�C��$[�:��#I9�<3��K٪�>�K��{�}�و��!SVL<�)o�I��l�M���L��(U��/8o��Nٸ�C�TQ�B�i��P�xZx��0��x�f��������-#RF,�v�\�
5D;��\�׉��R�Tވ��.ys�ݎ�6�7d���TZAS�2*�|#�*Gv����pi���|&~�&����*��	�i�;�gąq�9�.����{JC�_�×���/Q��O�/ҁ�vpw��C�ٶg����c=ܣL�&؊����a6���ضS阣����y����M常�1Æ�y�o�����̀2fd	��:ŉoc:<룃#ރޥ�t����>���?���3���n�����^w��8�	��=�����������|�Jtޠ�KW �*cw���]�Gw��f�����V�|�?��>����}����Џ����|�
�Um�"˥����ҋttio�{���0]�a��4��^��/�q��`�ʟ�\j��P�!$�9�0yN�|��.�\���:Ug5�A9p�k�eT=�ؑȕGz_��$��\E����qvi���Z���vB��q�JW���#�hs.r�U��,�B��c��2��\K�s|��;�[~k7𔚩P��k�$l~��x���2�"KT�}���ͅ��`K��=So��G�3j߬���S{��ͬS�$d@*ϲXh�����O�U}�"]���	4��g*���O�m��[��8��Ƶ�:��<���cuF�w�y�%7�hݓ³�1[!&�(؁O���`�%�����-� DHX�z7��]�Dm9#m���o��6>~��[���)��ؑ�c�4���I��h�{!�5���� ' �vN�{��x��F@��կԇ�_��q
t������=��H�r�~Uu��B�
t��]�;y��ŗ	8�B;_��r�J=ξm�eXˁ���$�;\����nZ��ǅ���5�z�I��]VL3'�luD�m�a/o{�{�*憎�-K�NVS�a��4ͰѢ������A���m�Y��l�=RC��:Z�061O��}�fnK��%�,����K����u��w�F[�z-mp(r�66��T9�[֙BVT�yy&�$�S!�	),{^@p�`v�|�Mr#������OP��O��ah��q�M�A59͕�������H��T]~$�b�d<� ���ikᇴE<�]g�����A�Ɲ����.Ư�7��Tb)|5�qۍ�Z��I�6r7no�bu9����%G:���b3����Vkcm����YFM�lK�U�I?�<��[�3���p�ʻ��	b8�\�ѥ蛇���?�C��?��ң���x�}�k薃˴�X�&C�	�rr�H<������w���'m�S������#�eA��s�a�������o������������?O?|�(8|x��?G�p{�K:\&�I�>S��(�c��D+)���|���9����86G��ATȔ��gZ�7tE*|�$϶dsɲ��4|��2�J���"ME���3a���³�i홅+`�o�"qq��3�x�5�!�-[w[��T�p��iR��I_^D�p.|אT�������6SaW݆~.~�z��-��M����&�����C!���p�������	g�R�7�f᷆M�GҚ�y1�v|.T��˅] yg����q �o$!������󮂶sPgr����{n�Ek �FL��CD}�D���!\o�e&]�YK��52�x��g0�m��25�|��H5c��]+�]�Eg����`g�1����G�`����>�ZIYE9�I�Օ�"��k9G��X�`(�%���%�K�A
*�eo�)����'_յ��H��A���
�v��1���q��c۪�y}^��	���3vB�k32ϑe�le4k�74_-W�|Պ��Ag�(,�,G���<�,�,Q��O�n�5'4���ÉzJC�O'*�9���>+"�`6Q3�	�`������%�Qis��<�e]��ODc�a�Dp�v��z� #$�秎�BԈ�k���*`�®Q�ߚ�(w���ӎ^���J�L&pӍR���G��7�ƏZ�#i��p�pw���F�q�c�[�cw���o����!�W�Y}�q���R�_3�jg��ܞ�]��*Xg9c���C{C�7;τ�C��Q�"�P[���Ec������yj x��{R�Ӝ�hKoZ�?ƙ~]{���%����xm�"s��,i�y:�':�|@_>�F�?���؟��������{��Z�����ƳK:p�����kX�z������O�!w�4F�w��޲�;����x�fzӃ������o~�~�㟣�|���O������n�BG/.�ݴ��O�1E�pqýOÁ��/��Z���Jo�Eہ��5��[꾒8������&�IF�Q�e��|Y(�<0��G�@���n�d	�+i���i[���b$�:��Ї�� �K��q#�^"׋è���q���s�n��f���!H�9=���a*�9J��#�9�}$tn.�m���g,7�Q���K?����Xօ�,ݜ��-�'���:�]���Q�P:��MFp7m&W����*mw�L�a?Qg����]T�����Ud��A�l:�q�� pm�V�D��Bp����Z��C���D]+~�4<���[��/��d�<	X���,b�j�m�0�t�𹔇���`� Ϛ�wճ*�ZRb��6��+��ʛ�*�1����|��p��⌅8�+�c l���jҴ�F����|�������s��gC�;\��nt��l.&z��y0@5��*�	~n��`+��?�����6=��捷~�l+�F)%ſՌ޺��tis����ra��N�4�-�9� �]n.|(bw��)O��Q�5�巠o�j\<%<�%T,����t5>���5!�
��rp^B�7����M�n#!�1aQ;���%���Ԇ�p����+�d����fY-#�)��b[�L�u4 ��y9�O��إ��m���������"m�՚iP��Kdo��Վ���C�a�4�3�I�9�|T&��f���ߚ3s��s�,�7U[�n�&�b0���r�vz2��K��Q�z�)��b~c�iE�e1���!U*.N�B����T$�.�[\�y�u!}�ra(��O{����먿�2��Z��O���$���=������O������;�.�*9
�ٸ|])vm���+K���������ꁈ���ǐ!C���U}���
����=�����������>��ӳ���n�V��C���F_l �.\�꣍1�t��N��LN�|�h��kX\rTa�;����<�/�!�1J	��V�Fϖ�.om
�=U�v�Jx���R��i�+ad�O�D�eծl�NA\���0P�P/�^����i8��M|/xmƉ	(+�����CY�U�ɩ��c /���({)�����1���~>Ww�u��/YpR?�����p�4�����N��h��<��Z6�e3͵I6�}��D�k��U��G�	�6����(��z���b�k�����]�hcT��o�"�\��mejֶL	���$�����%ʗ*G��g-�4�^�S��9tS	3�]��[2�)�F~����4�maS��`詸�H(XD��"�`r3� j�="�AQ���Z�'�e �;Ԥ�$`���4�zO`d�@_�zր|�u#�	�-`���Ė�ν�p��q��Lp���΂f�c
�����-�5�<[PNw�Q�|h��W�Dҡ5MX����T'�]y�;7�����B
h-�5 �[�T�+��d�~�b�VM���Ҳ%~+)
��QBsŖwkkÂ�	�8�a��{?Cn��Qr�0�(o�H+x�9�:`�vٓ�V��ſ���^l�m)���Q�י��ذv�����N��x؀fI<\r�҉s&'����e>�섊�\B"��Lh@�_�4|�Ls#�`��18S�g5X�آM�V��r��3𛍻[wE��oV�zf�ծ�A���Sk0We,�<�I�*�4�ݖs�U����#�����]�Wq�/"p�.ԣwz�VO0��Sj��u���H��7xB���/�S��D���xM�}�������O1�Pү�����#��G�ۿ����������z�]��k聯�x���D��Χ7���w�HG�SO�p�+A�|��9Z����W蕯���|�]��՟Ӎ+��F�}"��)
}���h�\R����6f*��Lc��O��tY�ū}��ǫ��@�x#N�{A����=�/eJ2\�a	g�x�C�#p�~���9.�ڰ��@K�3�"�Dzl;G����>
�mw��Zy�Jεq���!�Rj���s_�B>���\����t�𹭢�F��l1e)������	[{U�(Ҕ>�boݽ���W�����4�N�������Z4��6����uqràQ���m�֜����~v�oC_D��.��ǡY�E���Ι�^jy��o	0Br�p������L�U���d!�w��j�!M�|.ê�^��V{��^�hY/w�ed�,h$Ey��k��O��O>�"T�A�|��Y��=,QѹJf�R����ºT�(�n�Y����D�s��\o�z���Q��C�	����";��"����{�����h_�ω��qj ��y�b5^�?��9?���q�eڸ��h% �gH�9�Bȗ����e��*��˖;�'���5���z΁wI�|����J+���H0��:���E{(�U�ݴb��5�Z�u5�S�D��6u�es�e:���Ǌ��IY�#�
o���||��SE���A���T6^[�V���#�n���jF|�g��3����e����v}�����냈����=��Y�a12����
.1)�8Y�eOd�l�^�y`�$E��o��i~���Hk��d,�#�̴�c�!�t�-��t'{�8�F��=F��VZ�C�A���.�
=t'˭i�8��m���[ցu����_�E�x�D�(�.����ZmΛ/c��D��<޾���Bĳ�O��tq�ek�*wQʋȍ_xSUc.7���v�#E�Z0O�t)8T8:�t���z��o����|�n;8���|5����{���{�mt�ۣ�p�ɲ��]�#��C";���_e,��ȱ��_��߿B��"8X�kW��Og���::\��;O���}��t�K�%X�>��]�c��Ӽ+�I�''��SJE�SX>�a�?�Pr�W�����**2�t���zWi��bZ�+�f�겾o���;aYWf�4�Z#k��|���Z� <�a��6������<��K����a]��H�����lQ����]\G���.�kV��8�~���/}����S|�u���'�H;����ܪ�ҷ3~��k����`���u������>s]��X�~:͵po��O�A�w����A�9�[zw���_`��צ����!��]����_
&�K�ז̐7h15�1����#T�V"m�����o�����|M��WG	�g>�V>qsGp9�U>����]��4�1�� r�4Y.��
��H��%zi�I�M*�Oxg������:��@��D��Ȳ!��i�"p� �a�Q�j��'�
;c�s=��6��1@G�:Ѷ`H?�}"|.����q�t�p�&������A�ނ�t�-��9*�d��9
ce���Ƞ�PS�X���i��y#V��㛠���T�5B�f��7�+�=�؝��n!cr�"��ι�䷒�R�(�J뀦��&o�^�Qm���j^�����tn�a�&�樟�o�AG���N	���6�t�烞���x�g��
3-�&�<� �ߊ+�;T�Y�'�	��(�1v�m�O�z,w(�a��HC��[�c��u�:5��H�pg�'h����j���O�)�
� ݑ�¼I�9i$�H��u�W� &�b����	ܪj���\��m�t�`�'10ӄ�v�8S���`����W�#/��z��k��*�!m����e��\ϑ����[ܱ[CD��Fe�Þ"U��{�g{���>����!�׿�C���}�n=�F�|�=��z3��MO�+n�Lݵ�����w���^b�*��{8�^�x��}Y����9�z�ؖ+T]�DB��5��~Uz����щ��X��oks�y�q��Z���N�M_
CX���dOyUF,��	e��Z
eN��<t����J��If$G HE���2㼈kM���5�u0׷�#�J����ѭNZ��2l�g��l����J�����z��\9�"��r� �M*�S�
\�Ȋj	���э�:�tw+m���(W�9�W�N�t���ä^��6~���pG��4���A1N
D�5^�X�D�>��>����s�8.NIp��3	�TQ�Xo�5Mk�\�c����47Ѫuۣ-�Y�|�s4*'�F�v�s~�VF�Y��}wvB��,v5�>�Lr)8棝*;�1�h	�|��*p�z���40���H��fr*݃P�bJ|W�H&�)��a�7,У.�	���x�^+6�7�����8\�vsF]����BpF�2+~9�]��1`!_�P���fe�YA"��f�9I.���jm�r��-N� �L�T_�6�G�&�: *�rs����b�zx�t���Z���?s\yQ�@�/�kĦ�8�h�77g ��#�����N�+wF�b�aw���u&�Oħ�a���/��e�{�0���v.=���iɓ�ˇ�����J0�K�(k�F*h�,X�9"�]�}i� qJ�Z�r#F���?�_��$���U�������i�t�F�n�����iYYi�l��V�u��ʱ��o�(O/L����W�R"[Ioր�V�c�9\j�7 t�(:i�	�����lJ�V
T���@{��-ޔ<<� ��[�����=�����!}�w���_������'�H���nz��7R�j�?�[}��A�u�|t?��%]��0v):Hrd�)��j٧Ct��نK��?lQ�7^��.{t��1�F����vE� �(%����R��x��B��*#��Yf{��TT9b�QE�S9j�/�������M���JdBW!�p�i��/^���~1<o
�v���0��� :��IG30 ��Us�������<o��NQy�:�'��>іA=���cG��l��[v��>q�ȲL�}D�	2�_�����. !�������^�3��Ưe��F;~���O�L��1�h���6��4��Zk�������C���!�?gA�z1���oj���j�g�-���.L�A1t�\#m0j���.-���	#3m]��J����tU���uw'��F��0f=��]��v[���� ��K��q�	�T�0	X4�%��#E蛻"o�I�"������7��	��Z���J[��0v1�I����I�3�J���؎�.lx�sI�$�W����5ָ��\����V�t���P�כ"�Vl�U��v���5I���7�j��-�p�Y�VZ�fO��P�����m�]�Tь�xW]d��Ԋ�W?��ڂ]R(���H�$q�j���˥dlQ9`�B�IZ��H{H���U���dTԡ�b���M��\a�'�3�D���m���2�e�����iDҕ"��F����v��ZtN���k!m-�U�������DZ�L��v�W�p�h�%���*������'�[�jy�mN՗��c{�zo��j�$�`��-�G*O=C�Ɨ�9T.�:�����R�.�̀>��bQW���E�jd�x��ʸ���ߧg���O<M�������N���}��7<@���Vz��7Q燈˸��p�^!&1J��.�!���}>�b6ECZ�{W��/��r+��;ߧC��5wD{�ԭ��\�9�'D��48���t�������pEe��(��(L<@�2��.٦����
)��ỗh�m�ҳ8p�Q���#�X���O��<^�:�0\�����E8Y���4��A�����wql�]d77e3i
����۩F|]���;�twK7^S?�����4O54wo��5�F~Lw���k�Xto�$��ٚS�jEc�yxصC��/���d���3����u^'W�eMԈ��6s�XuM��/��Qe���H?�QmYy�9�����F�U���ir�DMy�3��+�����\�
V7zם(�$�.����12$��^#p�&8����g0�X�C�L`+qg���9��m���O���l�J�]Xf0q=͖	',?̐�n�h#��g{��2֎����Fa����^�����LkI��°Y�^ߡ��ө2(�';6i�k�t 	>x{a̽Ve��\��Rb�9{��s@"!�Y-{�Rf�|�aγfc�P��U���(L�8�۶�x�Ӊ7h������0Ze�5쳶B	��}�Mp�%ۓ�f��ʋDI�
;X[�+Ɣ�]P$4�j|)��3��vz�zʇ�!��:�`�W�}2�(���ׯ��i���xBs���X�:������syf��ҊB���0C���]l��7g<��V�7���aF�4��Y,����.G3p}%U�i�h����d��Q� g�c�(��5��j�U*p���0s�4iG5{G%�H�	���IʏӔO��G>H�>��8��sޱ9)8/����	|�FGS�G��7��o󖔲��Qy4�eI�ϭ�&~��Z������uQ.�/�7Qx687D�����B�!0�Y�h5W��>�te�����M���7�����;ｋ��7=F��؃t��7��bAn���v��������#6��ҾG�,9j>�ܻз����C��o�:}�ӟ��[��ʏ���}��o�L���U�����v�b�T^���VO:�x���~X�>[+�W_��ל}Z24����G��Z�5�d�`-�H���y%"�`1�cI��dv����{�H$�CGo�\����������[�#U}q�D��+#	��@�%��j�����Xyqy+�D;�j�u28��"��6����t֍tw���v$��vG.�tw�qi�㬺��Y84��Hk�i��<	�����n3�*05/B�#�^R���}quJ�Q�zX�W�=�T_�r��U�Üt���y��^\H��2<�}ё��d�l+�`�2O��f�q�k�dG-�'��|���%���R�l^I���))4���s�թc# ���f(�K{��	�٣������c�+���F�D��� �0�z� >��kp��V�m����C|��qV����H�-T��"��Hϲ~���s�m�1˨|���^=��gG|���i�ȁ#�N0��*M��0k�3�Q����#�?3�Q�O��E.	�4�w@[�`.,�Q8��_��!o��򔺔 ��m}�K�{CX��r����aد2/��lYay��$�v�t�%GA��k����i{K��٨?e�b�R}�Bi�A9p�b��g��
��	��J�l}�
�se��ö��M�zKK�
5a(v�9�ò.����^�E1�4�I��b��Su�]�f��A���$��^ӣ������(�P!m�G���A�`�:�Y�+�
t��&�S΢m��$�9^4B-�`p���	4O�#�Z[Su��P	�C��7�*�7�^��Ǒ�M�©�=0��^�ۢ�V�X'r ��C����<$홢fGG	�t�d0k_!� �w�0&�w��_�x�����':Lץ�K�����w��?�?L����[_s��G���v���.��C}�a�v����'2��]N$�g��3G��o�e�\{�u,�=ݰ��^w��7������>��g�#��"=��OW8_�)]��%-�U2�2��KG��6�:��%�#����A�le�]��	YƔ{��e�4�t&�\�Db)��¢�1(Ғm�ׇ&��C�5�ytΞ�+�����P��8	9m��s
cW��&�9�=Nvv��˲8t�%��H5F>���J����H�q\ָo� �vޘ�o�D�V웜��f�>uZ�S��e�p��:��a;���(7�;QÆ!�F�ְo6JS�Lk�[tl��K)��~���S�l��׆<4��A~y�.�r$'�u*�Lw�о]g�\>8&��y��49�/!o�^��h�]�<�Q�=���?�~@�?��?>���怿<���8ՆFs�Lw���-}�8a��c	_߻�WU�>���� ��P(����Ĥ�+c$�=��	R�^����y��9|��5IHE|�t�E7Y���5;�33���ȓ�8A�r�K��X�u0}���Tv�����`�+��r�vڰ��)�nMa#�U/�Lr[o��L���[L[0J8��Vìnz��c'JZq���P��cG�[��"�k<�l���c��m���a=p����}�L����%IqC7+���	6[�=m��v0�r\�|�1�)���]6A�e�8��ὼ�#ӄ�l)������}�e(o%*;'
�8�J���n����p����9��N��AU*n{V�;*<��P�+Bh��%�YY������q5o�"�r��뤑��kN=f�L�Ѭ�ZQㇸs97V����{�gC�G�ks��Iz0�x��4B�h�$&��3/�se��|b|L"�����F�.�Ń֕g-y�?	�7���Yތ�/`�Ao�Ή&8۩���L���~o�e�lDs��/��v	ȩ�!�?vc��>3�x]���gg�E��K�=�_D���b�d�G��ނ>�ӟҗ��4}��g�W�L��u'���{�M�Gw�z3��A�~�WZ�������� �Yq�~�ʫ���/�.�?���o?8�;~����C�w��>��W������������?G/�%��9�;ا�$���˔���L>�yYvQf0~<OA0��4^,c�Nÿ�s7�xy��Z�X"�d쏬E\�������� <>�
�Qt�au<��lt&���r��6}��ఁ�<�2�]�	퍒��3��4�ߕg����&�J:}V���{7�a��V��Dem�����p�8 �U�9ήm�������2��$�$E�����5�6���@�[x����?��,�_П�̱�:5�Z2hNT���.�>����_Ncd��xXE��=��a���C�u����%o��O9��|6�Ͳ(���Ԍ�:�dy�����L*��`r��K�¶��M
bW��g|%-�H���)��!��F��Rf�����D�cpJV��l�'-W6u�:{��7��2"'�8��H [��I0��N;p���s��A��������J���5�G��dQ�g�f�vAˠɆ�&dN����� L��S���/)*E�K*�ϖ�k׋ϛN�F��>z����x�	6l}Q:|�e4J�!"�06������¾�7�7�)^�;�oٙ�y.[�=�Q0�P�R��v5�3��<QyG.>+��\З�����H�U$�p$V�	�MEe6O���N���|��k�Ab�2�����d��嘆��;y8^xkl�>�Rk�ɵ/���Ӝ�9gO�Cz���Mk���J�ƽYg�����.˦��i����tT�l�ШjϩOU�lg,p0i���W��|��u�o9ءl)�!=���N��A�Ap����oeh&Z`�sC_l�u���KgW�o��|r(����6���u�6�Yp��!J����{b���_�_ڻD��=�Z�������>��'������W�� �瑇�{�W^�L��>�G1jF������"9qז��m�ӵI>O�u:5G���y�_�x�i��|�ړO��x���>O���G?�Y��׾A_{�y�v��Ч������bDb�x��Y��N�C��p��9�N�h�F{�I��2�����r6���|OyP7�x�쑛���n��s��c:,�6M��>��sB��6��B�;�p��8���
�g:Gƕ��2��z��8�SA��bѾ �k0�OW��z�͕=����'�6���S�a��s�������7�6a�ͮS�7f�4�cb���E�8o{`g
���:��f�e�0g�t�2cK�o/���wkh��Dݰ��&�Fk���\I�ݮ<;d�n?�g�nY��2�s.��t��/�j��K���V��"?�rv�X�;��*-t�.�&|z���':�R��ֻ��v��⬙�IJ�/���E!�cOF��Zk�R��'�0����^ҿ��W�M�r;wב�=�o#2������8�s��去�$���~�xC�2�����ݡ�<~q$��9���&p�!�4���NJ�p�#0RN�55�i�"H�\��?�Ĉ"5�'�J�qܵ8N�l�7r�aw	g�UJ�Y8qdv����r�7���M�~ƺ'J�C�^FBUv9�^e�v� <}���E�l���h+W�}B��Z9(��]�H8*��d=�������#TG���&�d砓���B�q#���»�<�hh�fU/u�sod��)d,��L(��@.U�G���U�Il�ժ" x=
�,4�]S�Q1���Ǝ�kyG�;��9�>�4W��m*�x�������r�T8�/W3�J��07��n���
�s�R����	�[�N��3���Y�6鬃?��^g]��'�ï�_����C��0���t%o>q5?�J#̢�L{�n�ZB�*q�Ϙ�-\q�@~7l:<-��Q�g���xx�?\�2,����]ާ�9�܋��3�	�_��S�Э/����Az����^A���
��k��G�U�mG<��ԭtK��3�i|�ꊠ/���%n~&\)��bD�!��_�3l����ѿ��7ѿ�7ӳ�>G���7����O�������Y�b��p�L�'��
z��|_d��)c!�$�,��:���=Ȍ	�C�$�pI�cHX��C�yp�d��/��:�~��)��;�Vu�����Ff��I�c3�S��5<��ǀCV9��v��N��ml����N�:��l�Hsr��Kemf&�X�{կ1;�Мic�u��:�3�L�������pa�T8�������M�/ak5ǐˉ4g�)}�i�PM�������\^������8+��C�9s`���X{V���M��-���P�5����x����t� y8ICٱ�j7ڈqꙦ^,	��F�N:l��F�{p��]�tX���#l�}���|�JY7\b���w�p��~�}��Std*ΛǾ����)��[q�P�ZoQU��=6϶��Qm;#��W�6w�!9��o�#0�k����|��Y�X��'8�ύ#p�:�I�|#����.d�T�z���=g}�:�~3,����?V���I�KQ�0� >ojxyr-�[ʃ�PX�;�me�`no�%(��ץې�����W5�V��#է�ث��++(|j�;�\.��ޠV,W�{�#��������$��Y���N�@�/�0�<p��[^��K�-y圌Ң̝R0�Ju��K�ǍY`�.�)�LyW�%1���~�80ww]�@G���<����}p�8tih~ׁ`;up����p�`f�.o�x, N y�7���+��ğ�s���2�6С����+`���F{�AH	��/Z6����V*˳!�u�3�L�ؔFs�c���~V~#�Ų�,�a<[oT!�C�� ��ʔ�H�J�o�e��sSps�mn���H��jv����`kV�j\�nB�oт7�C���BÁ��s�'9��Rp�G�HT����cI�����3D���s���?I���>K�������Kx�Ct�m���o�Bt���zW��]�[,(^��-^�޻�;��A习?$��.��U͇D{���x}�7�;y}�?�?�K�{��<}�?��^\5��2��-���d��C;]v8Qq��J�L��t:�#���1"�o`%zI�'�6���]y$��0�p�{8nt�SA�	���Ҭ2l�q���	Nײ1{�8k]&���+</�VfuzU�dV�Y���:u�F���a/C饑-���Y�/`�����i�tTwo�w#���S*�i[L@�f"6�v�g�~c0Il�$��deqo��id�a"�6��z��Z9jgh׸-�R����:{;����4���y��9(T>-���?]���[���b���|X�^�r�aK�
����z�q���Hy����Z�Az��z��5��_��1�g0������������H��r�3GG˕m�N�C�������u�{��a}I�^�_�v;~�	E+)-�-��U�<V����!���)ibO�8���1+��}!k��}�����[=�yo��By�_�kUve�K��u}��6)���v㇟�\��W�\WzѦZ4��"��9W�7�3j��pp��M�`�~��K��i!�����^	�)�u��|����,YkbĀ@;�&f���B>��ޛ}_Ԋ!b����G/��kU�h;�\1�kt��]�ߧ�׎�g�߇+U�rG{���rp��V�{Q��쿠��t���
�q�%ʰ�=��o�����j(I!o�zl�jG�]�|N�*�S�'�r�L�< p���}=�}�rQ�G��X�F+I�U	��O��<��C��I����/S1�N�U�w"i4����	ܛ�3|��Ȁc��9�I[L�Ue�=��I��,���o�����i�}1W�S&d^g3Joz���kSkn9����_#��y����1�w8s��F�eH�	c����[kY@��C@4zr�2���V8��*�ﶩ��T� 	�O�1��e4b�>���������<�����!��������S�~�3���<������=������n��2\�E<��FW�kc�A#m<
@�E2Y�w}��xWz��U��x�5w�o��m�~���?����L/�����!���תP����H''�,!�8�Tӌ�=V��Es]�V&Zi�9�s�� ��4r8�� '���T9r�3F��e����<��m�YѠ�	��|+oq\+��.��7]�+|Tzi8QN�"���=%dAݧ��{��18U���ϧd�~��z����M{j�F�l�Y�j��;�l�f��e�M�>���q;Sunx�l��uؓ���s��I���\��n�m�[����%�:��Knڐ����/�V5|�����>Z��e���ŧ]QM=�f?+��`P��7�՜�;�S>W�Xdg��"�"td�!Z���g0�ÞnX=�`����g?�J/�ҖW�vY,�.FK�s8u���p+ *�|AKJ�i�נ�]PR���/�X�� �i����
����
UJwG?R�eg���&��.b��ݷ�ZQ7�RJŽ���wҁ��t[�]�Loy�N1,mC5��ڂa:G%�BV �cx�29��:��H��D�̩sdo:���"MJX��9���'K��=9C0�(�9�����kK�|H��o��������kn�W�x}�?�?{�i��_|��x��:�ް[)�"
ގ��	jj
ջe��,!\_������uЦ��1�k��D�a7���@Q����0=��(Wq���`[��yC�X��z�6�#�G�1��Ҫ6R��qO�xkI�y^�j�k��uid��x~��Y�>]�|GP��&��vF�*7F?���f�1��4g��v��f�6�]�7� :��0�?F�`�2�z�L�L��p�0i��!�5�c��s8�G)�b}��z-�T}5�b�9��hۡ�({�z�-����������k������􇮧~�[�/�����>=q�詇�|���VZuK����%-���!F��A\l��t�
y��p��!����~D��|�2@��z��}���?�Qz~eE��N�/���DŢ�R�1@�Ɨf-��3y&��N)ZTc�����_Ƙ�G ��$oI#G�˟C.,L���Fa�廨vi��� ��𥝨����+���Z������r����vʛ��8��]��^�y���E�3������sFZ��ܴ�|����ش���iV��w��r�-�+�i����C�c���"�i��q�-ݦ\'m��]+�ç���H��,��|B�hdZ���z�T�JWo��rr�����帉b\�>�O��2?~飇F������>�X;8_,���ʶ�������|�-���_C�z�~z��W���=z�E��/�|�+��+[d}>D�P�B��`�/��=O۵k*��>�)���-LK��[���A	�K��.��ӆM�F����]�B��;�{c��g}��
'�͒���ho
��������Ȣy4��8��YEh|�_�Ƒw����3����4����_��!;*Jq(oc�(�:���g獨(�t�Z�\�p7a�>�쨿FW����·�_{�/�c���^u���`h{�F�p�]��;�B�s_���w~��p�Gt�bq�v�p@3(�ي�R7��E��e��6#u9�T�eJK�%�Y�&4�T��"�_3�<iɂ]� ӊ��p���g$�B�m�����l��%'�gޔ�5o~�f?�O�ydNL�_\i5]U]�*D �	?�i�/��L�4~��Yw���q4�V�>�.��Y'�IQg����4�9&m�vZ� "��'��lɎ�\ϰQ�방��(��B�4�M��%
ۑ5�S mW�K��Q�a֮Yx�]N�r'm ���	;%�,�9o�%鈧���!zqM���!��Zo�R��וH���2���]�hyiA�Y����w���=�������驇�w=� ���W��ޥ�su�.��α搜*��a��G}#$L�4��"ՙ�s���t�O�ɿ�o�m��?�W]�78�,ɯһ�#�[�k��E�X&+�0�l�` c=���!��ں���c�d)S��?O�lZ�`����\b���=31���s�m[vm{<v\�{��y5\��4�열�b�+Y�f��`�>�cᭇ����Б׸��$Xw���j�>����
ֳ�J���g��e�QI��*儯%�e�
<N0^��4W>����3j�X�gw+m��P��*�m�^�%]Ao����^��s�ي#�"�Rv��M\�ET}7�lH�%�E�zRf�d�G�[��<H(/���m7�)�bh~dM3�����J�̕ш���{x���������|8�O��p���P��kt�ڒ��&����_z�[衻�[o�B�2�1�y�{����.������������{+�hpD�t�wD�bB�z�m��+4*�Gcx�Ij��Q������A7<�}$�a˜�E7ӓȘ�.�4\�yJ���wW��.����-�0�&�I�1����{��7K@o�7|6�$��C#-l���˷���[^�P�5a�YY���c�9��g�j�D���(Rl�Ґ͝b��1Ht������;�%�FQx❼Q��[�>���q%�_8$�R^q�z�ï����'����n��hA��p�0b��.�w�ѣ�?H��o�����o�3?}��.�$O�3h���:�9+B��٦��Rd�Z�(��Wu�q6J����:3M'����Lk��V�ON�}�L��3��l����Օ����e`�����Oǻ;���(Bۂ����"9��H���q�-'�gz^Qy��o��l��;|u�O���J:��pƹ����]T+���iγnm���S��\\w�g��FSNCV���g�6�s���s�Ƣ��3L3�h;�;��I�]�M�)�c��Ўz(�ג�s��	�+W�gI�ee�sg�q��y�ߤ�m��kwV&�~�2�Ԫ󐚿�003��=�[�Ia��ĥ�������Cϒ^��1-�.��in~]�B��������_�
}�O�}���z�A��w�����tcW"_���)��;��AO}22�^�xR:I��#�ޫWio�����I_�ʷ���Ӵ��+��铽�~�����DvQ�N�/8+2�c�2����"����:�غb�X�Dٛ�8�-����6��zR�j�a�Ĉ���Z��i����n���v=a��g���Ƒ�u5`��]��+�]J�kp�@.�m��-/O������]A&�
/P�=��tv��������������6֞���ݲ-,��lG��g��s�|5�F�(��6dL*��nO�l��Yf��L��F�a�����O\'~ΠcE���۱����2��?_�Q�]����7�0Te\�i�j���3�Zs����zb��e�	>�p���~��`�N}
���Z�^���x�U:2�Y5�"�~^��F|.6�7������~��,q=��غ(Wh�h�e���Y}.�)����2�W�������C�{z�+n����7ѯ��1z�����Wn������!�����=�z����o��]������?���~�;��*]t�w>��xE;��ܸ�/i�b�<Nh��[J�3�0���ʣ��O�խ����Nkm-�ۓp��,t��!Y�+��oG���/�2����jN���;��q�k-��%��|�njj���'��.++`0敊j��D�[�����gT�f��yKp:���etϠX>0�r7������EE>F�y����!JFuI�k���+���G^O������=D��zk��18zw��2 |i[�%����x�5���]����ӋýԋE¹�Jc�5��|-���-sfΪp��	P�0�]Tʲaؔ%�r����avN�m+|�����a�L�:GY�0��an˪,�rW�$t��O�L��PR������e4~�D�`+
���?WPo�|v?��
�n=CcZs�V�:�Jo���e,m�Y+�'D-~H��+����hǍ����NiwN։}v�NC�{k�IPޛ�U9-��t�<�]����̡6�2&����p���P���{s>^���In�ꍿu�>J8o|
M��J���	����sDJ�J�b�<@�*j���z}0Ѥ�a}�GԮD�ۍ1-��뵋�֋���}\�Wo�B�_����'�}�����$=���������n�D{�=����Ѯ�xIJ��t.lp��N��e�.�C����ƻ�J�ǧ�DWWJ��`;t�Ƨ#��Ab�m��6Fgٞ��j��t�����|��Q~N]�z�<H�f�К�~�p���|��e��no,�0gSH��e����&9Rލ<_�׍(�Zu�Ӿ��ن��#��W��=ְ�<WW�������l�>���&	Z0�F���S�)ce�Dz��t��|V�-��i�M��p�O��Ѷ٬��5����z���t,��o@k>n�#t�xIC�;<�5:���Dh�$ɇ:�W?]���B��1���dNp��@떉���#�p���U�Z�B��m�{X�g���:^������ �d�1Ì�jpˉ3�i�akĳ �^O��!��4��9u�8�
��`BZ�t�9�K�K�S���/���!�����O>N�_�����+Wµ���������vl_�^�9��hI��wЗ��u����.�3�.��!W�I�����Z�_N-,��/�8]��Ryh��K٬"�yW�=��\�)O�\d��A�騹-�倈�¶]Sd����Z��x޺~\Β�ܟ��Y�J<5�yjp�H��K]���&��X(2G�E��(S�q�9�NQyA�ߜ�<���Z�y����N^|�s������(��e�5V�����vDt��-���ɻ_Ex��ԛ���s��d�0\2R<qwq�s ��Mi��Q�j�U���M�O��S��<K~�o��{�̣���ҿj��r�T]��Ԥ����y��^��p������ G�O�^N��vX�9���;'���i�J��b�u䜠o\��ө�=Y�1KIZW����Qoe����Z|�`ͣQ�2Ir���*�oԳ��k�2�І�}�c
�mW�JЌ��FB��vЈ#��71��n����9���4pG\��6�Y�;��fA3��1��Ò�7�&Xf0�]4�����3�g��K�F�&��W�&�u�1i@�4-!��!M���i���<��y�g���sOV?�ZL���'���v��>�����Q��i���7���{�'���>K��O�=�/�[^�jz�c�[ｗ��vZ�GC������z�m\z�����Қ�`w�ƫ:��t�m/�����t�5�����������u��	��٠Ĵ��)�B]�6�ԛ����ׂ�t�TO�ݶYք4l>] DD=C�anw��d��<e���@�(E7�w>@H��+���}˂�8�W�J�H-���*�rE���)�X����>�9�}�e[���b<�^?f��1��iyn�S�Ӳ;�|�ʭCSK]��A~öؘ���,z�8���_��A$7��V���J��(l�Nq?�����[M��I�H�:1�ʵ	Ǟ+�:Lir}� ����9���5�����c��蝜�{�JQ�c�f��Ţs���2�Lօ} B�K��5)��
ˣ%]=���ӝ7�@�x�~��7?A�z�a�����l��0\���`�CgB��9�����++����<A���g���cQ�M�:f��X��r6�������U���r��|��99BU����|[���U���U�քmH��Y9]��O�9O�� ���tn �jL�{óR�I���8�����gn)�� �C�+u�9	y���i�	YR,��GQ����xí�Z�!,�2y����]؄[,�V��!���ttH���j��w���z�1z���\��A�X����#������q$�:�ݞ���SYa��r�W�U��H���	�4���Vq������W����
*r�L�"�c�n���ߺ�<RZ)�Q*��s�ˬ���`��U~� q;}\a����8��y���!ƍ'�E*��|���lY(�3��(<J-g�Q��h=�z\I�F9��Ӓ"Ti�Z�$�u�/�YS��
�'��Fb�B��Z2j�*��#{o�I��a�f9lOᐧ��ifcVJCZ�c�	g/���&���Ϻ�5�.�����E�������4��7����)I=�uGU��ȁ��K��q�_(����X�u�}q�/w���]������̆1_�rA�<��]�g��<����z�-����G��G��{������Pǰy�\�s�&�'�@�a���EW�������e�1󁾃QN0w|��o��2Y�w��0G��H�x��	���h��օ�0�_q.��X)�%�<�Rji�/q�3h���]xk=�q����"N4�kY�n>��ͤ�@v\����mQQAr��x
�DhTc��YN�`-Ob�hl���Ƃ�k�������MD��֘��pز�����ekUiN�x֎}m����I\er=Ȍ�
Ω���>*�LǨ�$�u�/���?8a��X���bqs�6_L����W�.J���"��u"+�ƭ.���{�e�T�u���O�}�S����~YT�3캽@���R����EGo�~��w�����}�d��6DG�H}�Ej�C�����c(��8�׼�:8�#����̺������4�T�����<�	s��T�`�)i� eKD@kز]�"�Q)�r}�;%t����7ka[*Ex1��J��n�ZwӁ������� NL�1�c��KU8�BqP�{}hXq&�%f����$`�Hj�"m���cyys�|RM��p�Ń��5�I1 z���+��Sā3Z���������KgGGt��/����Iz��HO������F��p��j�/�\FOO���˰9���5���ʿ�Ш��|�Lo�u�#��]:��`�j�\}!��t�S]�ݍ�����SbD�R�SOS�NY��'�(�U�����.+7��\���V!*���"p�y���X�i��˵�k�� V&�º�$��JBc�^��Oa���K�~���yf�&�a��y�.Ҝ]�n+��KZ�4���
+'{ǣA4Q�$� -:�.��
d��=&qQ�p��3nO�A�_���X��<�<�\![�B��Xʝ�,�k����#�6���.�������|l�zJ!8Q�Ԭ38kU-BB�i� �W�)	��в�4�1<�l�RvE�Oa!d��7�UB~����]�#yS��X���Ͳ?<^}��S?�F�����?��g�;_M����=�<D���6�<���Z�	��:�H��pJ��[��^���?�o���t��Ɛup@��x}ˀg��"�zb�
���*�%m5c����p�q���PM�#���㠐�؁��p����:\�6��iʺ��@�{<87$zw(s���ӑ��jg"��	3�y�ҳ;:}���#pH��L�G�7v���ŕZ�%�YC�u\K��)�&�{k豪ܔ�cI�������}��Hd��U��K����vǆ�M����Hu�79��e�'q��<�(QD�B�o�y���}���[,x�_�R�ve#�z�ߨhG�<-�t�Pͽ1F��|��٨��-���(�����<'�����9�ɂ��F:�暈Kj���/�/�{UZ�,���f���j���/��gt���/�ᶓcI4������ܸ�(o|�+�������c��ݯ�[��7��?<��g8C�30�y!h�< >e�~��ǳ���:n��zL����ɔ�$)��x��]��Csުڬ���U|����F����0~��ty�Uo9o�.��xc���87�|�UKy����e����~�p�mڶX���g3a78�A;���v��4�L&�#��g�Y=|�A��Jʚ���ɏ��F�h�5�l�Z�Ӓ�_˰�]�vQ�Lbo0��l%��R�JF�m�G��Y˧�ă#��!-�-���+����_}�[�m=@w���\)�(	�A�`����J� �ӳ�5 �17\���#O?x��p˒
�]'�K�1
*_I�zT��$�]�V���P��KSk�9�âlъ=GP6�"1Ca"�[�+Z�q8�����P��
[��mԬ"1�]�\h�5�kU��;U�k�|��]0+�.�>��MA�tZ�E�Y��j��|#m�r �L�c�;��rp
��~e���r�]�����L�j2�A���k��!HS��y�ϘN��N4���h?�]t��a%�u^1��	;Sx��f =7psĚ�Ǚ�֦���Z|�@L~8U��lL�4VU�zp*M�7�3�1��J�Af�^�٢�Xg�s�mV����0�}�,L������ѕ��%�/z�t����}����~�n���ӣ��N���o~���Zo�x�9r0ș@��soA������.���ɖ�${):����D�f�MM��Ag����� �JZJ���E��A3�9_�V�q6I�ds���+oD�����[�e/��K6��jv6nۂ]ټ��(t�@1��0M�z����%�3|��Rl*S_���;�$����n'�<�6��ỘfI����Fڜv��c�����f.���c[T��:��/?���p0�T�����=�}����v&T�f1V�z�&�M���/�86hsS�=�+�N����"��~^�[ö�뜟��H9(̅�D��ɒ������|%%��Qg�t!��Y�����ҥ�z�5����g���t0|���1�x��b-CD�a�����#Z\]ҽ/��~��G���$������{��e��F����|%_��цN��?\�.I4th�������#r{��I�w��5-�L�P���ef�%�(��A3�_i'qa�
�W�_�c8�dZ�Y�,QC��''�d>��6��]0���^��V]~�o��sΉ���R�p��h��r�L���Dw�	<3_vҁ#3�8��3q�m-H�#+��
�L�E0j�8@Zv>���	BIr��3�_���k(�>/���r�޼Y����iܗ�\�>bQ��e�Z�Ե�Vч�-WL�p�,������Cz��W�o��{跞z��asr%�W
Ewm�1;�}j~P$�~���=l@ۑ�.���_=�ɶ��{���/<C���?l���힋� g�+Փ�������BJ���ǮT�T�Hi1�.��"�CI� �!��=ҁF��n���JM�n�9{�m�sSP�^�CplP�8�O5�>g KH;vx��s��g�E�79Kyٶ+L(��1sJ�l��c�5Z����|�4�N�i���oMLG֌K���W���8���NC#�nO�	;���H���o�)�c�76�kS8ˍ���c�>�Q�EZ�gp�����mH���x>V�:iJqM�+nTN�^�Ջ�\�i|0s�s�TG�%v�i1�(�I���ەl������V�]�\��������2{���џ|�O�|�����E�~�~z�C��׼�V�t�`xm.�	�aytv��@g��������gi��M����Y$œ�>��7�{"��\mR�t,����o���!�]k]J�IG!�c��L�=�]��1���&$�p/��\r`�D�4o5��:>-�sҗ���~�'���{�&K��@�#�{U}��8�� N A�$H�HJ<F3Ifc;f��cc��a�l���5[�O�i�ˮ����;�����JA$@T�}4����ˌ�8<��#"_滪(�^f��q�������pM�"j��h�c)lh�(tӆ��ztX:�r�R�<�fhXI���r���¡V�s�n�b �BG��E��E��ӿ�8p�V���}h|2�I��C�;4��*� �~�� ��d��eM[����T�ӍEY.���&�y�D'hA�5yw�d�E�2����dZ�:�\��u�)�M���V%�1xN#t��a:��6F��LI�ι91 p��h|/��λ����n����~�����1���^����~	���1H����:؅:}��)��n>�ފh4��C?���57�����=�+���X>rS�<���B��.p1�R��D���+�w��cODv*�#��G��������z���n��b�D�dW���M�_9#�����:����$�:�����|�5��[ʁ4�8�C�@(؂��ϠGji�� �2���#K�3��FтLyn����i�Gs@�� q��c�2��!Ocm�t��{��ݩ��6���/��������F���6�{��Y�
S���&jٿy�#�� iClB@Ư���svx)d4��^���?|�oFдTn"}/������"��i�&�`@R���F��@�M̈́UM�
��
*93a4TAB>����ac_c�KdQE� �������r�	E��s������a9�z� �/�&�WG:	]\�ď�� �%�+	S����a9��p����Dq��V�E�"�FC���CeC��!�9�?��y�/���8���e*_
�q
��A(��_7F7Ŭ��
��f)`�n���}vI�,n�h���W֭��H�1��㭶�]�����v��O�x�I��c����#w������u��v��/�FߩF`@��
��ÿ�����{�56�:Ơ�m��$ײ��B � �F�ٜQ�)�'�ĐNFԚ��D��8U�G����D�g��8�}��^��t
u!���b8ۤ'��p�@�K�Txg#�0�Y�t }��>aR��9��I���I���}�I)��e�ա[du���!�S?T�=T˴C�'�"���#s9d�py�DF՛s��Q�&�S� RZ�K���P�e=�&>嗴]����w-rS4	�>��:&E,�z]�)��=�h{��n��a����z������+��:�7�+��ݷ�m�]'��ï�����rt�ct��	�j�������� �ı��Nb`��9��8w~�ԙV�9�~�W��1�����*<Ӿ����DFQ�gy�� ��gCj$��a�7�,�{�c/�"��tL~h�F���pnh����}H����V*��|�{Y��!iH߸+F+�>E�k���84������K���:�H�ے��1\"@�Hv�,/	�ʔ@@V3rD!(���_�7��0I�������-�D�I�Dľ4��4a�Q��Q��`6�A��G�8w�>	�|�.���w���	�>u�����(ֶ�6֖�����;݂�H����E�	�p'���Z60U#��c��;���	T-&��-,�E([�	�r��y�{�̜���l��9r	�P�n:Ǟ�S,�s�ep��1Y�E���G��un�.�תyN�x�B�#��*��io�ē������H!/�V�����d��t�*i�<m��a}�ꓮT��/mj��
��P�����N���S1]�v�����A�ď��LX��A� ,>H�~��u�;��
Z6/����<��r9��C:�+�V5�(y��E�m����gr�'R�.gp�+J�#Է�r���A]L����������H�1��R���^�	�3��=.�����S�l�������s�<��c?��O�n�(��?���Q���0ҕM�/����������Z%g���q��A���'T���ڌ~������JAΈP�A��� ��.��.�<W_H_�F�#?�?ÖUѾu��8u���x��a$��Ie�f,9W����s�	�L�pD�K��@�S)�Y�ޑ�3$l.zar�2�\��)J��6�[u����Am[(���UIO\���C��,�����^��x�6/���|Р�X�������HU���Mg�e�k�^�q�7��PP���{���r��lJ�-jO��a4��	Pӣ������Z�}֩x�kw]J,���m�����.����믆G����������#Ƽ�w���j���8O:��V�`�,eK�CT���Q2�[���M��6��?�S8��;�F�ߘ��ݵg��Ҍ�S���D|�=FA�=c��1@�^�s�R�>B�2#d<��p�b�T�]�'Y��旯B�Il;�P������̀�"�:��&E�y0���{�}e��rh��!���H��e��5���p��j�Nޕ}��eV�[Us��˨���bW��P�L�$��g�OIW���/�Z�Li~�$�F ̪�Ҥ�	����#+4�/m�7�0�@�~S��a�`:k`��ښ��>v#���G��8u�l�Y�
�D#�Y�	V���`��8L�k��7�s7ne��eU��Y��7.�F
޿���/���O�
^m�L�o�Ș���`0g�Q�5��u�K�1拌<F���A��A�ӡ�b�B�Ks���2m?
3���(}޴����R� ��p�4�1�/�Ca�<�Ә����O���!�!O��E���-z }Hi%/9�Z���7?&B߫�΁��V�@��b��E��]UXVP�t�'��t&,4,�g�u(���􉓃\�yiK�[���|�Λ;I���}�]�a*��,!��A�R���4=���$�%3�hÏđ3���*�qξ��w�l��M���
g�����ф
��	U8��z&�������k�8�I�����х�e�K<�S��;�q`���qyS�� 9� �:؅P���� pâ ��Ъ"�XW��}3����u�.����n�k�ӤUr���V���6���\�~�e��g�=\�u�����尵=�����{��ut��4ce���Y�uSN�����=��̟�G%�F�	���'���D F�x�2���|�hM~>�Y@������;��+�Q�hBɣժ@�6͎g��f��R��ޏrR�z�D}\,XŒ֥�a��{2�Z�U���p^�6+C�0�}�,�0 �N�ȴ!�u&���"���@�S�4SnJ����ߥ��y�8h�^R*C��,
ݧ�ե[�t�R�n��8}%�c�Ѷ]�` ~�0���`֏�֫��α���NtҔ_�&�M��f���$��}�P�ڄ9e�
h�Cxg_�ߙu]ia!O�I1���7:,4	�u��� k��ȯ�<C(*��r�n Xq������'���X^X'm�grw����e��`�O��ó{{p������p��n��G�@/�S�N���^�h7q�����y����C�
�C=�}p:��C1F��ȗ�L�ﯼ��������z
�=v��Fސe
��`���CN�D��XYyFc�@�o�7C�r��(�y��� � �@�:�Z4w���ϯ���s�\���]��L�e`x��$�Ց����k���Yp�U��A~7�+ޗ��uo�����������K�=P �h���]A4��Hp��#q�+�$�RN3[1�"�H�T0�"x8�n0�$߶�oܢE�3�[	��	!��T�¢�jfF��	�W�<�ڸ�ڝ�xw�oÃ��
_��g��o��\~��V�0lӖ��L��������tKt�������U��*p.�߿x�{�u���g���1x��N+4L�l�ԠM>>l%��iǉ/�up�A
��8�1��cǿ7�Jғ�L/����s����u�4�z��*O �h�"y��̻5�B�*A�w�m��u�2�`���i2�b?KŖ�w�c��B�)�hF�P��a�#�~P�+��(�F�z᪘�B�*���羕�l�IX���g��ͫO�y�w�,qa@��4j���zTlv?��T�!I��L��%�.X��$C���'׎A��Z���{'����IP�`������+  �6��C���]��r�r�N��
�f�vrt|����Ѥb85��,�,bH��s*CXxL�}�bs�ɬJ�yr��J)�P�AY�͊�L��2	�;��Q��zX��EG#�S���j4�I����Z]��W��#o���m�Vjs<��:#c����Rc���hX��WG�[�#�]�*#�d�O���{�;�+��|���� ��8��iA:�u���ɪ�.��x��yStK�_A�����f��G����w��Bw��
�MO>Z}Cw�Ũ:L�xr����[����L:d��]��|��kW�2�)n��!�h��K�B�~���7
9�ye��0��<3@�?���IB�.����K��L��lc�����	yh.���.���nPv�@�[ �mg���+�29���#=+��r��f�SǢd��ɥ��ڵf7wmNl�&su!B;��r��K�<��iJ��*J��(R9_ai�b�����cS�l�5~�6~�$u�|�&��]T�u����M��'�>	_{�A��G��S'�`�6�ك�@������L���a��q�X�j�^FO���u�*�N�4�3o_&mho��.���o~�|�g��;���L�����mGk�A�%2:���: H��ć)�} �� ^����\��i���X��E�j�tPB�����[�[�P^�tuAYQ����a�d����l5G���fNPM����A���뙗EX�Љ������ǁZF� qr/�~�D1��in@� #:�"�b@
���y!E�~�� e�1�70kW(�ӢxE��&���l<niث[�<mo=��l��n��rߝ��{����NZ�m=�{И�q㡣"��$���B`	'��k� �)+�ߍ�Hp���P���^��vg���o�~�s���g��W_�Wۺ�&0o������F�
�#�Y�#d�C���xW�x�}�N���"mA҄@ʐ�@Y � �j��?o�3�碰>z���Ó} �Z�<������B���x�|EL�L�J��,��h��r�GR�+�����E�͋�%]��P��B�Ef´+��@ˡ��$B຾�idyY��4�~��l~D��К
�~��԰[���8@�I�C���$�㓎=/��$#�{���U��ޢ� �	93� �8eA���fғJ�\��ts�<�A�êI{=����^-�DCc�2'��.���8��[�Y�ߕ����x={
��'���hbv����l+<���q��B�4���iD�/6��Ӎ��FCP��)�Ӥ}��ea��h�tvS0��^���c*sIA���\�8 ����J���0��v���ϵZ:�C`�#.j�1C��/⒩F@x��k��G�(Ṯ0��R:]N�GZסw�~y����+Q��M�q#u^��]:]��~�z��7�U�U���Z2=�N3�h#'�/:V��*���^�ɻ ;i�`Н!V^��B��5�	��ɸ?C�Q��c�O�L��c1�a�|4�lps�{���"M��W�����T�l:�#���Ǐ����r�]p�98{�	���Y�fw���f�!����ۯ����=�����T�Hy�~g���e>�h�.���^8������g�ɷ^�w�1�j&m��ؑ��jTE/z]{0}�͆^����=%�A9GǾ���!:�H�}�݃!:LL����<$_m(���U�؃�!��ew�c2�U�?k,�k9�뭞��T���f�xb������~`7a�q>н|j9�(F�}Ή ���Y�J�<cy����_#Cu��_���m4A���ͯ�X�_kb#TШ�.�;3P���Q����k��_�n�嚫a2�j�VH�����tm�0&�lQ x�ЩK3��eT��o�۠1V�����\�6U�w�<����'?y��,�|��[�`<j�0��9����6��c��C	�	��Cr=C2(b��O┦H@����~.��d���V,���i�K]�G���J���պ�ɗ��0�6�|*���ޜ�>��r�.n�Sit��
�ih$ʨ�Э��9A���Pr�S�N>泊�i�����B� ,�?��O���Z�B��_��h9/�{��ѡ��4��g_� �^J�0���H�|����Uə����Ų]KK:�⢎w�	��I�T�Z#6c�,���CO��Fi�l�ϑR��eD,)2Jہ(?قK�� GUG��W�TP�z��}^,+B3F�]�d��cž�c�vq7���x��umsWc{�4��eZ�i<��R�Dok����$=����2:(w��f5ksr�4��B��q��n
�.daԿ�z�B���.�@���Y/K�oo(���D���b�Au��DO����H��ͩ��f�@���4�H�!u�U*��*]����IV�w�rd!]�fU8`y��DąO2?p�Ne�N�^�ҋVs��� qe�^�D�U0K[i馿s��2�wZ�o�\�]͜�΁�ʑ��{*d��!^�%@�)?���$Ǐ-���r{0�!��q����Ln>X���Ɠ�6��wf0ڝµ[G����o=�	��}w��'O�=��i�)�Ӱ� 0�VW��o�1�Tj��m��o*4ZpW?Vw܃����m�63x��s��g����	x��W��Y{#�ѣ�,�scd���YpTހ��V�i�̧,H��bJ�Z-�P��؟d�G�N�I� �9�!G\�rT.06u���cQ$��6�B��� B�IB�l3��L2 �p�sJJp�N���:�-�a��	jg��ܷ�k�Xe3�tx�E'����oJ;�b,�&��w�$7�@��9�#
.���Ϲ�u�-��r��`Ov.l�>w��,xӪe��war�"�~�Q�ݯ=����c7\[����ʹ�p�yKh�%���7���{mMD(l�*�oT���J��L��Q���M��n~����?�1|�̯��s�af�ql��ݲy����Ϊ����e!��D�s�;H����ri��\���$��z�h�OVq�(�;�����x��Q��F(Xb�K����,Zg��&��R�r<�.V�\3��ŔI^�fܷ��:DPĕ*1��tp�	���#W�a�8@��F��J#E1%"|)L�;��	�[�C>��r:�T�*쭭�b9*�>a}��l�Y�t��d�?��
��qs�z{@��A:�i<�p��� csu�0�Cd� ��ǣz`���ɷ>�ɘ0gD�.}��:��
M� ��5�1�p�D�5Oh]�r3�'�7�҆Q�ޠHt�I�C��W�(<1G� �Wd����+[��?7��XU䯫[�L�<�����^�%��������R��ċ1�}�#�+<W	�nou�AO�6�|�VF�4���,��U㼅�3_��TX��~У~c?ӹ��^���(��'�Gz��d�Γ��;��4N_��+~_ٽ��!8��e(~}d����-r�w�'�d?R���A��a�=��\�j��#�zr��!��Ftؐ����l�شo�Pջ��*�t�|-T*����!�>dF�-e��v�� �?O ыFH���v�E�=��6a�^N5���S��E8�����:��/~������O�Ȥ5fg3sw�+�l�������4� ��À�-7�k��}7�Ɛ��c�5�k����L�n���w��O�>����G/�/��O@o��Ƒ�y����Y�0i���"�g��O���>��a��C2c�Q����u�x��f�u7��kSZ�C��S�G
RLN�u!�L2����(�b5���tpK�P�v��εy��xV:�P����d#G_+�CXȤw�� ��Rr�����(�уTd�;eB$ �xѼ��-�AA�T�H���J�OA];�p���w�y����o{3P;3����[_�~��{��[n��G�9���Oc��A �� �h`|9����+o��7.�1�#=�j<���v/�Ϟ}~��Y����S���Z�bo���Ʃ��'�ZA�\�f����ʸ!U�	�vڐ�J�5�:�߬�=Y�0��C������&������t�	�9Sپ�~)1}!λ��hL��$.mv�i@$�x����1�VIz�qRE�N�/���"�m��2B�7�?h?Ԛ��ҧ������0��+�u�����\�2�˳��n�>�逤{��?�]m4w�qh9���(~9��:��(Xxc%�}�3ޚa��y�J�+o�=��7o��&vq��]K��a	���=��B��^���R��4��B��&�ϼ	,�t0�����l��<��ػ�IN���VX�����!�7\��%� �&iLj�.D�o7�~+���V~1��A����7�A���T�eX����%�*���!�0,3)�k?)gi�]�8ݼ�����`����R=�t�G1#�AD�����:/��ύ��@�Q��:�'���Hz��I99�Z���:�.�e� ������}��.�%eݧ���gt��p�@��mU[U�K���9��ļG24V�]�����%�pT�����iI�O�D���{�o�4�,ȉ����3�}���B�S��'�',�R�ZB��1l=��،7�P/X�n��"�(VAnf�G"��{o�L��j����ׁ̞L3�Asq
G���z��/	��.������h�^�{{n���z��S6O<8j�`__/����߱!������������|W0if�ʹ��'�����g�O���;�`g2���*�3j`�ۜj?�!He5F�
�����k�`)�ǹ�=F���\��	��C����q�x9,JRtܡܧB>ɚB��J�>�3]tCz{�-R��f�#Ѹ�&:��g�bw����'��yC�CF�)ɝ� x��מ#o����qWuCko���Үz俐��.X��b8�5 ����v��/�h�	�痄�!C���2J����7j/�8*�{<YDل{B���	
�v��Q\0qB�]䳖�&��A�+E�
v/^��W�L��[n�����sw�7^y�mmN[��
�r(!��:c�h���>��k�6W^#���۰Y��B+��ʛ��g���=�<�܋����۶w����MW[a��+2BB�v+CXy���MU���R_jI0.d*$,�%d8y�:���5�Ӊ�&�9C�,�s�m_�X�3��j1y�)#9�t�ؔ�J��+b�+�5�Q�^��B9٭ �Q��$*��4G=s$'+�wZ||D�.�Rv9����"\~��	�A�y��nsa���>�̷\X�6
��j�.|���G-:��;*�%h�tL��c�H��u�y|���a��M�:H|�W��U�DŇV-ߔE惤o
����2�2�@���7��"�p'��1�ޑ�����(�%��0J<|46�s��t�&��.��麆hW
�dr���yXVcE�Tι�-�zDZ������FR��!�g�������}Y�ou��(���z�1b�8�r:M����T�F˅�Z[�S�Lk����,�BГ$p2�i��r�,�C�!���ؚ+�`�箜�!+���B{+�@4,�M~�#��R�)�ž��^������މ;c	M8�0��0��˅u�7]a���Kð��E��Nӯ.z��e�+�kR�^��v'*���UCe���Q�{0�Y�yd<r��N���4���$&��A#��R#{�qd�s�<L��pÉc��>	�������?
W]v�z�г��g>m���_�����ྐ3���FS�d���q������������s/���Y��/��'^|ޫfPنQ���'0u;�m���`*�:��a���X�k�h�I�K��H"�Ge�Ln���oq �C{�G�q�`l&��hڿ
kB�M�X7�G��'T�^��aC�������J@}��Z���{��$g�"�[�-T��]�B�Z�3�UM�̍;Ԁ��AJ��C8�u�����.6}89��i�A�,�%Ջ%�$<���I	��BT�UT�#{�ı�_���k��Y+!8;wO2��}W�^�����m�O�7�\+4<���86i�Sf�T�Lכ��ڻ����� ��Cf6�t*�Q+�J����6�m�����ɳ��?y~x�9xy���dǎm���	���
)���1RG��/�l$"{w��0��v���6%��QsWO�c<!���'_�8���δ��d׉�Bu<�˵���.5�-�,-����� �"�Y:���U�x�!�%F�\�9��ZG�	>���,����0�GT�{߰�H�:�.���J���R|Z����;)/�����6�K�3uY���S�+�D���9�8��)���?�P��Y�g\\��!�C�0,�ɪ��;�� W`ࣂ���2��E��[��JW�/��aμ�:�.IY@����+	�.�2K��O��RӠ��hͩ6�(:ku�Y������xd�;�Wi`�R�`����3x��4��R�%�!��٨� �
lD�D�?6��nÆ�'T(`���!m�������BmI�F����,e�!K1O�39h:�%�}�Iɥ�a��E9X�l�N�(�;@,��L��H�<�:(сl~$�[F3���0����������B_�<�C���Va3����;��l$G��c jn���t��
�O�'�ӻ�f�~2�}��`�$̧A���ηfC4��n����B�Y�fovgS��j�����~����>��4��U��V�ߛ:#l�t�k���:Nk�\�ӹ�^n֬���n�AT������81�_����������/��g_�����t~��V�H��^noe�j4�����mu��ܕo�*ow�B���o���D�T#��T�{0i��������j>���9(��ȼ#v|���Dc�f3r ���y�h9 ��3�\Q�P�l0�A[�ª�7RT�(De�vuGY��TdQ�?�B��C�tŦ[;)��M(G�=�8���*�m<"M���.�+0c|'n��a�up��,ìl���0���u7�8�q�=��|
������X�Ns�XA�����W�
�4�du��0r�����#Zd�;״��?{��?��`�P9v���ͅ/jf��r��x�]�b*m���Q��L�2�a�}K�D@�1�r�@�G�<�q�<�h�W�c��mj��¨�L�)�WM~��j�*pV�w�k�
�uqdu����In�����!A����)f�5:� �w���X��3G��G�I�%~Ӆo�4P/}J)�(̢T�7Պ]_.ydTG�c^^P�(�9:\����c6��E���f9D�
�aT(O78ȸ��S�p��,~��u�X˥C67��!nO%Hھ�Qޣ|I�t������UzI*է=r�[$��x���rNi�����Z�m�<3�x�����h�鹨߁F1ƕb��^���>�G�����߻o�w��c�۶�	�V]N)����mM9��@ȌE_	L��R�p#����"��<2�˒�N�AC%)��TǘY���1H�	^G�b��J����8�.(�H0v�D����qG�������s�������H��
�Ju��Y�J�h�Jt�k���t|�qVIi��C�e^�Kx�9�%�eJ��tE�vNg���.�&�\W�8o)_�6.�L �Z�_}����s�]cC�.Z^������J��ӝ����un�!l�М�^�ߐ@�����4��u4d6�f��FL��5�;�l:��f�����:��g>�����k�����q�a䲩�J�5�n��E��r�"�7>�#�����{0#�Q�xL�x2O*�s�(�>���o����ݭ	�/���`���x}­��l*��r�7�U)A6p�е/?�эѺJ�=�ɾ@���"���L�`�c��.^j0~�3E�^g)s�W5��I�W:i\���!��P�d��hZ���|�y�q�p-�2�8��)cH���>��%ad�s�Y�
2�\G��F+�\G���؆���$lvY^u
l��Xn���!��1D�(��ٳ���G��T��ū-�o,�o�q���M
��ష7�z�"\�=���x#|���K���^~&��M��q����KX��t\d����M{�.��,�������()�4�E�kP����.����\�R5VH��#�S�ޯ�
X�y��
�������I` Y��K]�S�о�h��L*��<"m���F�1�H9��@�a�9��N$�]��#�M����OI��wo��}���(@����H-�~���i}'��}�m�5m/[laa��ܲT��J��AX��0���N�@g�������/���(��y��itQ�E�F��z�+U����ʡrB��!mw(��N�:O�l�W����0�~um^�R.���6)��NW9W��'H\0�MU|�CzA��(��2�!t��Y_���P��C�T����@�%��"vg�{�R3�{�����BpN�f)3q!;�*�-�����}�-$%�q`a����U�hF�*\����܉=��j����t�vvᦣ��[������MW����1�{;�������߀?��������N���FC��v���G��D�B9�[0d�+`Tnj������	S�О�?�-�;�F5�-�/�r2��t\ �hT\�xl���I�ڧ\� ���ς�#�&�}%�D@ǹ�e�A���et� 8�
K	؇�$t2�CFz��K�)�5O�)�>�[�8��}����!��}d��%�EX�]@��6��+��7�"��p y��RZW�/�M��Z��|� ah^�R X��<�6?��Fn�4�O�*���Uo��^p�TJ�5�z��"�0�1�?j��T�� ��4
�NoB���!^iX�=�J�"W�`��������.�v�qx�O���<xםp�\CbƯ�v����~<��Ak���E��BفG�	���7T�$U�p�3�6�,Q�@#l�kZ���.�ѭ1��Ƕ�U+ڴ���y�P��^pF����e�B��خq�MY�+D�Q���Gf�x���s�ي����s���������
�F�i�
���1�R�.@4���!7g�d�hUHZ9���5cw���4��6�yۍ��/i$�+�yy��q���*�к��S�
.�#�	��_-"mV���\���J�`��: ����s�%�G�$Dx
��o����E��
��9� ��u�%0m��=��^Z�~���&��Fj8Y��櫯�����7�n��#0��H�mNw�F�}|Y��BօHD��Ǥݯ��V���w",^{�E����o�>q���Ms^6&�%��:�X{:��o�׏�����i"�QP�A�r��Ҙ# C�kdP�`,���b��BBk�*�8�Y���:�b��yr������������ ��YS��!6�/�;_����,���r��W���i1:
�T�$���hxF�1�+�G�{��A�>�p&K�H���5��j�a��~�	�䐕�u��w����n�
[1�����D��	o��ýW�8�2��LY�|��"ע ��MAQVM�|��e� �%���s������	x�i�y�3kC�8>�F .IjJȋY�����#�p�R>J�$����@DhEs8�7�5�%(Qb`1�Q=�g̏r�kP},�S��B��o�V�
��\�sm�j@�5�ӆ�����[n�o��qx��;�ګN�V5��FB==>��N��n�o�����9��g���f5�F�ӡ1�W��F�}B���hh�L`��鄱�1���ؘ���j֥�ԛ�K��lقH}׿	��M?1��o� {j�D̦�#�VY�/���B
�A~�>��J탧g��6p�����[A����H��r���fXN��Cu��֕g.l�,�i"��w(䕄	��gI���I`�u��/�=�����嶘�C���C\%�.Z�j��Db���Y�^�gÔ�v�K!W��NRC�ޯ��m���@=���\Qds}�ы[�%�e7@m0كa�$/Tg��������e4ك1��8�xB�[y���vk�zk��f��G?��{\q��t�T�����VXsyn���It�(s���MT{#��q�j{m�*ȇ(�u�I�~�ԉ6�k�:n���(fmu��`�\��+ 컸������!��)I�rX�ۃ	��O*+���`'��l�����P�0�C:��ݘ>���-�a��ܡ����K�kQZj�6 �%V��.;Zn�-2H5��k@�FV������¢qPգ��8<:p69�W�Oi.$<�S�t.�#!�Ą�e���ě.n��͢
�Vc���E�ü7^�0�x�e�L�.�\�����5<x�u�O���w�uW�t^-���ح��Pib� �m/D�<cW���i�mc���)筣�i/�2�1}����Ե
�����w۞T0�B=�TҜ3��[|��Zs�|n�^�*.VH���2b�B��(0XdB�17OrB�GF���F�w�$���%1�:l�qF���UA���U^6	%jDH��z�8�Ě���C����5OrB��Ѣ�$H�p.�^:G8c�Hgb��/���d!����9 >�h}8����M��xׅ�\�R�\|��u��R�	z��D�Qf��.��C�*y�	�>J���n�P:Ѵ�2�S1$!�TʢM�2�Cj���!�Ul��C�ꤿ:K9b�%�JR��`��'�L"��WŸ���<��{�D2���2�2��~�^��1>�_�Wd�]�PEY��N��t��n��D������f�����+����mk{O���ҡe����T5�:1���/��������_s�$�����E�H�HcE�
h�y�@�*&+�^�ԭ��q�Gbz�����e{*>X��^�كT�����p� /e������b�o�o�N��z�\$�W��𸑟�<��7��<Z�6$��g����7}��E��{!JzǊ�C��\A�a���0��r�y:�z�^A[u��H�Y����a+����1`��,�ҹ:��.k҅��_� &~�H���<M�s���b;�W4�M��v����~�Gq�Wb���
f�8~��y����u����]���=�%������SG`b�-�]�m��43�C{���?�@㢷u�s�|9ә+Y�7;0�Y]�1����W� v�-:z������ʉc������6�5�ސ����*����x̛ #Є���z����@���~��}���`b2a2��Z�a�c�DE�����5M�l���y�M���`)�a,7B��� �0ʵ��]7i����Jd�Y!���u�i����PhࣻV+0��D��\�������KX��+�W(Nj�p�X~V�#zu|�LHLX�ns�@�8��(6B�\b]l��Nʹ��/��Q���n��醖���*㞫�u��Td�D"$( ��!�S��2��xfk+��&�V`i��ۃ�ϝ�Ǐ��5"�Y��1;ߨ�=�<�
C��dۊ+N��� �o5o�o�+7����3�	hc�@����7�З3��!�
�6s���Ʀ���"	f#tQō.*��Q	�%�OޛaJ+�d�!!�Í[>F�R6�E�b��ky�����c�)%��a�����DAU H&�\*�	�`��P��E�|:Fs�tX]ķ���w�3]��+G�O?���'Uj3�E���\_��g��<�Y�9�F���ʤ��r
����9�O�e0�H�A�T\5|X�;i�<�%!�I�%ካm�R�N).�UN�n���Q���o9O)����W�Ղ(�����U�n6��	��1Geַf
f��c��>�U��o�������O�9}9(�Bl��{`)��m�:�J�����
����o�}��s/�M�=b�;U0mu�%"\uo�:ge�{V���D'c��Ѱ�͢��,2��
�r��u���A�>�:�}����]A���!,����]�{� 2"w\{����'Py1�\J�x�&ǐr=����&9���
��mX��<.I#a͐�aJz����Pʫ�~S
���؇E�󌙕�D]���������C ��;M�ئ@n�-��P��K��{��"�����(C�\��s�C"v�7R6��fUD�t垘`�������	עX/fF�v?F��L���o�y'|��O}��p�5W���`����<n����:G�^���P-�]U���|ײ�*���^�&[F����]8w�"�:y&Uժ�z
Y�����q��~kcL�l����<�F�Ud?/L	��q���iߥÐ�!�L7�>(�D.�$Ӓ��F�� #�R�]���Y��r_�癃K���}0������ ]?�v�{�m5�VY�P�V4����!ᥢ��S�L��?TcԜ���� �k<L!�e\a�wJ���
����z�h��Եe�v��0`s��N��>q�u��'�/?t?�z�G���x��kpK:[��mFa?��S/�"�k��?�<�;dKJ*��18�����[�^|�m��_����<���k���o�]#�1�,�gs6���@2�F0�����_�Z�*~Ѱ�|4{�uhvF���F�He�� sߋ3^{< �L�S|lǱⳠ�/�͸)�q��'�J�K�e��j-?��g�2<���ul�d=p�s����8K�B�!�_��7�h`]���D-��'$XvY9]7Ҡ܉`�[됽æ?��9W\��'�S!��O�]x{�znF7���̅�Ń8.�}2�Bb�G~ȏ���J��y��_�+�|a�8��6U-��R��@�'r���W�+ۦ`��s_�T/�RB#J.8u���ۣ��aD!��#N\��+��x�y�C������P4�6A%�"�4E��t׈~#�Ὗ�� ��M�#{��qu3{?�h�}��{P�:�U�>}�M��4|����ړ���tm<s?�Y�mt�)^��=.�?��-W�>x�G��2���j!ea@žt���(=-�`�y�&c��Q&#��x�]@�O	YF���<�T�j��U���q
���˼"8�t�C\��~���zl��ɦ�.!2E��Q��5$��?M
�S׽Q��*Vݩ�S��@��7�D�7� _��K��b��Q���AB��SFW8�])O�vg� ��;�RL�ƨ���#���!��������	:�w��M�Ӯ>ϭ�b�y��k�7xs���/}�s�� ί�3�=���A#9��g�=��<�A�!
�m�����h�G�y�л����ڂ�~�������?u�z�0^�����2�b�_!{0q-��l�+�W�8�Mc���#�i��3�i=��.N���_��ξ?��Y8�;����1\}b�^�b콝��r�իv�(��<LM�w��{�|�Z���Z���}a��]ރ�`(��m_�+��Bޱ}��tE�xar��3�y�|��4�6Vz�g}dUzMl�<4DoD�9�����a-�(��n���z��$����9���\X��%V�v���9��3h���!��%Q�}�"�Ef�B�8_��aC����즛:r�	�%�t�e
�������7݅[/?	���g����p���dd�G66vZFm�zU�
�Z�&����x�p���#Zx�6�2|�����&�Fm���׽YϽ�2��w���x��w��z;�ؿ�ށ���ྛ?ͬq�
Y�i3<��L����vw�鑶��Tt�����B�%���
��>B���)����3�����o���->����&ҬHd���s���s`ӧ�r�Ūʍ��.
G�����P��c�+ �ɜ8i�����, ��t�M��`:%��D�Y��ᵎW�̘�.0�T�HT))�AJ5���[���<����h}���Ï����G�8$�|L��OX��Δ���曬���x�AubB�s�W�Q�2�&�~�/�už��"��mu"�nZ�]lrc5k@>g\�P�i;y�nHi��"eQ��S��@�Lt����b�..bJot�G�9%dW�ޓ�+��*��V�o`�9G^��o���u�ܸ�N�~�zQ���]���6��M��=�?�q���Sp|2��5��GcRKHm[��Kx&�@���1m����.;y޾0�^Q��	��s�s�R��Hӆ|3���(�#����E�%�+��-6��n-�#��\]��D�\A�q��89z�t���?��(���a�ti�Hk�����n��b�(D?��sf�|Q�K��*�$��9D��C��]�s]I�F����n܀�C���Cú�D28��IJ�9QM�ڃ�+%2CCǐ&�X k�?��d�
��K��o? ����8�
�=��J�WB@nOK�'�럒AF)^��}�+:�T�~�����|�.�=$����b��U�^I�)���u�B��^O�L����6��H��)�߁�p������k���>�\q�z�^����[���z�	eq�����vF"5�hf��V�⩌a�,�=$�f1�x57�0�����������������y^Q[0�g��[�f;p����g%6B�)��vF�P�Í`�p׭�ц=<�֭�B@X����1Iy
�@(|� ����z�7RF��B�D�cs��)�C`<�H�C��������S���>�Ǫx�㡨v��(�p�����3S�TߴtN�K��h���8`�DQ�eGJ{^
 �/������ꁃl�>ez�!|P �@$���3	IZ�^Kr�4Y��G/3N��>��MxJ�-v4�G��^yR�j8چ=tם���G�>r�2��$P�œQı�z���g� �G�6��JO,�z�p
�򂲛��ȸ��K�d�^� �z�u��3O�_>���7��V8���s��mG�\֌a��i�4�%�TGF��F	�5��u�(��V�V�U��p��q �o�F	=M����4�[~J(,�j9�d
����^��x}���q �ll*b'��u���7K��5����?�pe�!,	\ 矩���W>5�/Q��ن���	?n*�	�4YfS#�"�E��Bfb�Q�]��K�,2nrU�
���p����U��9����ݻ�h9%�m`�$��.e��[cQU���NY��x�8�2,���C�P٪Do`�yr����D�"	�
�XcUf�	��0b&�5��G��̉�c+pH0ɢQ�9z����h|�5\֞p��I�W�ڝ��#��뮇G������-W��PSw�f�l��i�U+�;画Po;�zI�xS`�Z�k:���WfS��W�0�.��6�B���e�T('�밮�!�JQV��j\H�
�M�����']/1�
1)(���p9fښ+V���Z��z��"�#A2\�ƽ�o����Q�$��tҟL�I�2��<Kz�E���[�0�O����H����X�:~K�Q��>��n�!��b�u��]�������spya���1nWV��`������uz�����9ºB�5%F��&���6����5�����.���l7���j:�+�&��/< ���}���o���P��3�L3
y��*Q�*�����;�=݃U#ק#4��Xl�Ej�������S/���œ�7O��8w�m�\�1일��wbr&��5k�Z���x�M�p=�3���sA�##�tM���i`^/ɔ\�]�U����Gr�Ҝx���	�^Y�.��X�x*�(��T�Q��t�����!�>4c�k^�@JĂ.��x�{�m� �fL4ڤq��y��iH�v �|���p�!��[]*H>:�h�\<;+3�,�4Q|��nH�4�%���v�v3���.�q�U�Ͽ��ޣ��-����g�J�!�	&��Sk���k��7�K.��o
�P��L�P2�暺�9��gΜ�����ݧ�������C��Տ�B=1��3F-�7F&���p�0���
��)���Ň��)��G��
W�v��4��r�w34�\�<_g�̈]t.A��X�\r��
�ý�8�0%A���Y���M�2D�7�u"'����pa5��7M?P�*m��4Q@$g�(�(�Q�>p�DXO� BYM+C@�����;yŐ���Ei��J������;����;��Ƙ|��{t�Od�Sa�ۺ�h�)���a��!Y��8�C�]��ʅ�s >�ˉ袕�%Q� �l� �('�H��=���e�� �H����8��y�,l��w�R���r���T]e����W#�k���ģ;;p�'��_�|���k���V�1:�]0ޙ����	xY]�\�2��_�WX�P{�f�i��Mx���`|�X���ڜ���D�a-�H�+.�֭&��sN�U�>	�Fv,�D�D��l�+U$ϋ��6tes�������� m �Jc��-�����U@�s����k��cpm�@.픴�0��y�����B�.�(���ɋ��$0pY^>��a�y�o�YZ�`=����!t�>�t�p�W Y�]���aݰ�S�w�/['��tۮx{�R�~]�o]��\��u�+Sm��\������q�W1�҄5�5�s��s}������������M�½w�#Z�Z��O�6!���9O�M���+�h��Z��{���u�Ad`�c�G#h����9��3���{�,|����̹xO���c6����82�
No�qS�nuw����j��֧*?>��(��^��Ke���N�N�̙�7~���l�ݬ0��z�P7r���Iq�QR5���b{0}ͻh�<<�,zސ���<C2��E!�(��utu�7t�B��\��:�8L�S��8e�CX�|P��+����P�t��$C1ް�B^m���q�(��B���=�?���õW��'�����p��
�������=�ֹ{{IUY���吥����T���o��I������2���
'��д��n������d�\�N�?�6��cc b17��#�\�]�~�;_y�z�!ѝ0[l ܂��������F���"XT��#�Ct�z�p#��]rܽ�0��ݐ�+��7�G�yͫ�0�웦��@t5��DK�f)F<'�7ˬhm���@�ӎ�z ?]�UP�U w���@H}.^4��ʅ�t��9���^�.Y���/}�|�+�FY��QT!��<g�Y��kn��e��^��!m�R�\��4iwEڏ& �n~�0�'�o��zl��F�po/68�~����~�7�qqr^�}�Y�%K�d5B��S��{>1_B��H&%Ċ�A�Ef/�Q�3 sΉ2�'���H���Sq�܍�?�k��	��5D
7פ�Sy��]��+�+��n���©#ǠjZ��x�h����V_2�S��S�����AڤSѨ"TN7��G;��Qei�O�yε���T��8�*�5�7Ѥ"	�k!y�sy"7�
m�@�\\jtxfL��z���M���_�Ӧ�>_��CُvZ(��$����P�'ldt����q,�:��wB:*�J��o����e���cjK]�=�!M�,J�t9��>4&��0��}V�Lڑ�>�a2�P݇�"�@�\*�i�@��>F�Q�S�}�%�A��iN�L��w�P|i3Q|�]�ht����A��y�Mr�e��J���rJ~��DL����D�x�օp�W�����{�װkw����V.?RW�����7���k_�#[#��N;�V`��������浫�&�C�x7F.7���bxU���V3��K����'�7�|�~�x��b�̶��X��P`|�7��Qc6t������n쯺s9Gޏ�>Ķi�������54^>e�s]��UW���9��p>�r)���H�NS�$v��.h(�
�4"�'D���[x6's�"��%��
���ʚ���eY�D�7^�r0����(W�τ�P~<�[�����V�v�vK�}�A�s�ec*����i����s�#M��x
��D� �F��ݍ�\w�q�\vq�ǯ}��o}�ZV9۳��SM<�d���������o�˷L޺���H�R�fV�]<㎭`�߽?}�y�/?�9���/�K�w��1��:�#���q�e���q6��!c���UI�y�Ԥ�נ�`XP0�.ô[P��i�L��vMP��;wIN�b:0U��(3/C�f�bJ�������P(@F�hj'Xũ������\��#�]��+�(_1���.0Jlj:��9�,_�Ź�:�3�3���%�q�a^,����9j{���!L5.�x�59�A`!xRE�AW���q͂��0-W�K]$�\��74U�i��S�g�%�{�p���.���ya�<���G��t�:ց+���@��l��R���9��n%i�|q/֛R����ʵ��)[�����Ky���$3�d�ha{Ⱦ e��ߩ�$��;^ɢ�dd�����h�a���)	�l!0#�G��.@z�J�jh�]ψ��Y\���rZT�>�ہ��G����o�n��T��8�Ǖ�F��urB���ݘ�5DgԤ=�x#��3��~��	.&���&ޣ�~������FǎZ���J�ǡ�C�-��,�<�=��7|�0'����ېW�x��ٸ��Kn���Cб}δ_7 ��Yf�f�H�)�zo	|��X��Y�9�)r�I�M��Ћ�������}�����&��aqNV>?|'�r^�ԛ�<�8 .��M�����Z�ʰ.A;A��>����c�T.�e/3�6}t�>zQW���m�D�J����௜��X^�K�7���N��n�x��$bqe���{�́v���=@P�kt���O�[n(R<Jyϋ3?+���� &�Y�(�����>�/��KZ�닲<~�_Q�Ȯ^0[+��B[�Y���ש1�o�ÿ�/�w�M��M!�� Uи�����ÇT�����r{u�ȍ葿>��l:���������?{~���f�?�NZ���I5�(krR�C��p���k�ہ��I�/����=�"}EecXbnq���D��X="���3�U<�� ҂L��P�G�i,%B�Y#��5�*��� �o8t�xn�a��8o]J�j<kOQ~�8��`$dޑ�E�O�e��76Cmr}���QC낵p؎����Kr*q�<T�9W����1$7��(�Yd��4A�h#N:���� ��Y�9��o|ъP�j{r�< ��o���!���&R�]t�+:X|����c*��=�5r��1�Pn�����}�-��_>��s��W_��Z�EO*���G;.�<n��a����V��u��§Y.�,
�R@w��Q�c�ML��	-�T��B�C��~k<��Nא�L#�G�"�9�R4R	'H
�!nl��m�"���.>A��rQ�(�兾?��i,;��Ê��ޛ7|�i��'�(3fQ��dA��������r�8�%���&t��\�}�jF��;�3�rPFI�� �t���M�b�Q���.��bæ�A�X�W��0�+ݕ��TE�Hs��b-��.Tt�Gڸ�x.uu�Ǣp��8�Knal��;E���#_�?�*/xY�l�󹪚����ǆ�����Z��3Fr��}N�IXf���s~pN�iD���N�� �iٚ���<\�r��<�_Q�Jxa�$���B�IE}ȧӤ<�mxw��m����?�S�^�s��a���Y{.��Ǐ�#w����gᡏ���oY]��{κIV�C��I7�ż����^`��c*�t�@oGϻa�L��+�x�o~�������wሹz��J�szq�.��.�F���,>At�|��)�g��s�vB��#��A�)�9*'�4(D�Lx"w5��OG$tv5�{�l���>:��p^��s�l�P�ӄg"|��l	��ߛ�\?���e<pTv�%S�WVp^2ޏ1���3�|��~�T�����e�l�r`� ��¤~�������i��O��I<M�I=��%���P�$��kN�!�5l���L^2�y�iH��8��14N=r*���Ci� �r�C)���/����V|z����VR�����i�
��9�5V=V�ҷ��ň*ۍ:�-�,�S)%�h`��`�ߏ���ٛ��6�����_��ǝq�$x7�aG8��;��dl��=&��=+��BZ}�����;p��W�~�K��3g��7ނsՖݙ��6����hx��,���c@ceuk���XI_Yo�*z�Fa#���4����a�i�^��B�w���Uξ~�%���ȁ��\��f�O���x�:BQ7�s�P���Ԙk��d蝣�t���	:�}��;7���h�>����Y/��a�X��������h�1��deJZ�.���`E�\J0D��2�]j+�9�����u~B��A����l�}"����=p����6��=Ƕ��e���Y?[`����/�6�M�8�7�+Z�fR�t���*[�{q/��&���௞�|�_�+�؁	T[�(�=m����w�"�	��*d~C�
�N�#�hh�cJA)�m��'zmlcaj�����O5:� o�`+�L4^� ���@�Z�a���D��p��Z%�>���=�$��:D���a{����B\=&ʂ�/�B�2�g�BCݟS�xE<`rzu{�gs��S�T
�T�'�h��t�cK�2�������2:�*��qY�6���OrxWuW�Sdz�Sw�,�;.n��Ƥ���e�6V�T�~�@�+� ��MA��1^5F��$"�D Ou�� �?d�d�}+O�u��y���#a�z��K~�C��Sn��\ɘ�+�r:��2~C�e;��kp~��G��g����7�xF���i*a!�Bl��B���%6�;�=k��c'�ӷ�
���N����GO��[�ֺ�Fc0:Lc��ړr6W����E�.�+�Ѕ��)��v���]�b� �]7�ʹ���{���;x�6'0��?|�*Gؓ���IT��|+<�Y�(��>��$�;ݜ�⒫�CN�I��%:�๲:ؔ����|3ns%�8��������ܤ�| ?GB�/F�-�;p���Lʠx I��	i�h�A'��a>�C�|�k��޴P���ߩ~��a%����5�Qi4�C�ij9ǀ7Cu���e�_��\;�e)��Ø��W��I���J��>� W��Y�%e�\�j����w�m�����*S�;J��Ӈ�����qd&4���c]@&>S��d����7{&���?u��O}FF����QF�P�Zk����:�LNh�W剟�1���H3��w���߀�~�2|�g�G/?ﴑ��U�  ��IDAT�.��-vFzj�Y<����ūN00Y�q��>F��ec�
5��,��4�Ul#��JE��iwԳT��~��c�Ѵ�él�YT �"�'���<<ު$�D(#��8Ta߯�#��dA%%7��)�rÓ��R�n=�,��U!���<�%w��O�8 �
/�ְ�&AC:���+TT��>)�끃4t.=Dx�"�I�#7{DR��Or���2֤ĈX<Zk�Y�8��^s�e�c[�࠸�./D���j�kB� !J�񃲡������چ�>�������g����s���0n���\�R[��l�kQ�I��ܩ6��$��ĸb�}�BV��ډ��JǴ*ė�fZT�:U�<�?y����
�=#N�@����B
 JD�BW�07FHR�IƉQ��\ }��i����A�A7�`�	�v��kT�X0�.�Y�x���╫ ��9�R�	u�=�)��L%#ۏ^�V��@e����������<�n��e_�e)�s�"��m�(��Q�]�3��P����u�8#��:�]H7r�
T���)S�� ����؎Z�Z�,A0�� P~H������i�Y/�Y��QZ�
;���ag-rQ>���Pc$4�ɕ;Y��(�{�\�"ܕl�k��N��8��ɑ�XX�j��%yx9��c��|�!>xoF���A����x�0��)��.\wd��F��'��9}
��F�����]�3'��U+^��$�u��%#�Z}ǻ[�D�\yiNյ�;�=x���{����~g�}�Ǐ��{1��]����GѮ%M���^�@�t%���Qފ�O�(߸�%d1�C+��D�Y��עƇ9��q�`/�nZ�q4Vp�����	�UA!�@J� �ڮ,�B���	P���M�(k�b�W�>9�D�5��~�+F����x1(6E�x�{�
�Lt@u�>y�F��,�'t�7L�yW�t�U�����~i��Ⴗ���A�z�j�E3�G�M�(�7'#��='��DdMn%�!tl9�.]���<�]�yF�<kV	���N���w7�	)�:�.��5t���b|�5���?�x�r�-�\	��s��q@�����m��|J'��T���p�he�7v4���~	���_z^����m��O���EF#�C�`�������q��`&#�U�<aX+��w�jcG��7*���	g׈q����A������	��F]��C	V#���Mtj��oB�A���@���{0��K�[w�"	�G�*Ltg�z�*v�`�\N��ig@���Yu� փ�o�SVM��C׌��ZXʀ���=�>��V�B&�*��pWk�(���4���rBD��H��9�:"{�1O����]���XY&�[��n�g4���U��i 'ƨ���Q��Mf\3�%�3x����}�o������ͣ'`v���?�U_�j�a֦�ʺv�./5��5�P�uJN/�s$>vUE!A� �F�~�run��h�o�{�Z\�ѻ�4'�5'F�y� ~�Qi��Tq�t�!�t��/��Q!h���U7u�z8j:x�o�z9:���B�e��	q�pZ1:A�:�N�?�w$�HN_9����Tv��}i�R��^9P�* [���T��0[p�q����9"?_F�8t�F9����*��x�� |�t�.W.�3���¤��+�xnؘ���-d֎4A�r���N9��شǒ�
r�#�E�򕝌��,5!	�zy����QQu�<�S�X4�e�s'�6l�@h����Â��^����>�Ud�̕�5��#���+���v��p����d��-�nu�ٞ+�1vWڦ��򮌣�e?d�q&Z�ƕ3R��H���N8r����55��9g^|��O�w��vq��[0;�m����s^��m�`���=u2�K�Y��>�Ҷc��ǹ�5( ��ؠ�nj�|�r�r��2��F�����a��h�S�t}`�rEim��o���q���M5��@��8"��X$�@���X��:�j��/���u�U���Q]Gg~�yS%HY�ԁrMT�7
yH�G��g2^Q��$�N�|��kuɌ��i^�>WR~@��x&��2�d@.�M�<D��y��9�8��|L�,V�{�����6
��;Jd��%�	��:�I���N�]�=�B�}�\.��nJtX�k�v�^��`�q���E����9K�|���"�OgSx�����?���p���М8�5i˜AՖ_���vF!W�Z��
�#gM�c^k&��+U���;/��:�O�����n�ľH,X_-+�ky��rY��츧s3�;h��+�fذ�r���lvթ���1=��-����S��C��B'~]擊�v"tM����<��5Z�2��/��{z�0\�$��AV�U��H��:P��;p���JK�����s����"�tU�؈9����I�l=H�'��p5�	�9�e�j`4n������;����,4��e5)"J,����B`�A�`+u����1�q�ix����߽���
��bdU�V@�4����U�X�,NV����@_�J!�&���q���Tw�lV;�Ea�9�m���͛$��gJ���ÜZ����4=i�R	��2
�7���\���ĉ��Ō@�B�ox�"�v�!�*�@.z�l���7흛�����;��	�G��Wc17G�&3:N0$�����"R��Ho�C�����2	���*Hǲ�ģ��+D�Y��dYN�;�j����a���"a��J~bM.�.�X�ذF7�(_���s�J�⴬U�I�X���w�����՜�w"���ٱ=��m��4%�ȓ.~�~ȍ�d���w�-��-����P�Pp�NA�� //��l�;q1] o�,�aot�ą����v�} ]7�JI�pN�5^�j�f6�fzpaNLg��kN÷�� <|�]p�5W��xjV��w;5T�X]���Q�Y��t��PkBk}��z�����R�kFcO��.�d��XW���o���5���g�dGv&��z﵃�hx�0 �z-E�K��g�P0��~(�O�~�B�C��vA)���rw�$wH���!ޛn��a�~��n��yιyoݪW��k�Я��Ms��'O~������p��Q�;��J�`m�_z��A�Ab�H�z7���[�n����V���\Z��f#ezd�K-��Gj3�������u�E�G��hE�$�"����9:K�^X��Ɏ�f������D]1Z�A�;M����{�f���g4!RV����SMA�P���~Q���2C/ꂮia	���QE2&K�.������}�N�oꉱL�����M��5���r\ۊ�+6�"ysk���#�+TG0وo��3���+믌K	��QL�`�eҘ,&��g���,�~An��G��M�4F��)���� �t�}G���W�b�X���f"��r^�Ӣ��摍�΃SE�$=�;)V���{8�a�{�y�N����b�²C��vC�do�����^���]�W'x�E?wnv��)���>�Ȇ=��✻]����ED7Y���o���x�6	�Zr> �2��g��R��mR�}�Xv�߁@hud��9/h)
p,����+&b8�g�x�-!y����F��E��HU�+���9�O_z6DvmP�����������2z����|3�A}�5�D�i��8����sH���#ـ4.I���\^@_](�q�K熖w��v:�����`Z�,`뷀"�ꭥ��,�$�&��|Nݵa���r�9��*��I�"_����G^:�[��<
z�6cRU�{�RQ�%2iS�(�Yo�[Y[�Y��������_��a�����z#H���F���8a���D�6JI�d�P�6����tꌣSd	�K��(˧���&�C�}8��h���{A�oI �sQ�ꊲ�f 9"Cb~֪vC�6�hn��~*%&��\7�s����D��� ܗC�Z��\�=̪t��xCVl%}Ntٲ��6�;�3�F� �1�k1FRG|��4/��'^�qSr�Ό��NӇeR"	|Y��'�)~�ߥj�����Pf��9�����;k�{�n�`�Pߏ#��AK]����)�#��*_.C7ālM�J~Qt<Q��p[rb	ur���K�/K�7�
����M�0�1'���%�����
����InNL�^BZ��olGR�J�8�^�?z"UɚxA�?�/�ΗL�{6��חD.o�^Ak�G԰`WO�A��ht��SL�M�kT����/�s%��Z\u��8eמF�¸���6�z�N�V�"|�6�t�XG2��q�:\�6荰����{�}7�G��w?|O�9x� ~��8��x�L}��:Ƙ����krQ�	�o� ��%��N�{�E��w!�e�d�e�c�kg���>�NN���>�,o�N�U6	4n@���it_�~N���
��u9�n09N�N�LJ��Y�� �k��A��wRߑ�,��AY�!�g�5��(x�~cTz#;��@���A.̌��t�S����>%a��F}���7��NwQ��(SⳜ�;�1��3
CE��(��*���4B&H�+���cR��H	D>�j-eav��_G������F ��ųRt��\�v�A��J,eB�9��Y�z�s=[ڶ��oI62$�R5ƫ�����G��͗��<n�=��n��h�ǭ܎��O�y�ς]rm�.=�4���%�ίރ<s��G������u��W���a��Ft 6L�x5#jE�w���Q�KN��n�r''�����ӓ���8��t���א���M/^�H�n0�$��ƤO������ rpBњO]�C\6DZ�B����ף��7��|�t��?��d���PZ��g$g�#a��O!5���Od��L�_�_����p�r�j&q�9�RC�*G/x�Ji O�"p<�o��C����.<Dԃ>e�4'ӟ��6�)���\���Q�M4�U'��b���?x���8m�j#S4�GQ�@<�����n��e>�Z�I�N�������v7��=#��-W�7��/����̋������{�)0i��	v���@���p7�32��ԓ ��N�yo�&�Ԅ�q�Yd"���`p
^�f:	%,PYd���c�F���셹�=a��ků�2�[�fx���_�x�$L���p,�@��r.���a;�f��߲��'���pm6����Q�;,��z�wD�'��Ð���0��!M�h"=[޽n9b��N��e�l�*|�5�+̸����L��B=�ms�ρɹ~$��������3�}�H��1䝃D������9�=�<2�,�r��w}<f+���#Eiå��²�>�|U�Kh�t'�T`'�m�����v(K=1@�S����
X��i�P6��*[ӕC鉠C*�`���L�S'��PNq���̓l2{�#�Ky�!lr��]����:�5z��������r��p�%ᔱ�o&��c�u�PaR��R�ڀ",�#=]����c}� Ґ�8��N3&�cm0i��i���Op�͟�������#x{cf�
�w�Q	wa�﫜�Ϊ��FeHB���b�.'����j�Q��Q�R�/����ṑi�P��E�Q����^^�fG,L~��}�l��,3!�G��R7�Z�&:��'8�� ݝ��䩾-��]�|�1�m
�-�dQf>�CI{���9���]^�V�������o:�^�V�I4#�Z�%�!"N-��Dm����Pb��|Z6Z���N�yl����>-U��)Т��B�A�)B�	�3�	�S�pI�hK�Cd9bu�;�&���2�U����F>��ҴY�\j�|,�=G��v��j��������-�	��H��O#�+(f�J��8n$�:y�E��h�����o��Ǹ�����*�WO7�D`�8Q���I��N,�F�~�����3w��_�x��x�����=�7�k|ܔ=i��h��U�o�I��G�A����"O�ȂKO]�I_��5w(G�{D��tp27�
�8#X���Ű��x9u��bm"o�hR�TP��c�m\[Zl���i�I�m����I���Z�G�(�3��4뙶��H��Жe�������RIn��<7�~%���/;���yT�U'N}����A��,XЁCT�;H����dG�����u�ޑ&b�N�3�/�]��Ώ��1�@))����u |Ή�Wx䵗�W?�	���_�Y�#N����į�pV����2aB��@2�bj�b�\n;�|�r�y��;oǏ�}�z�9<x�5������*���\k�Tg���]Ϯl2xꌥu��n�بÝ�܋S�F*$25�"wL�S2L��]lٲ����uN��\c�&1G	b��O����++�B�.Y�B$�ȴ�����E-��
Ӆ�yÁ��|Z���9^�e�0Ɣ���J�i���6F"2m�3� �&�	}���ٛ�P���Fh������Αn�����n��j�<w��"?K�P�.N��^�%���ZJ�\hM8����vS���Z;s��
�r���?%V؛�u����E�<�Pr>�7�b�M��{ygC�����X�J���F��v>�4�5�'�g�����ǥ�Cz*-�	J�&�	���G�=8O$�E�<�cf�Nk*��՛p1e(��WE���DZm�Z!c�s֨�U)T�tRc}c���uT�Ns����[o��_�n��J��мl��>��/a����k5�`�֒�4�\�Z|t��Ƙ�̮���.4�ʨ�;���ï�?{8��?~�4}1�`u�����7�N�.��#3�i�;U�^4�V�ĩL�rѼL�Q�]��V�`����{4�'���8J��Q���&&�Y�:�3��*����s�`�t��6���rн~�њ�l�����"%g�����/E4�C��I��r�\!�%���lP�
"2�?�JS@�)Y�%K^.�.�X��;�z� kV�c�6��sݰ`xߧ�(�����-<�����hHo�)��JPR}g�����:b�n���xC�ˑ8m�i0G��zq��(]�$Z�k�}Y��a����~����,��q�-��yUc��D�D�d6���㮪:�G9��+���ӱ�5��_=�S|�w�K.��p������G�hi����&���k(�~}��Gǘ���ӫ��?�x�~��{����|�~�<~�m�۔�c�j���L�ՊNH6��t�xmc���a�z���y�ďp8,<��5n�f�\%H�IÖ��^�R3<�1��!��4$ܡ ��sm?W�#ʢM�wq0�3�rf�&&�lI>I��9�c1�m[C胶�E�E����XK���.��B;�]W�'����"s�`NR&��Q���l�{�v�*n��v4�#u�V�)� ��B���6����t����2�?�$�Vm�
Y+XE` 6���$�Pd�`���7���7�'x{m��������� 1��ɓ�B�O"�f��>RF�("
�I�B*;¸�%:��̷�����};~�[q�����wz��~����a��h��h�\<��?������9pDO��p!����-uB��o:r�$<'E��<���Ck�7�쩣�7-L��O9�6	j!�
�&�� S�,܈j�.Z�,����,�[��?�����@h0�
�����mp���c�a�~�	LT4�k���6�|^VD�t�~G�݃�Lvt�n�>s�*Z���$@�,�D�VP��'GQˤ}"R��d�6�Go�F��Ʉ�ָ�I�~[���ާO�xMl�\���es���ʦ�RuUc�b�Q�F��Ͳ^�wCŗ�����0L-z�\f����Q>^�**9��hZ�+)�C�ul��R�u�p�׹뻼ќ��c��q_NK�T�f���M:�	b�,[F0R��t@��t�-Ox�+�cA��ːa�~�� �.Z63xZbozm�Kኊ��L�ْ���C���盰Y�kzf�3�w�ht������u�CL���	��q����p������Ǚ�v7�=�N{Gy��(hMv�B�h���	'����9�Uǵd���^���O���o����}��]�י�ڞ%G['ͧ��F>ʆYG��6��w>j�	wf'}!1��y|�&�i��(�z�wRER�~��՞#�aF��6��tM���墐6�%����OJ���n]
D%�ƍ-�h��US�X6� ��mA~����p�yp��n7�e�=�e@EA�Zu�����
�8{��^�Z���	'kD׵�*�k{��=y�zo�b��2` �Qy(�ܪ�3׾.0�����g��"��t!�E0D���GPl�JƷ�s�W�W���Z�t)�a+�?!�����wt��g�]���2C�{��r�����BG-��.,l�lY"�hۋ�Aa��F�F�{����ԫ���UhTE�Dr�>YM��1���<T��1㐝��������N9#lfT���6���u֤�'<3Q������^E����GQ�8��ןw�=����œ���o��!|���q������Tkk5򿭧�>��]�y=F=�Gn_ɆKV�������S��E��`l�Aв�e����֠���=��Qo��N�LV	/������2i��G����}#��:����t����'?�f�?o��7��[����b��ު�J�(;x�
>��B���u�����M�F��#�N¢��m��0��50vE��B�"P��*�VnAQ�I	ׅ"|�JM�wU�.+�5&0Pk�OV5�|��	]��������� _��:�8�aR3,��C��F^ȨF��"2RE&��^X�Iе��W�#�{�a�ּ��������y��p��w�<��8���l4k�.����d��xA�E�
w27BJ5�9#KF2�C5��u8MV�LhVܗ�Nqe�/�-�ǿK�,�ʦ�����]QX2�-X����=V���f��e��|�Q��0��>�+����9�����h�z`+7�\�0�h��5.-��r��7 �K�f'	#Kַzm�9�3E�F/#��I��֦�|�s�"9 r�iRd�"��@�?��X�X���}ʴPW��"�+]��L�=�⑅ԥߚD/��r�w[����3�;=g��E�����h�H7򗜧�Ч<�9�nl���l��c]K+��&�x�(��鯃6�>Ul&�����d[Qg�)����}�cP���|#_�f�r��B"x�E�w�;�*�K��Ɵ�|����H������6��~T�ow-ɨ�Q�][�mW\���r3��Z\r�iX�ArQ,����Iw���
��#�j|��(s�Qyçw������b_����.���O�O�	���5zδ�㚼�3��ϊ�32A��E���B�����:� +���m�l'�(�U�m�2��'�.Մ�iZ/B����y�ri�]��hǶ�J��ZH�K���/I��	�鴃'��L��$��T �d�?f"9O�#�v^�!��,��
��{J�t㉎
�Z��`�-��Ȗ&���̄.�VzW��[)��w��CϻУy#h?�'yc�B���.�w4��^����O�L=�	��]	̷QNY"H�6^c�f�(�MR�&�	�f�����pT$�@��D��O����8lQ(�;���q���L����K��2q��C:�
�_o���!�l�)���pS<����_���������5�3��*2�jw��e=�i����,�	���^�&~�=��Q�%�����<�q��O~�><����#O�'�^š�>��]�2rQ2F���nx��k-M;⽎#�>�L\/u@��8Wm,bj�=�[H�j���t��#��g=G�@ �9�SD��ɂ�sZh������U����^�@��|�<��6���C��R�.'E}pjȡ�*��;<GLF̄�G6��i4H�"{��E��a����}�q'{�Eג�egz�z��O�mq����UϚ�8��?�}r}���N�^�chl�.B���2Th��^"8�������9mzJ��W#L��ԇ�����?��=����q�g`�M]{#c5��!dF�$X�{�(�/��MK�_�<G�rd"QvQz� ���]��/���Gx������^�O^<���~�~2�Y[��z����'��~��L�1��I8=G-gr��U �6J�~��ܹ�D�ɛ�:<0	˩�����Z��䫜����1J���=���5y�1�-'����,;�VX���X���*
�u0�o&��b� �5��9�![l�h!�A�m�s�)�@�B[�M��>]��$h,1�#-��K6F����-�����ki���Q�.4�+F�yAˡJ�D����Z��Y�F�cE]�k����#ߑ!�4J��޾0��'"l��V�U�'K�1a�5z@ܘe�'��C��ƕNB��{�N�s�2؏��js���)5�MV>�D��'�y�I�x"���GQ5(��	�)T@mCd?�v�����G���E�?��/�˷ތ�N?��;Yw�CV�"\��k_F0h'���`��[���M��.��d���B�T�k+Q���Y��ve5��4D��x6���������19p �sU<�fbG�S󙞰^�*�ЇJ�C9=��*�l�z�2m��c�ډ�����0	�s�d��ܲ�J<�F��&�~��p�'���s�f��6A2]^!i�G���{\eJ�T�B����It:�;h��?z@I�³+�����w����	��u)P˅K缾S��R*�2y=Ч��M-��)5ը���Sx�	 ��(xB���ֿ?s`��Q�1�K$�T�/ƚ�������iz���@QY(�J/��J8|`qs��� ��/q9.��G���R���f谦E����ǈ��7�F��������ڿ���O�W��k��Y{���}�3��2g�s�,�`��7�����m"�r���aBD�����+�ݧ��O�M�����/���?�;�s�������;:U���~�T�0]7���;�S��I|��;JLgC+H?��,Ը��ȕ���.��;�7����0؃�0���@�S�5�7!!�Ց�����+�^P��ԡ{��ȠŃ�3��iy;��Rj��H��<uT���w+b6�����4�7-���~�s��eC���MND؉����P��:~� QtM�����Cm(:�Ԇ�r�h�\d�&����ڃ�6����k?}�s����o�������*FΞ�"_X
�?�+�W3H��t��&E7	�&���G�����>�x!c�yv��ݸ��+qߍW���?�3_Ə�z��0�����^ooZ����̓U/
L'M}��U����J�����a�6��<u�S%]���W�ՕE>A����~�!m�#��(��dDiy��&�H|���5-6�a[Av~\�knV���0O묘��塂5HF��@�	��O`Hd�ш�v����S���&%���8k,פ5
����S�v�&���6�ʣH������.$ҿ�aI���վ�g}���Ca��%/�����O�њbm��N²!���<����L1Gni�`��rSYș��)��|�<��ן��;nDf��Cѩ7"��SX�v�Ow�I����ݲ��btl��݋_��V��}����/���Uw�#̱I�29;����1<�c�ʑ�n���7k�����#�����Z�u�y�ߪ������ݳ��F��FV�7rר�+.����s4��@t>�N��1`�EO�����a)?|]nzמS٨��r�x%�8!��1(s����Y�|R�V9�񖜨��$l?�p�r3zjm�"-�2ii�
��z��QLҕ���?���2���L�\��+�L/v�H���һL�\��0�j��5U�>�>��(Rƒb�YT9�̣�,��L/�Z@��s�E@���g�5t��T�<�0Yu i�^��*lg�Y#ϭ� ���l�Kkma}��$����]�e�L�=�9��I��#E������F�Xod�ck�����W�[�?��u~�kq��c�Zi�9�b9�N�T���]ԋ�$3��_�EmB(y6�ճ!�re���ʳNÕ眎߸����[x��A|������k*5:Ѹ�0��ht�u|�A3Z�'C���ɺ��V��
��"q�G�H(Učh!]͂d��<=�(<�MO]���+�zꧽ��d���-0q�M�Pb�e���Wn&M�)W�#�[H'rh�b�N�fü�-Ϣx��/b�S}ҕ�'��N$�DKf�<i��|v>��͵�����hb��Pq���(1˔����H�K��,��.x_��X�3Ιd�m��x<jn�bcu�N�����������^�/]w�r����s�Ҥ��Ǧ���XGt� ᄮ�𡂉`�����N�y^�h5�N����օ'�8ϩ8��[p�7�h������{�q|������	>>���Y���бa�{f��ǚ	:���z��)E�a�D}u�ǝ�Cϓ��>���/�Ømً;���=�Ah7gZqꏬeąJ�3�QnN�>�@uóa��R{�2�v���Zv�b��
˖h���3]�Č�Y��h����rNAs�Ɣ�޿R�L�2�WMϔ�����a9�c�YBVMl�0���	�ת��7�XC�i	�v����>�;���;�3n�XO������W��Hɢ���T~7�!�g�V�~��d���o��P��ܙ��$��J^��`٤�!��v�H�M��(jE
�뢤��w�ځ3���a&��Q��_z)~����ś��瞅�>�pS�d����N�n�S��B�)/��b_be���x����G�0�Fۑw��zY1�	xr
q�m4�\�06.,��tr��#ۄ�;���H'���?��;�q�}�#!ʗ�8�3��I���4�ى��<i��]�%�����g�P���9`���cO��b:��/<B�/k�ǲ��Q��Ͷ������9�����lZ_a�W�� �V��z�l13��u�4V�WҦ�PN �҇����|����ާ�tA�*r�zؗa���m���P�h�5��|<�I� ON"�j�tO*�K\�%���fK|�`<$
���rwʶ��fE���8�9�l���mSxXZ�E�M��=N��Je.ɤY��i�>��`�x�4F�7r�s��X>�V�����p��G������}7^�3�8�߀dՑ�[B}�.�����q�E��d�#H����r�������ᣯ�kS�+�9��>�z�8���^���8<p�78}��Q|l��n�%�"޳X��cI��.)R���A�&Re-��M4P):%����b������=���v|���|-���0U��m9"`~g�\"���9K��d����u/B��(ƌ�)�W�](�}��J��}ei���l�{fR�,�~TVPҏh'O�e�ρ�v���!���cm�@����qz1b�����Lp�}O'�wQ�#�d�<��
�a��$X���.����Ƙ�Tx
|��7����/~����|����UW��s���q#m4�(�B����	��y�&'�N�=QM�ۗ���m���%n�Y�*\|�)������ﾋ�^y�?o��\Pm4�MC}�ⵈ�Gפ���f�I<�����A.��to�Pa9�&���b&��OƑ�.;��1���26*��d�(M;�fG�V�X�����ZH8�)y-rj(�y~Bq�y���7C�(���8 �R8�H�u��XX6��	Z���e`�
t�)�-�b��a2���8B���u`���DZ�Ʋ������+�쬆�VHG��FI�B�0�q�0�١�u�W���s�t���-]�W�-���iJ�t�d�H�E�!=��[	}xn����U7���&�K��Y�/�E�#ɳT6�3���a%�T^ԑ�L�lq-;�&\��`l@�P�Oz�dF�[��`������Mt��:0����2Y%3�b��84����m,{:�G# M���st笮��.�}7݀�n�W]x��������x��_�_}��u9t�Aķ!8a��WE�¤+K<T&��
uB��\$����!�{�-|��Q|��kq�ڸI7	W��umb�������#���v��W5�3jU�c2�c(i�p�Yd���*�XV7t�GcB=����;�f�I��m���Z�J')��'��y�~�)3t͗6Px�}�\��
�m,?>�ZR�j�\V§�@G�Y:$�ڱ"�$���#��8�G�lf�J2x�/�8m7rmrہ"��T^���oE�X�xP�K��7Sj�6�E袡�p���Nip�|�&~���%=�����²��e�ED���uN����0��o��#V��/���R����Rw$�I5x�۸y�"M������$���ɼiu�.V׷�.��Y�ya&E�=���(&�G�Aa��SB77S�0�Hw:��(�pq��ǎm�\0�>��v�Q7�^ߨ��^��?�
������+/�}�\���_�N;��U�Z-o
r�N��l����c����IN�Q.���^��Z���F��ܳq��g�w�Oy�zO����~���&��x<~'_��i�����H���\��iy����E�I2�|�um�:��!�$�e�Mb�)y�t����@���Mc&9H�>#��^Q�k�~��m�Z�XD�̺/9�q��4��ܘ-�����S��h�@����v[4\�+�k[m��3f��u�~=�Qހ�tm�dhFs:p�b>m0h���x�nitCKI�Ǜ��*��L�K��K�r��$��tJ2r�o���(��������nF��� lh:�7�� �F�'Gq��K�Ƴ���]�q���}T��/<�}���#_T���V��7
�[j3c>�퉩�l�q�	�kM�k�<W�}~����'bm}��T�CU!yr���AR񮨉3ĺ��#���C�hP�o6Y��^�&��v�a�\����D<]�%�)O�d��-=��1�U g�>�/���˹��<Fu,ùk`i~���$X���q�0���h����rĥk��PXi��"h��BV*���6��7�Ŕ�vw�u�'<v+26�ozҫ��]I��`Q������G�
��ݨO��~��|]����a-�p��� t-�C��?������y���|��PYh����=ΕXۛ�8/�S���Χ���&Y��Ѹ�`�����j#W4Τ�i0����)6��(��I�I�~��?��瞅���q��w������E�p��u਻��
:�Ch���mЭB��:ݗN�D��Q��ޟc�VM��#�x���I��s��_~�!�?}ϼ��:��?��?�Y�����l��&���7iԜ�o�Q�������0>[�|mCv�{jei}��'���;,O���V�q�#�H'�(��o6s#a�p�hƾ�/�|Bc�}	zL߆β!4��㶐��C�1;�$/S�6,�~B6�����M��!�!��v��w�l0�)3�����:��)o-0,g�mZpཥ�,�Yq�B�.�.��
�������j�4/U؅�6�>}0��z�d��nâ�'!�Mk1|�H�Q*uk�T�J%�U�d�*lR:"m���HZ�m�j'�|�ϴ���V����Ji�n<Γf�����1F�4��,��ǆd²�G��l�l*9g��]ލ�>�r����obt�w���w�~��}���G���Sq���񏮿מ�;�,������O�a�Y&�f$c��v���1AEו�9�ʜ���.�Uc|���p�%���oÇ��3�#͝������X]ɮ(w��k�wz���U��(�@��*�&y��Tj&�+���e=�]�nJ�7�\`q�$1H'2?�,(}$���6��EB��aw��*�}0ݶy39�P�HĮ�6J"\	w�D�gs�[��e����a;"tH\�~����2>�x��98N
]�_;�ļ�$ )h�0�m.�a��
�lJ�[��q�!���p�I#�W��Z�dx���\��4r��Eh��IC=WF.`����p���K��^�9+>w�%��;n�Wo�眺��4�h�_�X ٓ�D���.�@F[�أP���NTO�bF8}u/Vv;b[�;�	Ye��u�o4���ij��0�'G���JW��8�>$Cl�n!�N
���@Y6Qk�@_�l�?�%�F�Ir-
�:�g�H���Y����?�1�~Q�����ᅝP��dܖ��p�½�lO'���霚/��.����[�B�F��=�LY����{X�5*7��(^�(1.��j�C񿬬)��C��'Ӭ^DQ�C��e�����ί��2K\Y�~�+������, ��=0�x&'�CZG���p2(�� d�f�SO��|�p:�ү:��,��7丞D�!���ĉ?IV���`d׏amcW�v&������-7��.����ȟ���iw�,����(F�a$���S)Ɉb��նvF��>��x��8x�~v� ���<v�-���1|4cz�y���X�6P�OEe�*�b9s������މ�N�)8���^�Oc�52銝 �$��X���o��r]�Pҩ3!pr�%�� O(�Jj�P�yįw�z��*N��Ϗ?��%�:XV��ݒ3O�N��,�����:x�紤�H�t�ܲBڮ�y�Q|��m��)c��Gd��t��ӭ�S�<�_���Km�Eb�6�ߴ�4���U:�i*ڵ<y�����߉
tM�7A;J8h�p�R�e�Ş��sn(m΋z?�e E?�T�&.�Wˌ�}��@��>���b�q5)b���:Z�mT΂���e�8��5\+(�㳅E�IK�od����a���E~f�xj���\��x�TS�rz��*����<����=��N݋�_�����q���={`7�~jCd@
f.'ڃ�Zҟl0�P����a�G��_��J�Q7�C��c��S�2^�tڴ�ѫBt�u�VQ�smܰ#���M%���^�=�PE�k	{./�V��NQ�%vi"�qR��Q�VD�g�����K?s&s��L��~Z�1�l:jF�����@1/mX�y���]�9�D���;���Dba����D�<�+`�۽��y#E1B�WpVi����r�8v�����q��:��2��
w3� ��͹�M �`:�u�2)�b�����A0L&�p�Y��>�<>3��V������p�]YAu�
�� ���[�������ᛸ� ~��q�u���}�0�L}��'i��k�|f����R�1q�"/��vP�,�����p�Z:�I<�Xl�C|�'S�:�p�[�}�(@�{���p,D��G��u"RhK��^���!f�Q+J��C�6�e�`�i
[���WmDaR**��˲�@K/Esm��m��獾U�7��r'������9���Y�,��f�|#���u	�7q�[����C}����K����!+�%�j�����)H��M��m;9� ��-~�6�xU�0R�i�jԧ殒��g@q�����7�\Āa�`{����Yւ�
�)��K���R�[V�H��oH�]ǡ��"��EÙIˡx�h!(�5%zmS=9�7Hщe.��5)�|��A<�己����IS�t���Q�t���O�_��6\|�x��3펆��.s����$3�pI����7�!��WU2��9����[(��`�(^x�e<�����g������V����Z�)���sᇝ���"X�}�!�w�x!��]�b�	����:��&f!�w���"z9�\zV��lϛr���6k[�����CFV|7�o��P�Q���*�~1���dK��3�%2<�q]�^�l���M�B�Yf�9A���+lh�^�X���g��`�sY�)����"���Y뮥$d�'�w�t0�/�e�;����]y��Y���lWsJ�͌ϒ^���<�,d¢�ͼ��ڷ(	�v�.z��M���>9�u�-���$*�A���[|L�N��(�|`Yz�G�-�'RW�;��R��,9���<.�G��dT�����!jU�h?T�Q�yj�W$O{0��֯�K��@<��4��U\�E��gN�X[Vv���g�|	���ؿ{_�n?�ꢣ_��V�`c���:�}&���6���:C�<�!�{E{0���ْ���W:�o����i�
f#R?M��A�MzU�ޑ�x�iK����r8�x[H�-߃k�}h.��s��i�L�+V�Q��'{qkm�%Zߥ�J��ְ>��Uv�n�����LV���1>�@��S��5�K���ۮj�<��L���CU��8Uk4���x��1�4kˌ~ӥ/0vt�}��Tə�,�6M$<��g}���҉�R��4�ڊ��2�ʣ%A46�y�z�7
�	g4tDn�b��Ok|� ��������7]�/�t=.?�\���#w
n�tR�TQ��d��x�V�Ĭkƍ�~� l3a�r�0�8êCޕj��dTM6|c��"G� �� 3R���ɿ�q�L�)��?�Is*'�
J?fZ�1�b��@}�:����E�-���3�a����,o��]&h��\��P�#p�����r�"���|�Oo!D[Nɐ�>'����r�B�	I�1���y�K�K�?����q�wa+��,�S�r�e�︺���R�p`kTiRR)��yހ���8�z�Q����<SYnv�+��Ef��p%M,�˽&����TuV�KG�xuqW�ң#�<�˴������:��ˈ-]]
]���j=@_�.�>�Gn�k���6pi��,h��*�4��ec�1����g��'\���y.)]Ĺ$�Uh�.]m'�9�������xU�����qg���b��)'c��.�JI�`VN*^(0R_��Tp���i���Q�>�`���������8}�.��G�VR2<:�"V�`/��F]'�.�%�'������w��7Z�+X���6�>!���:���S�����S���_4����
�}@<�g�C���xl�u�+�U�ޣ�Q� ��(�t�Q�D�X��*�1�����x�WY�H)N��c��g��'yWҊ�cڛ��blT�&�,�Y{���p�2<:�z?l��f���jZq��VҨ�`��8^a���m-x΋&і��ߝ�B4U6w��׶�>d�~k)��؄<h�o�E��͔u�P'zAol���VYL�HtY�W�"�#���5��<���%E�'�t���P�Ol"�<����n�5YREl�B>�m<�,�b�D�y���t�zV�E��7��ws���$�������'S/}.�#���M�vt!-G%�Ϛ�@i߃oX�i����ظ�H3�R�4��	ya}�q�3I	4�6��^K<��]�S%��xu������Y=2U�>`����8����1���O����Ư�z=��j\x�8�Z�rA=�N�{0Jp'�:��,?���n��d��6���Ц�jٜ7?Ȍ�W�`e#\95AG31�(�&�[�>C�pV��A&��!YҮ�������c��������Ms��.ـIFLc��R�,����{�@��f.�A��+�Ơ� ���春?z�N���w�r�<�d�a�;pXk��ڡ�ێ��[��!�7Ӊ�)���'t�	6ˀ���)@DF%4�9�fIK���TM{sͲ����Ǳ B�WArG�t�+�1	��P�0X1ߊ�0��S��+T�m�=��1<����q�r�E���]���x�;u/��*�I��N|y٠E�ط�ugㆁe���9�ľ��T�4W ODY��������N9W�r�|�M�bTcݮcm<���܍tu#T8�W_���V�/�Ě����yðzs����1Hg��w��c�eh��䱤�]yJv�-cRX��c�d�c|j!�aaU[.�����YPRj���E�=�{D�H0��e���3�~����L6��&�Gy��ِ��l�!a�|��Is�£�g���ѐ�|䱳���Md�l�i�2}��a0y��O{Zz-&<ۛ��'M��e�����bs�
��]��K]�/�����a�yi��6b��̹$:��F�@�������K��J�Ƴ�L��1�w����tz�Cv��6<u�G�T�x�!|J��y&/����M���\eI(�ʰz�<�y~�Aל��5�>3��к�O�Ώ�5�Uf9@�U��� �AF��U�g��FNU_��<&,&�I�u��#�����������0M�cM�q��ar�
��F�d(��xp#vD9�����Ȏ�.፳��(P�>\ǡw��ϼ�<�"�x���(6�u��v7YFXu�=ƐʾUt~7!*��;��>\��;���Z�>� w���8+�$��w$�2
#�0�u~f�^C�	���C�S8��M��Ҡ==��k�]���8�WY����q�%�3��O��i�i�yPW�y��5{�R�G��B���N9��@��0#І�TS �ˬ�Jvl%`j+��qH��5�mD�͂m��@w�Ĵ�~fr��b�$�q�Q~��ln/ǿ�2��ZBgYV���OS�l���?=!�������(�9�G-��|I��u�{}�s�ۥ�h�Z���|�NA�m�U�����؞w�#�~ך��p��)�ؾ��i���B�)������UN�C姑_�dj�ߐ4��A�3^��Rԉ��O��w[���X-����:'c�Fa�cylG_:K�uFy]s��aE8f�Ā�Q�g���P�X�9�;��{+��v�Cz��q�y��M$G�½�Ft&�Q���p���
\d�����.��Z�}e�h��o��|��wq��?�{/���y#��r�:Zi�~�y�[TtJҹ����&T/ީ�6^Q	:�XǷ��u��8�޵�W�s..��G}���fݬc�9�78m������ږ��AH�g\P̙�n����`D�8�R�R>&����r�h�g���c���n���w�}�)�^�e��ZA��2�wu�[۲��-����,���擏�Oc�m��'���=�_hL^�E��'�k�k#���בfPd�9�_��R#ϱ<��F0�����ꎓ�S�����t�/�����%�Jk_5t��բ�:F�&���>m��ڹ�ƈ,)���9�X1yu�#c������EgL�-t�����?~��x�o��Ʒq�E��7>w#�f?�;��	2��0�*S�x�ß3�4���4�Z!9������E"�.����k����O~�7pՃ���O=��~l4�l�.��\زiI\a�&��Q����8�6S�ʎ�޶�ÊG�1ٖ<�Y�W��A�J��R[�U²(����I�ui(���ݥ���-�5O�eB��3�(F&�W/Y�9:,�q3��K�[L� �D0�S&$��}I��y��J�	iO�0�����p���j��-��m4�F��1Q5�(�sA��h�ʮ�W�-ú%��PBB�۔W(I���)/@�+���O�O�,^N�����ʟ����m\`�7K��){	5Sx���zF��ꮵ]J3$ߐ��*��������B&�S�{�<,�g:�?	u��nv9."��[.A�\5�<� b�P4�͞��#,{���e� BrW0:�e2mt��G�ǿ�+������t�i1l����2B�)�:���g\�N��h\�Ty��Fc/k�8�Co���^>�o��	<t�^[?��++��q�s�1�F��*�]5�����PW6�l,�i퍱u����/�r~��p�?���8tj;ʟ>(��Im8s�Ԉi��<{��<�d/��L�d��-;�C�oA��.QE�l޾e�'[EW4��e��ڶ�`ļ
�c�w��i�ѿJٟ��Ƙ�ˡeS���hy��}���m"1�ƅ�g���$D���$�TN�oYg��_���{Y��L�r���MX6.&���xk�+�$e&;"�?�#��J��n�tޠ�ZWџ#Sx�˝UN�y��=����2�G�o��':��2¥�ݷI���6S���:2񀎑�5dϿ��ڼq^����Z�dP����]�6�����C��b$G��^\�߲<�}��	�F>�	%�5`3Y�m{j�*�\�S�_�����Aё_������(��^BЌ*�/�_���:�d\�ul�<��|g�W������v#n��b��{w���)>�����s��Y��Eoq���θ۱��e��58��o7>�~�^��=�>�<^��c��k�V*�Dy����sZt>BX�U�$�p�
�bΖ��@�K�,�
Fsm�_&���D3�׺�P���'�gJb�;��#<8Z�֕��~Xı{�t�N���%�=�{`hs��d:~E�p��v�s���/:]B���\W���O,v�pk�d��z��B2T�J��K��z&�Ӓ��=���ќRx� ��4����Q���rF�Y/�����<�8���F���xu���k��������]�/���\��.� g��/8}��K<ö���=�Y,�}R�� y�&c�����bE=���1���|\q�9�������_�cϽ�_<��|����p7ι����"b8#����}�]P����L��KNjڷl}�tSc�*�O�0&[ZK����k�i���7�a�L4Zl~���s'A�%/b&z�/]�f+����'��J'���@��͔�2����|-*�"m1��>�=�M���%�Ӳj���:�4l��#�-DR#�{�1�7$-sۨT�6���R�%n_��)�K�op��ڌ9ߝhP2��2P�DH�2�ߧ�CǘY�6��!�O�.��ڶ)/7�!�����L�a<5yȻ��Ѿ�Fv�Ee������O����{#ׯO�G����rFҚ�Vש�SA�NY!�	��[���N���W�g�ŷ{�}�)�0k+���(먪I�KU^��F�nr��)HS��T��U9��ʙR���!O��r�S*����Z�"%u"I3Y��ϩ��/m'��"(q��,A�{[�6���r�z�[�["�֦���;�O]�&�5�$��"hN��~�B�A�W��Rܤ��p��ɝ%y��o���)�6�D	�X3*.D�+�ބw6��p�#��w�[�%P��PT�8ۨq�J]���UKQ��/$�KQpVA�.��v��ZR25�M��t��gP�Z�X�٩�l!��vu�l������n���p^��^^؁�X��):l�8L:`kzZ�'O���ōr�;��s)�ɇJ�W�E)9�$(N�*�K>�rqI�� �(�Z��e��>�h���t�f��C����c�Ԝ*�Jx���w5i�Sw��ԫ7zǦx����O���]|�j?��J\{�98e��C��$��v���X19G��t�������������vׄ������­�]�Co��G�~?�<>�s�����]�;#��������ǧ�m5��G�YH6�:ᦧc��h�zԡ�n$���w�ʺF���������c�;�i}���f2�i�&D7!�66C�t���b�xÂsҁcXfɭ�H���&.3�X:g�"\���!��2��� �gR$���@��RJ�5���1�f�������Nu�t��"��g�F���q~��v��Q���o�?=���Gp��g��k���^��/���ۋ_l�\
d��&��ⅻ��f�R�UQ�J�6u'�l2�e�6�\�o���v��mx룏�����Q99tG>����6�k��p�NW#'���a�O��DO�� �$��'�C(LK�'�-��A%0w�<��k��RH��FJ��eB��r�t��vm�q���0)��/ �ˣr��4������f霹H�S�J��IWȷ�w���:���
,@n�DfB��'����H��)<#_��=-'=�5����G���W@K�+V�i�\��Y|Ӥ�S9*Qp��GL,-V{�:՜W�+�)u�Pno�<�&=LWS�/�=�x[�(��*H��,��� ̯Z"(9��¯˰�G�f�!*�t���%(����ϗ�c�k�ݔ���,���=��֠�|ON!-J�)j�|���%5�MO������K3�qf]�O~�7q��Z��'pW9f�� �5�M\���C:UƝ<Rc'���
�j���dO�t������>��M������nh��^7r�0F�T.L��mq:��f�5>Ȇw������S��$�.'��O���S�7����H&*�����̓s)q\��K�S��I�F �i�u���k���E�R�PԚ�N�C�e��&I���$�a0��t�Т���睡��-'Wr�bC�7��o%z\��I_dI#m��<�)�ڸ�L��6&h��lJ�2 ړ���i��#��Yl�d;$��U��,���ɩO��-��%A%�7-����Q��t^��V��A�P���ZS}�=Ի~��yRi��U��0X��+`"5$�ư�
x|F��J�y��2à�i�қH��� 3�w$�Of��C��S�p1{[�z/�?�v�R���Lo�x�՟%Z�E�»"��{2���&pG6¢��,.Gms4�{~��EA�y}�@�Uu؛q�Ê�h1�l2��K��̓�q�w��.��\��_r!���"�[u��4#���k�������|w�H��<12cwP��L�Q���:��F��ۼ���3q��t߽x�����ǟ���}O��6�=���j�2�+��$!$�����OV��Ðㅑ�Xt��k4�ӶE]B6�6Q�.0k��HE�H�В��T���%�5��R\�}�����A�O���Z��3��V��!#4�*�um�������?:AG���$�{G�*���F��	����A ��f"@��(�k�2_ �.�N}��)$k�`��QK����'g���:�ʘ5���;}C���tt_��88�bd�p��5��άb��zd�CC�0]��6^�F���&Ϗ?x?��O�������ï�v�z���F�p�5bx0Ϫ1��@���B�����0�m�Hݔ�ʐi���g�G���Eq��n��w�����x�����S/��7>� ����Z��v���X�7���kH�"c�Щ��ؐ`ǝ<���̓ٽ[|�T�/M=S�����k��W,�is��Qڌ>�R�>o��ݎ�?>V��r;�CR�L�L�H��}Ȋ����V�_׀>ֆ�yL�Y�7���uv�`^����+�=�}��6IJ������̜��gu	�ͬȈ���ή����X�mQ�J�Fn����H�������eDt5�+7獳d/ʯ��2�g�ܢܡ+["tͺ�����|Z,�t,��C�Q��ҍE����m����ݬ��F��7z�>�M�h6�Q���İ-PrVX����}�F�)�i���*sޱ�y��)9�hT'^sA��y��cR��\�/1���U%�W]㓏?�W��	��?�G�d��2�Q���w��[8D��d��hh��W���{�9�Ǉ��Co���G->vz�h�qu�K��t��̘4x�+SFQq����A����~؟�s�El4ζ{�&:8$���D������RϢ����9w�}r9К�iN)���f�[���V�/y�~i�C��(m�w:�Ƈ���t,�9܉��|�g�LS�"[��[3_?9C���s��DK�ψ��.��7�&_�6��,�I������dSH�Z��(��ݺN �Q-�B_(?m� ��bM���K����bhkI���x[w�C��5�A.Z��\����涄��x#5"�e:����4e="��eH�Le��=�n
�8�BZۑ��/�,ծ¶ J:�=�ꝞN��1���[���|{X&�6�q<ߏ�����3��E��f����t����9�Y��}c�u@�}�yQ��<s���1{O��! ��O��z���$�T�����u��.��,z��j�B�L�/YV����6򸠫�"��e����`�`�w�ϪK���f�W�4������/���1n8���]7��k�ƅg��]~ǵ�{0���Ǐ�`�ȲG�<]E�QvF�z����`j0ݘ��KN?��W��?����[o�;O<��>�^x��q:׾�C�B�ز��]��+�&+d٢br�71�%����給����=w|��Uv���Lx1���?�3U|��jI�k�/"`�E=龎|v}~n����r�D[}j+� IO]�Rs��l6�Ҿ]�I������.����V�� ���?γ�Z{�.S���T�3E%A�Qzߵ)��Vx�-Լ��WR�3��a��Բ�pT֦�Dc��W��x]SB��p�
]-�[Y��rl�B���|�<��1<�����>�n<�|������pə��=�x�l���%E���B0��w�;AgF'K��l��4?����d�S��u�D����3O�%�܁ߺ�V��ƛx��C����������M���17u�8f��:PYㅬ�;vH�?q�7�3�~�?�8ٔ�O�d5��:m{f��>��,�%���Xݦa��K����vC��}k�6�Z�6�tU9h���\녫��0A�)[qlL����1�
�P��?����-�t��ՑH��,>Yd��A��읬�<�u�|�Id�L���D��<;{��'�ur$b'�ͯ?����,�MIF˖��VYzs:��{�����3_�E�C��+]��q�J�-�\�"�=��p�i�3)n�7^N�V��(�w��2�umz���AG�X�3�"������-�(������.(�YV�7�!l����1~)�(%|��fpӎ��ϒ�Pe:Q�#:%*Y�e�8���ߧ`�Y�+5 �ꀅ�m�:��ŮF�@#�'�d��h=A�G�[¶�䀃s`?v���������'>��������k�j�a��FQ�CNGv*�{2�rCv�>8�2ø	\-�8���y}��)F����2�C�04��dY|�h���D���g��<��ȇaX��5b�*�Z���uym����<�������`s4��?�n������-��aƼj�Ra�fXI�휳����87l��Q�Cm�M����M��U��tJɲ�T��D`麠@�ҙ���X9܄E�&E��;�E�H!g#��b��%B�'}Yq4��-���R:���ᱍ��w��+���V��G`�t�����[R訬��%Aae�*5���f!y-λI���h5��0�&���lHbA
HR�x�W"ڏ�!��������0T*o�%f˼��>���.��~�P���:���tO�efTf�"Kw�
C�g5��p�W��,ZG��o��Y�)D�2��%{�E�g�� ^?�.~�o��=උ/�����_s%�߻{�����dg_7â#�dw��x��́(�Wt��N�U�m�VI��]��S�n��<\w������W^?y� ����x�w����_#i��������^?�RF֝B��o�h�k=�L@�ӏ�0�XN�c�x�:"���a���o�A���N}��É$�n�$�~\:3�fd�s(��1b|��8�����W��
�t�!�+.�e�O�v�;?��y8��Y}V��m޶nqsa�~�:[P� �aRb�N3��e�@,���K�CtYD[�1���$?��~���ۼ -cDY��4ʚ�_aI��l|�N���d�z�&�*��)���&~x�U�������3����=���%g��=��|ԌE+*�1
��R��+�Q�F$�H�����*0����5�	pj��SοW^x1~�λp��#�ޣO�O?��N��ru�F\x_���!�I6(J�:�
�26�9�K3�S�d�y´��7�/23Aa��tР.�쾍��-*b�2�6˸��*�������'X:��B&���[���d�2�wJ�7�==�kTK�w#�t�i�n!"r��7�N��>J�C�붅P�?�+O��4�Tr�d�GC9�c���%�����4�n�T�f��œ��sk�@�@P���'"_��ܙ� mhr�}�٩�_�!�K��KI�$���A�[�H�e1�5����;[�S(�t��>���~%V�ct�s�E�Z�Sb:%���ս�Y���\��,U�X�*=�2p�a��)}�l�G!��z0�ys��͸@L�O�O�r�h����\�����+/������|�#����6���]>��qt��N�	�\���3?���p�nPkj���tv��Au虤�1�����b��NQQ!&�#�5�?�ѕ��)���*f��=���L��k�-�/J�
���8���j'��h���g���r�����6t[M��;(��Yu��Y'?&����E|[iC94�ӆB\_%���Wl��s�.���s�� �0r=�f��״�=�	���4�/"�I�l�VwzlD:crz�Q�i�b��اhJ��9�47SU�'��N�3��_J=��M��N�)���;��[���X|���n�߅�y��mj��i�^q$���͖ۚQ>�J�\�J�� C��dV�E��t��M��Cѱ�ރ�7#_.���^���L�[�PA�1y[=�y��Ȏw6]!H匘����!W���D��1r��S��c�^��q��w�o���/� _���y�e8k�>����Qz�
��2��e�N��V�/�bF�YŶ�^��h���	p֮}8��q�W��w�<�2�������Z�g}2ize��I��L�P�+�2y첎��=���Kk�����M�F�X�	'�ᇁ�>R��5k -)�ǎ��%�pp�L��/KA.(��%Tl7��P�:�.K;v�j���ɢ��N�Y����J�+�l�Z�A����+�h&$�Nq&!�k1f�+���t׌6q5������, `��qPJFϓ�C�*Oz�W#���Cv����C��uN��J������z�U����W��7_~ �|�'�B#H���n��������iA=��׹�N���dZ8��Ϳpp���kW�e8�O��еC!"��r����ԕ
�^~1n��
��O���^:��͟��_�ǣ6&>T�"F�/|�3���5���'|��U��zn�d�yP�0�~��;�im�g���6ҨS(�� E��K�}F7���o�^�:���$K;�M�esHn�0�穯�u�e��������8��B���DrL�̛Q/l\H����z�a�##9]ވȆ�BRY񺥮��(����i��+׹Pf}3�aI�ȿS��q�gMdt��S�ز4Q�������z�t�S��R�����l����Q��w��]mK}��L/����:�f9���DS����G-b$+㒿��Ж�������-�6�o'�t��9���fp����U� �/���'���\C��VR,�9��V��Mq�n��n"�'~��y�)�F7��ao/y��xæ�2�%V�i8}d��s��l�Ò����_�x�=��w��noޯ��c�p���O?����2~v�e�;Zñ�
���fҔ=	!~�f���a��1d�y�Ӻ�)��΁ݵ$:��x��?2�$�Ǿ�Q;�n��M�£���<�ou�h+�*fg��瓖¸��+k&���&�L��-�	�I�2�\�Uհ4�cy�O'�����c�%-r�p�F;�.�q�����ID�#���x��D�Ch
3s��D3�fI"?t]�\�5���R�׺����d�o�і�t"��	�tɊ-�T|^8�Vq���P`�NI�d{�^d���t���q^�����։89����HLg�o��/��O�)�)�7�n���t*��L�^dy�n}�9����!��<-.�g��r�,o��w��C���%����t����huC����龶s���Z�� �Uv� 9̤��g�� 9��6ȴ�D����y��B��U��mt�C��y��ɗq٩k��5��k�݈/�����ҭuW�o�2���9�p���[|=6D(G�׷���)��{W�����IĥkpΞ5|���;n�����ȓ�w?z��&�i���S�$�x=��=�Թ|hY��Q0Y�Y#֝�m�U��6�#iz������hu�h��ѵ��a���́1��������Ƶ�~��S��gg�t�d�����`�+T�t��M�!������x3*�z��א�1�}`��|2l�,�b�����fO�V���t|/��4j��6p�΋��m**UIE�L�BR6~y���YhA7�V��a������\y#�c�+��ꈊ���]��0㷚�_{� �q�0.?}n��b|�����F����3Qձ5�P����yc��H����F��>w�����s�/�|ݖ�ub��k���+��M���_|�G����^[��]�2�!�a҉�\� �����E�@?�fa��V�s�P��ٓפ�R6p��Bh���>�6:��f'��F�*;���UE���R�H,��
EEc�W0�h�s�R��	e��/��K�}�G���u�CF�N-���%2�
�S��y1)G��k���SR������OV&[޴���ʐщ�K�f*��U�t}���n����+`UV��uAdG[_�2
�^|��YIC}/&�Wn��i49�X�����V�����W�U�9Z�+D.[�l�����BG���@��c�R�#��з	Q2juѣE��0Juu�S��u���M ��dĘ79ݦϮz

��)<�($F.34V���v����|�x�Ng����D�:u�c*kV�֏!E��|e�f�j'/������-���D[b�������o.��u�=���:�b����cy�<����6�f)����W�kww�J���Lqƞ\��\|���������ï�o~?:�sx�c�>���ȃA�p�4�F����������gЕ���:lV�uI�2ʜ�U�$:����CsddEp�J1B��6�L�	�E}|���䋢E���R~ t�<(1h�҅
�>D�����e�r?���B��Ά�-j��,�~��^Z�v3Tڟ9uSƚ43U�q���V��<|[o��2�N�o����r>��Ah�^�����%��&Q^��f
�m�72�e�h ���a��3���K�79�+m���5iҍ2���@��6J���vY��Q.Y���
o�v�hSqz��|pj�q��kzW���G��w�P�-�.�x�ڐa��"�{� ��>.��g�1/:�Wv�����Y�=tiN[�їW��W�Mڙ���Jħ?s�wV.�lӗF��,��C�i�Zd�����]����Spۿ��J��B�֞�7&dY�_7�W����vb;��?��x�\{�~��/�mW_�3N��('�d�o��G�"R��j��!Y�#� �ɼ)|ڃi��u��#�����/����_�:���S�d��O^ǃh�_�P.]���ԧ$�0�ߵ2��[�r��dorE`�0Dr�Ĕ$�v��+J�%8�i�?�u��w�\bzF^G]BBN��L�f�F&��/���W�0����A=���{�o���N�W��7  g�$@� 'p4II�,Q����m��L�W�YV��������CguV'���d��n�nɶ,QI��8 A�8�$8���޽�rj�U��T�� �"���԰k���w�*[K���!�9zK�s��,Q`�s�}�!�;'���$i�$t)&9FR�A3�?pШ`�4�NAd��J��Zh4�Iݹ��ڍ�$�~�cf4k�d!�<�t���W�tJ��Ԗ�R�Cu*��pW����z� �쩃���'pK"��w���R|a�V,i��:lX�,�R�Z8�]uh3{)��8�fE�@¼c�s�����q7��e��?��,�AL��G͝o�ͽ�J�BԆ����!��P4�u��� bπ���w.E p��.��)Ŧ�"����b2K�����0#F���1W�>�8~���d���x�ox_P������Z8����g�<���;���h���0�@��~|P��)c�C'dΜD������S����l0�~��cm�}�9ΰ�����!�7���p<����<��/��D��ocY�f���8��XS�C��#j�����f�Y��g���<]����ڗO�S�d�g�<��/�O-��6�A���$��)�\&�s�dt1�b���$�C� 'D��#�/��</�fF�F��Y:�w�3�?���I�V�1��3u��D�I��o�xO�e=nB&r�*�:'����|���|+<?^�ۣ1��w�bi��|֪x�*�"�;Й���;�fs.�����ҶĂ����B�
8�����ō����p��჏N�gO>�?��x��w�~��6�@,.WZs�O���0V'ٺ��i��x��S��G�@�ز4�����3���Bh#l�2U0��<��Ǳ�Q���m�î��7�'��|"0|Ų0|��w�;�G�H2�:\Q�
�9:�6�<���9����^�5�r��h\P>�Nu�� ��
�>2�1�Cew�h�3i���uA�G�~>.�.�;1}Q�u���5�CgR�'G`S �yHw����[���Iw�����i�Y��%�G�۞i��dq>�)��7W*Dr437ҏ�y*�S%<�*�+�;rp��<"z��f7b.\��zɲ�z��}BT�6tċ<n�z�.���:;�J>��!#��-�1S����Bo8`�	��h^���q������S�k�d����O����}����z:{ļ$+ӧ���g�B�q������w��tɥ9k�/�Os]��p�@Ǳc]Z=ISS����ݩ�YQk0ʩC߷�(p�z��w��#���?~�\�c;���r�y�e�{�%�2܀a1����"�6.㘩�z^i�u����'ƌ7kGaw��+�J��������Ŷ/�gO±�qF����8W����L�����IL^����\1ysΊv�<,1�=���:�c� ��?���m�s�y�uj
��[�B��>�}��'غ�4��I��'p���=o���F��0,]	�c�E8�y�8L�Ɵ��OD��~����n���X1��ң|�4��5�^�œ&�<�D� �y�D���m�Z�l�2���La�����h����$p(HM����0�wTړ�g�HT��8^	�><�g��#سy3�y����/݁Kv��E����d�CYX�׮4�+\�J��>E��Ԟ���J�:��p�y�mx������{ذ���Y8�5�g�k�n��Ju�sG��HȐ����p�%\��������ZI����ƌ{��ȏ�Y.���A���_������qfv�����}�X�(>6R �)}�{ze�x[����˸i���R?e���E�E.}�rn�
�R�d�|�9e�� /RbdT��HKc�^F7)'��E4�K�)A;���<�i�a2NO����B ��Q�Eu靚�����DL�Q7�Ԅ��;�=� ���1�f�y�'u�$�,lfrhR���y=]a�T��UR�NBk��d��r�c�͟�bR�{�}�Z�T�^rl^�\�N����D&^�ux�9|�1��8#�W�Ai�K!��lq���?���ï�?�ַ�yI��a7H�1YXy@Np�t�Czz���~bǴ�#�3<*|_�	rT��b���u�u��-{���g�{�>���}VzΩ��åJ'Q�c-O͝�B;9hǍ�4'k���Zŷu(�<m�c��b
���R]�d>�Ks4rح2���kM�p��s|2W%H7��H��su���� �-G��N h�&���x��q�Cuq�&L��ݤ��\.3���I��<"Cv�DO�˘68Zu��T6G������\\��	o��n��O*}|q�/D8c<�!��ݔkhpډ��3Va6���k"3�DN_�P8y�e��Zܩ#�9���;kD\N?"^C��}��Q�ML�3��Km��P'�S��Ҧ��ĳXbĿ���N1e�E���X��˙�f�OM��&�i:�m�Ef�Kf�_�&�G��:Yc�^�w�9�xP2�D�'�9O������ð5�Ōے���^�yYn�4q{E����@X�'�S��H;�c^�l��!��rE9�o��.~�Ml�������o�v+�z�~l۰��r<����!���W9��_�)k���e�	|3Z'O��������[��{/����%S� \H�5H�;`����_���|#���}�Xa�9"�t��H8�����G�I���Cq[��69��@M���_3ֹ�`�o��Rb�V�S8��tNH>'�s�nͥL����q?����]�}���<�����m�\�"��#VL]�1�w>t7��5C�����*��m����=�{Nx�l�C.���*EI�B��J��ʏC7�V6�i9�s����G���o��n�W^x�]�#�֤1B�4�zsG�G;~���vO{ ��
a8iI�Tp�)�����_�5��ǟ�s�GX��UF��v��6�)��W8R�n1Σ��hA̐�d>�&����g��fɅϤ�)x�k������'�<I�ΐ���>/=�#�D"3���������;O�6��YD�ͧ^GϗI!jj_N�A5�uE���8o��(��ڋv/���p\��%m}(��y��G۪j��r�4g�� jr�ϲ�a���L)�!�k��UILg6Ð�9]���9z��D�>U�Dylr,�����n�>!�'�fr(͍�Oo�,��k�9�b���C�$�<G�8Yz} ��2���AIEQ�H��:]
����������G�����\��
�����26���B;�0�ᱴ����\կ5�6bl1`�N T���X������տo�z#:�~��<��Q����//A,.��*-R��?��:����S8�i��rb��i8��+����%%�z���;�՘[G�
��a2:N�hb�E@���P��\esβ��8��0����ޮ�c��'��'	��P��R��}C�|F´sg2��)ģ[�=�h�˝NV���SC�z�������;mĺ4���Sģ��	��4���kݘ̅tWiq�,dm�M�8�]a��"��ju�Z�.�贀x�q-B:^枊0O^�i���9��̋��0N^/K���3(���t��<-/J�l��l�A�T�o[/�(�)a4��ڎ]b�0�f�|�̡W^9��.i�g�t����8 �g�$�IG�j����L��g�̊_q���g
���
{J�-��VJސ+��Z���JYT閆8�!�;�!��wq�����y+��o.�~.6i�sJ�r������ۏp����u�����P፵UlZX���~3�����j�p����c�4�7�{�חc�t�do}�_t���KX��p���\���Aq=���wuٝ���m�hR�ҷ�|F;�	N�`�\�L����qG��p��.{;�'�	8>jb�	��ב䛫!AɘK8Ѽ��q�#�@�
��K"!��M�.�KO���"��%��1�4Ų����X�F��Ӱ�bȅ*�7�P��o�v Bӥ�V́�W�]Z�[ �g?���a�ڼ�^~n۳W_p�۶���lI��|3 �;p��(�ԗ��}�ʶs���̡WM�#
��!<0wo��J��W�};�.
�H�������.�����"[Ł*��m�q�ػ{J����H���UJ���\W����ĥI�q?φ���x�o�BE������N���;hx�1E�}���S�����Ȃ������=Ή��,��6�S �ұ�Z]H6��kc<#��%���R��:3c�[ܩ�paVV��"�M�B&���Ry�����&��]���������$�;�r;���R��&��r���>?G2���zH[yuL��$U8��L���1���Y7����L�l
�(!�Tb��?�{�;>���j�	eX��(]Aɣ�ņ�l܌?�e<���w�έ7���*.�r.�3���D�2���8�p�~ڕs̭��B{"ย���n\���v�y�ux�ͷ�ȁ���_���}��"N�씓֡|<UIV�QC}��9C�bFX�I\Ohzʊ.ͼ�@�O� ~U���0����=�6��iq�/r'�t��l��m�� zGGn�8�&��xz��Ќ}W��]m�<X�EN������o��Y/�c�.�&-c�:S[����E~���nGb���A��Az��+�o��0�_�t�����@��\@U�dH^�T��W��]���~�_��!�K�N&,$H^Q��˲��"����	^4�1C!{>�ߥH�O��SȬ�>�A�S�K+���"j_���G���9�>m������I�n�_ӍY��5�"0
0�1�o��φ��J:���`�O����`�c���`
�N}�h�>��X��"�$l'BY�L�t��!̩��x��)���8��'p��sqǮKq�U����_����T��H�)
V��^����9�f���0JsŤ�K{���m����ҙ����!��r'
w*p�t�L�Aֿ���@ȘR���Ǥ0L8����%D�ùi0���!�͙�ޥ��!Q��
��CCJAcJ���5����''m̸�(��W�LT&�1�ɇ�8���S��ދ����0�SO���>u������0�G���*�jR�Ҥ�ǝ��� ���[�IO;N�9�K�	�q�ؙ��8��<�,4R"i^'��9� ;E��n�whS�B��\p�f��u�[;c!*�=,0x���{'��;�a�g�T@b+��jܳ/.;�<lXZB16���LXݍΆYx���n |����q�ƧO+�n�r]�:�)�6�2D�m�'q��w*��a.K�;P��nS�������i0�Ź�B�dF9�`�}�� �Pd�O�^�f:�}�������8\�������-��[uu)��2�z0�&)��5��o\F��hn����ڹ��بH�ԎPg�s�G8M�>�ڕ#ٮQ��e5)2���6�PAy���AW��QG�o�L�xZ\���� ]u/�L�ڲm8��Q�A�������㱥�l���3�Yj����Jb.^�
q&3��1-M$�@}Y��.��$B'$
�,�����-��|y���9ǝ��j��xZ#�y�1�YiR��������&D�1A�x�Z��ŉf���9��:�@uH�V��J��Ӗ��$K]�� n���g��	�� 51 ��}y�U��#r�J7X�@]O2�8g	oW���c��ϟz�\}~��/��K/��Ҳ>QO�V3�|��Q���GFF/|-�dFO7a�����'�*�*�/��.؉���]8��1<�������ko���1>�╋�*�!N�$���+���)�.;ҫTy�JI2W���iO9��J'����Qw�<�>���F�cc��X��~�t*)/C��4�U���<v�"a�p�#���s�u<�֟ 7��"h�搒c]yX
c��S8���_�`��k�ܢ(�1%ԐF֕��D�m��/�A�p�=�7���q��ڰI/���*Gx"��S��Q��ykY����v��u�o��:�*ꇔ����S�<��$�40�'�G,(�'����)��Xn�9Oc|�<A(�lN4愰Sļ�^B:<ߌ��]������"�U+�.����^�q}`�\��r�=�&�Bǵ	{��C$"�Lh�!nE���w�m�j����<b=$�/���e�,-(�h��	%�a1L��h�̉m�&M��6ɓ��H�3s�S2.G~��� �r-d<κ���^>��y�4�'�)���f9���w�����y�������1,���S�ݨbta��5���5�4'�I�\,p��/�?�˯~��^=�?�n��"�{�5����8o�6,ca��Sa�����S��l���W,ش<Dy�$����E
��cʑ�*�K����5��X ��,=d�zW���MẑQ$yD���z<�b�V���&OH6q{X�m.�I5�����J�%iy���� G���;u_x:%uQ`��4N�� z�~�X&g"��Qs��8h)`�z"��!7y~�_N�7�\e�<}`����rt�"�FA� �D�ǵ{g�&�Lxv�O�h`�1rJ�ė~��t7K�]]K��%(-P 1e�1_� Y����+I�}Q`���J~/.��x�G>:�_��1����_�߸�Fܵo�߱ŨR��+rd�|R;�o�[�UsA���/]=�d�4^y�],We�%��pmN>�	:&�	OW_	|�K�D�QK�.|N ��d�}�O����Cgo��c)��&$�!��1/�3�����G�(�Ǒ)��B-j�[�d���f�%��8/�2�Y��%s`�)��$�m�+UV\R��/8�"H��~Sz6�D04t��'J��?�熟�v���5�D�����F/K_��ҥ5�=�]W2���+znW銢pK�d���HM����Ze�8�g�V�����׉T&����h�z��鑍o�s7HS/�̳�3��w4[��M�[�yO���M�K�>
j[�)��ld�!!2�� �k�*�<ftu?�.���cH��_�0o���=��g7Br�{�Y)�&�=~�
Gs�>��H���zhkOw�$=-�sJ�6B(~�8���%���#��ï��];q�W��}Wc�[��T)�KsО��5$|,`=��'k�W��*D*���ί�W|å�K������8��[x����^��G�'Nae���S՜_����;b����4�')��p��Ķ$[���:�� �Nv?5ow'sRPCظN߰r����G]Q��&�8!�$�C)"����#%��%c��:3�:]�׳k��.ҔO�b�2�a�لp\�Y.��N�eqG*����.�[�gm?)9Ѷ�&��/����[�_�a.\���;,�ak��-Q�B�ϩ�@����a��c\�u=�p혳���[~|C��g4�K��dX���E2�k��ʄ+��R��z�(��5az�q�1_��RǨ|��9ĩ���J-�M��ԥu�F��K0�i��or$��[�=[V̖�	g���Av|�h^��5��Ʈ�;�����s��/v��ʝ$��
C4���d28>N��Μz�C�@U�2��1��taR���6�Y�C�qT�{.�(�|Ƶ��]j�3�T2�[H��`�=���N�X+G+���
��k�㾗��%߿_�}�y�M�e���|�F�ӕ3R��=�NAѢ���v�mU��;|��ኡE��ªlz�$Wݕ)�.�v�X���>"���KFz!�"F=�\�qX��+�w4,ܐ��wN��eM�}�������i���h�+^=e�*�	���9��Ɋ��q*�3
)�y�G�r�1�i,��1�	�P�&�
��Y������)��9M�.m�b0m(0�L&�qŔ+aD���2����+�i�']iR5
舫UAc�Sؿ�e����
�R�]����#]�+��*��o�F��ѣ���ױ���K.�G|�q�ո��-��=?�6	w��]�1��[�p��c,-X��P�g.��dt ��)��Z�.c+]���?x��%7�8E�?���>~L4����9��#�a���s�ɬXD���k��L׶��y�����^��2�}M���5�|�q>=N7�J�7f�?� C���RJ�e|���B�J+m9Γ��Jrw����.=�3�B��Έ��a�U6/sá�9,{��0�)���H���u-�2x��0E,R3�6�|�R�et�n|�ɖw��'�鹝S�R��Y��Fֳ!x�[\�9�K)�q�rVk���F��3�|eh��=U_�Y_绹�����?�?|(�n -
W����\:ư;}�3�@`$�QI�?~� �Ó�s�
�j7�س�/��^x>6hG���{N��1"��\1��􇕛�H{��8]l)����K�k�]�N|�'^}|�����+�*��Ir�0F(�[4�K�9�>K��cR�6RG#��x�aHa�/����^M�g��P$yAE%��(%��٧��`11�;�y���CDTGC?F9�ܜ0�ب�i]��%Ҹ�-����V����(0�s}E�Q�g��@l/H�0>f����4�77E���e�Our�bU��"X\�R^G�J_`,�n|u�9��I�,���%�'��Fp̱�k]��_�v9}'��������:�U���N�I��̰j�q�{��y��y��Ȼ�(V<dû��ʕs�i�o
�p���g5�5�*Ĩ%���_S�i���^���C
[����	�s�N	BB�#K�#�g9�F�,�;G��.���5�������|,d�~�xb�i���Rڋ��u�*��4��`
{܁��I��o}�J��PbmP���iy� ���A�ٱ7]z	���
�t�s7.W��M�F���U���9�#���x��EU��ie��͠,�F�n��}����A7�[3���YDI���t��H���D�f}�l�u~֑.�̏^��a���+���4���tV�֊��f?�l(�-aB��mNh�3d��	�,��c^! 3Q���NW
�'C�i�h���?���Y&����T���I������Y:���]0�a����o��/�کcia����U��O�ơg�ϟ}������Ҟ+q��;��4X�>�U�lKC����n+�B{���ǿ����zV}�q�|��%bC�A�[נ�f��o�����&���E�&[�]HڕW/%��f�-8GF�Y�����<L�+�5�X�C��d$a|}��>� ���da�?��v�;����/���A��(H�>g��i��-���xh\��W�s��H��qɞp�w�J0��AK �9DxLy�0C��VLZ�O�AKtQxS;3�#�4�a�)fM��#��� o���]�P��+T~\��~�ZD�:@���WF�"z�DgK⬚��R�,�=]B^���Z6���˛R��s��d���w�P��W�C�g�u�myfu�h��QS����<����`.^���E�7�R��j��Ǯ��s$>��0�qA��0I��tUJ,X^ނU�p�z����GO����y��;o�mW_��n�P�_�T��|WW7��^���}=A��P'l�A�08��]j�\�wU9]��eqw_�_��||�8���F�DK�{,�B�(��5u:�"�ެI�*I�m�8��tH���E�(��s��H[_�w2	���8\,{��ON�����g�N�i��� &�Pc�I��⅖Y�.;���Y��V�0� �>W(�g!,��qڸM���sv��.�������Y,���z9, Й�桬����zO�9&"Cz9͂x��τ�u�Ln��� k���z+&6��U��T����ߠ .W�r��Ts���]� �h�m���Yٜ�u^翇z������*2��s��2��C�g!@��B�@��k���<R���T>*Й�0���f�9��|��<��i�4����4'�Uxi��U[{0'D�ݳ��Zr�i�rm��%���V�?s3�� W�-�z����z�ťJ����٣�}�G�8���� �ܾ_�n~m�����ui�J/�H�Ƕ�t��r%)�ݱ����G�O�pe�^���:Sz+�dxB�v{j�-�kuha��1������^�?���s��)��W��$��az�z]���^n
t)�ڴ�f��M����il�������.�k��@��ȁ�7۳��O�Khsb���~=,����r3�k>b"�;k>�1��]�rW���������j���Q(IN#lf@9R�"�1Z$���_���-��<��,h��R� ���Pi���	}��#�|�8���|�׏�e7�k��⛷ތ}��֭��3?0Z�q?�l���XX��w?�?��9���
�>��^& ���<Ie��gS�J+�}s�,v�Ttt3oC~w�r
;�K�8!$윁ܽ��	vS$�:~����$2A����,�3m$7���cK/88L���!ղv���{����^?$H	�oh�x|��.�?�4���W�	4}��o��ᅱ��@898��X��n�!�O[�����W�t�y���U��i#axh)�����'l�2��`d���̸��Ei�_����p�Il�%�ϒ�;V��8%9OX��"����@p��e'�����"OLB�u��u�w�>6jA6��$����}QJ.{�_Է�']���'�O�언1���I]�C��.b��8e�>SmG��EB����)��k���1�/��3�,B�o]Cm�wH�ی��
�:��*��m^���BJ���'Ux��RFNѾ�,7�I'0��|7l������ϕ۵��Jm܈_����.����G\�an�y��n��
����K+�0<'�u!��'�d�[O��a�9�"ދb �����Y�FeL��R�$�JV���h��Q�dvi�L���d��YldD��<��+$�\�?�-^�~�ma/!p�IhA9!����vxs�Q�ev��#����tU�{��!��uc�'Ϭ�EvA��&n$m*���Q/�
��ϟ8�ˁ���m
���J酕��i�&ׁY�I�E.>�>�a��r Y?��J��ٹq�R&�=�q^���{�v�4|��28����3'�G�:�U���5����6R,Okv��u%�,�&Ǖ��]ȴ��,���#�X�d.-�2��'\Zڼ�e����u\�4�ϯ\�Z���|<���S:d�Оg����=Yq���@Z���%���>L�ڔe��]���b(v��<4�6gL�����e��;�@�&�w�r��-��LU�'q�b�<�1E������R�gv���4�ޅ������-9�t^�����ĵ4���%RD��h}�-T�SЍD0�2�ҭ욌�Y[��� �w�gɕ%��&��;���6��k/؆oݺ�ҵ�ť[6c㖭k���v>CS݅%<��K�����8x�$������"&q��W�����Q������;�:nC���X��%Ŗ�{Nkj��O�#.u��3!�6��<l[�M�>���)�o$��(1�����$òS��mo�!�MhͿfw-�&���ˁ����~��K�V�fbǍY��4L��*e�)�M��23�=S��;
fg��20��B{ӑځg�g��OgH�Sm�9�)�WHS;�Q;�Ӯ<z͔���B�l�;@�ˑ�Ì�Ӓ	�D+��v����vC�K�d]^܀U,�*���y��sصyn�l'��z��y)���Iu$�����'�/�O��0�z�ZZŘ��Y�Jyiwy9p$�0/n����Z���]h���!�#��.}|�ȿ������ne���;��i�3_�L���~��EB�5��+dzVrz����/��������qxw�N��P�'A��_[ࣱģ� �K��q�i�u	�R(��K>wlLϦlz��s�;z���� 7~�/X��F}��_%@k�X/��*�6^�F͊���`�uyKK����)�\[�h\�,T��r_�Y�}f����1��$(g�]Z�з�Y���aAJR��.°�����0h�ZJ�]�w�8��D�RD�)�U�)ׅ��8I5lR��&�{L�I���ws
T���@eY{�2d�p�C*�I可��]:ƂZ�8��_2�����P�Zb9_O�e��Q+�'YfH���YJ^��-F���in�i|t5 L�0 �%ї��*���Dm�d���UXȃao����-쏥я��Rφc*�5XT���/�|�{�E\��_�r'�z�>�>�]\�P���;kӮ	]t�hX֨N��6���j��J��p���N)�Ufn�ٺ��F՗Q%��S�N+�Lh�2���}��~�VN�������6��rcT�.�h�I����2�:�Gm�-�nçgO���_�E�r�Z�З�����ʩ��}�K���u���	��Q'�"�o
�t�Q^?o�=H��Ffr�@N��0��R|��Q3g�n[���C� �h!��8��E]g����6yҜ�<ܴ���@��b��0wL:��� l'�&�D	�G��Qi]��k�ߑqJkkcl,�u�F=�?>}
�NW�u��'1����|�G�r"Ty*��fͨz?� zQ� ��zЬM1^�fk�t�
������~��m,Qoe�e]_�.�z�V�e��Ǔ��M#?֡z�X��O��ks��e��4v���ş�i�˙�+����S��q��:�4fC�YK*�o�|0���$.;���gNO��M����I�͢0���M��X�Sx�f'k��7O�8J&�V��@(�5��/q��K1�S"�*��=��.��ث+��"�tu���e�OY��Z#����98]ͭG+���O�?��A\w�ܹg7��z�ڱ6,=m0������<� ��O�k�������k0�[t��x��[k_��7��!l:�🔲�ǫ���̂����ޓ��;U�2S5��^�'���g�Є�s�nsx�>�`mӂ���磣��1�z[�������i�*/�֟V9��wA��h��u�B��6�}�`�}2�m��β�o�x��Bk19-%�ی�C�l�
�cK��&�\�#��D3��
�jP��]fO�D�]R��(_��^!
�Vϟ�d���<��<}�o>�w^���?K���ٓ��׏��� ㅡY�T�zi,��^|�ÒhLYָb\"ՙ�>Ӕ���tS�U`L!��[C�kD���9u�����z�
���熸Y-ص)�i�  ��5t=�IZc��%F��}�G��n:�U@�@��Ƒǖ����l��_Fς��@���.�~v���7��1��拷��ة|����[,���A�ٌ����k;V�p�R�V�M��g�&�{�͸��k��8��k�8x�<t�0z�=�	ֆK�,,(�NbM�����4�mhL�cʥ����c�L�/���x'5j��b'�{��U����87�}���9r������6�g���X�L0uSv�Y��R�	�J�����Ay�^�E�I�Ǒ�|L�es��d�tx%5o�X�0��I����š�SG*}�؞*#.�:�|�h��`�`��$8��wqA���D|�}�.¥	������t�s���^v�Z���TW"��8w+�;���X���I<����}{�o·�ߋo޲����ӣqՁ�L�kS� �ө��+�%�r�Hv}�5�y&�F��3u|�r�K�V�	��PK�������m,]ea���tm0q����-�'SW��󡚝(��yTE�F��`v������p�ӘK��8����vxŋ�j������P-'GN&<���r��;E����or"�yV���a��EsZӕ�o�r)yz0��}���OO|;���c@n̥�o�F�L�@�mfqm�t7��F-��F��s�T���J��K.ǽ7߆+.�k�N��G�#/��g��So��+���e�C�G���\ɛ�ڂ�\)-�2��v2��ӡ���j_���N	yg
�Ũ0~'j��E�P'�F��:ey��g�ԘY�Yr��Z䞥��Q��A���α�OQ�x�F9��X�u�I�MJ�ɽ��-�M�̡�X��k�-�L��(ǫ�B̑�t�\l�:�'������mz��WiqCaO�+-Y�]�Z#)�sFQqb\��wO��7ǿx�q\�mnؽ۷lպ�_��x���,bTt�B�5����.^��6����VM�"�a{$��H0�鰕tW�yD������/���=�}�r;-�+�B{�?q?��J����2����+��]�_=�Z�C
B/�}��y�e���{�I����6F�r�Qۋ�C �P,�Z+�� �b�"�l**ύ�����Ο��'+�t�}Gi��e5e鏺�p@�K$F�E<{�$�|�9,x�+��R�ag��>�(�KEɱ��-�R���x���M�F�7��/�w�D������q�R�<t+����g���igm8M����}�%'6y��u���32��'��g'��a��c�����9k�'�ǝ6����>����K�;ଂu*+2V��d�ǧ�U�����*W#,�Wq�"�_��=���8��m0��R_+u�����_���!=�<���Oౣo��1ؼ�ǑޡV)da�[��o`w�ԩ�HCɎ�.�ƌ�N�t<ɵ�KΈ���;5�#�e��]��3����A.m!�$������	�r,�9�X����]v|ZB��9���yd2ik�(z6��\ �;^&6V�ȸ�'�D<˸�E=��NUdF)�.���C�\'2��N\�VD�p���c�N��1R������e�,��ɓ8�Ӈ���1�p�|��]���+�g�Eذ\ɾUi�mV	�.���0�㵗�;�`�"�7�nQ����jѸ�K+���K/�5�<�g�x'Ԗ��₾�Q]!���Ѳ^9��"��REQ���+����d"�Iŀ7%�2	Z��)V�
����V�ga1C��9i䝝��u����D�A0�LzQJ��K�9���|��vl���|9L��гMM<8�۹)�k�5Ec�,���iu�;�y�N�<�a:OMǴ�"P����h����!P����f8g2��H�X~
��R���O}��T�������˱8X1���{/��������ţ��'���~����#|�V��}���j��^Y�E��=%S�{u*��DW�t\��k��-��[��";n��"��tA������]��SV�&��i�N<�SJI����g��Y�7��0#��2�W��8�o���9S��m��󨵉;�J��2�ph�u���j,�#�T5j\��0�r=�'\R�:�rx-�ӷ[�1�6��sU����8��5�P,���g��~+j%��s\}��j{�:K��3,��K걋ʻ�Z^��y�=I���S�#�A�\�	��d�^���(�y!������Z�Y�#p�F���w=|�ڱӅ��� �)�Ѩ 9!Y�ؐ?��UK����'pHu�vtﴁ3������D·X��L���Sj��t	|E�T��#"�'�n���d��V�$�ќ�G����Б֥����8����ۀ���0U��`�:��, ��Fio�6�����鲔P���=BCJ:�i��
D,.U a�� ��R�U���ύZB�>yZ1��cN�Q��mC�$�c8}-�N�(6��Y;
[7�)��5A�.�O$�ӈ�8Gt�$�����ΒN�S�)��7w�6v�w2p�K�	.)E�&(U�0���|�?����4��\����w&�%�����Zo��ٓ�3 S�����Vf0���0VN�:>���U�3�4G��:q�p���n�}����*�]Q�e�,q���[�ތ��|#�x��x�ŗ�����^��k�xa�+��QC]a��S�Y8R�Ne���0������%��V�Ld���c�Zbё�����>F}���~���ta��pɿDl!5Ze��^Af>�gSL�9d���9ŵ�I�$���gbGtn1�O��)Oh��\QH2����1Z��Q�Qpeì�-
�Q�Nb���֧�tM��W��'�kb��yȊ�dût��9�����>�������A��x���Ј;a��X�)U�b�Ӌx�j���.�?���O��]�����]W]����*?�.R��|>�<��F:Yؓ7� E�Le�����Ұ��o�	7\y�r���~~�^|�=�85�hq���7G�K#����m�Ի��O�"�b��K�c�ku +�]���&9}��Q�yK]z�o�x]�y,����g�5������	����7r�uV�}]��/$�=o���d�sv�T<'>�(��4���m��L���x'*\��@��{�>�y����1�`yQ6��`S^և�21�=����	c��hU����o���w�m�T�7��	�f�+�='%�+�y�%b��K���v7�{镊�����y�~T��./�
�Σؿ��R]�Rg�	P���^pz�E�Q/=O���Q{%�������k3"��O0�|�dOr��n2�?�E�����t0]�]_Q�l��|b��8+�C7��<}h�[�.c;'���&�̿3����R�I��yt:a�e-�LA�g<č��R$Z.�o�����$�;��,F�V��g�B��urT����C�d��`J�S`���p���M�Vk0rh텅sQ���D�
��]l})˯E�I|K��&�R>��CD�z��D*k�M<��8�y�Oˣ&M_���&g���i���Y��I2[��	Ɨf	bd��άd����ρCuH!�6D�b�5�����0�'V�y�i�Dp�����v��ӆ �9�դ��7�߇�iB�0"�g85s��5ϫ`�tV x��'k��д(�R�ü-��q~<B �����Ŵ�b�*��\��|����θ��S@|e��7�X�9�K}�;(TDm�\3�*ԡ���.)p0�۝�2(��vaON��G�&�HU�������@�X���"#�B��+]�́��B���/��w5�I͚���w�/���6y��+,�`���3ja�v�X���z�к��h�3P&�^�P�y�D����c)jS01��R%��Ԯ�d]���ق�ٖ��RD�8�Nb�c�c���������<m<E�FfF���Mc�kk��o~�\q����P�=a|�)�j�Ĳ`��b�΋�w�/�}�z?9�>�*�S�vq���v����E���;��Q��8�I��Cg��#ߩ���IN|)��zs��|��	��"�G���H�ݦ '|�;PuR�3�jڐSیB|^��Y��.�MZf[:�������"37��۝�e�--8��B�6s��lG��#�x��>� H_
����ӘoFI�,���r�<���h�+�K���g 2��$X�v'�de�pm��a�U�������G���K�uj�P0ҲKb��T>�T`����G�}?:���#|e�n��m7�k��0�MJW(-A����X�m��b�� `u����Sؾ����݋�^�ﯞ�C�/z?;�
�<����t�K��̗z+��@�8���L�fw�9�����Λ �
�Ҿ�f�#=���ǣ�f���N�sP�Ō٫�V�p�t��&���E2�;r��]B
���}��:��3B�D�Hǈe �}�}i}���Zc�Δ��d�Ҵ�ޡ��A��I#�%�9��Ϛ~�gt�\����'p����۾����"t�r��M����;�mb>�?٘�Z�V;��x>�?.M�Gkغa�~��aX=��D{	� ��g�T!�-�
�ܻ��ۋ?��]x���q������ٷ�ǉ�%��XVȨc�����
�C��䄪SaǕ�:��w�b������1Vp���L�@�`��*��}��$�c��;C�	�X�!���؀�b�y�C�غ>����	�'��Iv���i��)�d���?󰻥�c-}�lKӉp��\2�\�c�m�jQD"^��{�F���/ǩ&�����u�Μ>EN�{�A�v �=R����-r�=+z�nE�H^.��)8)����q�H��k �����D��М�'�4z\PGKӇܚj*ޤ�ȧe����S?Q R�\ZD�D�f;�}�6$�&'�	�7L��v%[��]���^	Su���I�ӁĤF]'����d�4�k��s�;W��T䆨�K�cl;�DJ.#e��ϕ����sڭ0�dN-��2����jc,)'��;��y�H��3�p�r��(w�عФ�dt�th"Bd���s$�6v)z<?#E��EF��b'�tR�c�F'u�|K���^S��I�\26�Z�K�.l�GY����`��)�MAo_q�X(�e!�r�陼O"HO���m����K��)��I	J7�◭hX�1��u�%��d1��wI�#M�e\���=��CI�d��9������Mc����i��|��	岕Q���D�T�.{Q�CL>�o���㊺�r���U���D�E��5�˶m�7o���!F-�(�y�n`�����c3N+���������;o��/��?�:�?ykK�/z��B��J�OB��v}��f��c���� �!�C*]��O��/�#�#"���ȴs����LB��ð5����.Nv9^�����)��!M��a�se��l��a��#)�|t���пgR���hw�p���)B��2������7�����7ɴzMN^��F��Y���0T}�_
Lٱ��w�'�)�4��s�q����v�kHJ6���K�i[�^����$e2 �؈��%�'��GG^�_<�vnX½7��=�ތ�w^��K:�rU���@�J��k��h�e�]ۚ��dz�I2FOCri�
l^\ƽ���k��[�?�O�z��a<��8���b�&,s���1�w(L4F����`�H�H�2���c�؃X���ƫ��H�,�+�9�D��Dt}�`�P(#�zD��J`���4������X�T���Kere/nPٯң\��=Le	�����9[T��*�k#���g�����F���s�:Ф�"7v�hl3w��0��7�`�u27�:�(W���vC���*��aJ!]=�"��ԫ��ݽ�r�ܱ�6yl��0+��^�V�	sa��Ͽ�
��5��_���~�	|���p��qB�ъ��k�F�.�PYZ~����/��*I'��E�y��L��>�7���vd�߆�DH�<���\u$Hm2�̳�C\o:ی^��&0Z<�Sq����,��H5���K��iZ9e�����I�4���ɧ�Ʈ�m�z˗8v/���%Sr�@D��i�˽��8P���\=��Xz��h��x>1_o��o���@z��y�)�Wګ#��y����S6H�q�a���8�z^ej���x8�:�xTw�qkk0q�0�D\.��vk�릹��s����ՠ�cV��s�t������4"���	��u<(�=�L���F_��z� k�	�+��W���`A탤˳�5�}V�J��I�*M������Z�k�3��H�����bqx��������l�����9���>�,!�D�&�����$� >EZ)����t�	��ah��N>���y���;�`���iCmW�Fq��Č���-�\/D���d <W�t�jQ]�Ȯ�������������q$���-|�?>]z��]�	M�O��W)
�X|��fJ�j3��K���[�A���������R��	ϴѠq|q��y��"��֔7��q�����67�3�½a7GU��xT�/j�¼��2 }�!̉-��{��v,-�k��ʒ'�=��Z��;m|,�԰2z$�ea~��[�������O��Y<�ڛ�`�$�A9su|� ���Y ЕT%�h��)�aN$�=��1�H9N	�J�;y�]k������A+�e{,������<�?Y�ySVM���w�<��k���ě��g�SDY��Q�K���B�:�!Y����f�m�S��;�r���K������l��������5d9'~��{�D�#�1j+a���}J���:��NEA{s��������ɱ.Cǿ�a���82��x� ���+ػm+~��+p�+p�y����*��Y��a�.{��~��9a�,���R#��+�����qBQ�h���Jv_�u3.��|����[��d�����z��:�cP�X�+ �5+cs(�q�E�UkO�7�C��us/�{3�/����˗N��tQ����)� �y����k�pN��Lg� �C�.����3�kna���z/)Y���;��\8�ԏ���Gw�bJ!}��$��If��1�P�}�e�>?��� �"�ֵ�Bʹ|ǌ۱�+O�s�e�#�-S���	?�˜��_K�^���0*�{�q�o\����{p����_<��?�"^z�]�*Ug��y��%NۘF�݇�u�:1Y5o晹�ʔ�[��[��vÑ��"�5A�۶��Ө�m�Q�~ZӴ=�rkX�IkS���\m�R�q�H�m=����L�w|ή@�]-��+�˞��<O״��7pG�X;��a���<��[d�[rIs�]�[[$N0F��Sw��e�H�M�TNS{r���W֒��`2܊[�n�`��s�O�Q��Rg30m����!�׀s��4K��o�ѻT��$��-����+� ,$�>�������GR�t��t(��}���N3	Ԅ]���%���p�|���A�;�_�v�'Jɳ"�.z�w�9���LmHh+y�b�+�*�#ST
 D�&�uQ���uJ���6pC�ڰ���j'�YJ����>�E�p�@�2�ay��EHy.���N]1��yP�0�6�8�B���:}0]}7�>�՝� �w��Q�ݱK��K�eBH�5r� ��Ww��6���3[��[��]<��)�"H�Jք|�7p8�ن���z.ܴ���ޗ7��Y�h�Jʤ3"�'0O^!���҃�T69~۶kl=C���1�|ta):Oiy�}���-f8݅Ύ��(w�H�#�Z�x
�i�9"̜*+|ǀ�
�[[[���l�PE,U�U<��(�['����9d&�n�*�hU|��s�}�V�旮�ﾇG���~�9<���x{�����Á.C�7)�:�rN;q�V�dt�M�w�E�A]�����X��渽��d�J��E<��މ�r<S�eF|����n!�yUS��Mܘ"�w��XŚ��g�:��d�2��S�v��Te���i�+���7~޶�&vZ�4�D��Avi��5�߱������\Nҕ��A�teg�1򀌷���.e)G�BbQ��2��waK.�\,�\�Cｉ��z?n�y!~c�5�s�n\�};����c���:Q�\�v���E��.�%�0~'�p4�ea��1��H嘩���ō���+����ON��S/�
~o|�N���@,,`4�'����iW]5	{��� .��ε�H<Oe�p�c�|���u�+�-Tg����wB�%ŵ�?i�:^��9�����[�2�<�(Ӵ��T3^4�F��tV҉I�^�oj�3���0:����ii��T�X����s*��!���g�u���_����>�s�e2��/�j�,W�^�y��n����Ӕa���ߍÅ�Ny�ҝ6��i�E�a�����/��K���s����G�q�V�aP�<���#!��*��B��Dw��+�^߾�N|ƹ�E�-Hoe)���F���Q�z��(����i�9�73� �L'H�	�)��m��x��ӂRd�>l-g"�Y͘[�ġb�2�~���#Ȭͩ9dYP'fZbzCI1���6�H������
ŁaL?�V�f�=4�8���ɄŮAݮ�%���v2��Y��uڒ�Q�F�5����B�}\���	��n���A�95�(d�G\�� +�q�Nx�ѼA[zy�2 �Wˀ�C40��������j=�����N|�m�W�N�m�<[>+ҵ/N�ȁ�s��s:���n���b�,@���7����]�����Cl�ڙ&��@7��5pF���#v���|d��^�B��I8a�GBr�*���i�4fR�{�ù��h�Nr����J�Qfe@�Y�5G˒�BIg��R�noY)�li��9CS�3�p8[ѣA����`�T�z(k�L��S��y�1�ƒ����� ���3�Ic���	�y���Y ��bLyO���P�m�/��#~���!�c���/R<�)�З_K��|�)�3m\�u眝P����G`���F�:�n�:~ SyD��5��JL�l����brj���O@*-i�GZ5�YQ~�x�	n��GЫo���Gܲ�|��b|��/�#/�O=�<��>>����j�����p�K��9g������lZ�#�e�Xa��_�K2߀�a=�ߔ얏�����)�PA�G��:�f��}�hٓ�3j�%ę�Ksa�ƃ����7'HmL�İ�H7_M'[�Լ�s�n-ֈ26��~�O�3/DX%)��p؉-���Ɖ�!�4!J���Z����˱>�	ry������7G~�K6<�;w��ߺm?n��
l>g	���J9��Lj�H%/K#[����cl~ޡ��UHm��Z�:��\�v�Tu����~�>|��}x����:�����^�1�Uy-/�0cP(�[e0W4�드�Y0���K��Hy�mL)W�Xa=C���trZa�$��G�m"�
�[Bf��)"��T?�M���튟�=�K6�/�|���.�'p'����:����Ȋ[��o�^���,Cα�o�5�J3��S�>J?�������",�����6Pl�t���\?�����jψ~�FwE�j���N���%�)�]ߘ��ed�~ @�'QX�L��B�p/Xڄ�܂;�ڋ�������_<�G_oW�~,�(*}Gy�+�G�9Ҟ�ᎁ�,]��,�~�g�(|=�<�����옲y��J��d�{��`�_�1[Le��/��b:j\����x|�Ϭ�٧4�@u�d��yI�mjC�
mv5��.�H��q�9�e��|�z*+�e�����-y��$��x��ӛq�"�%��4�i���"S�$+���``s�؜���1��l��êelfӬrΠ�
պ�����+,�&+�1��Wz�p8Л�
�Yl�N�3y ��Ɲ6���h�T̫)%�ْ�j��P��N&!�`��D��{1��ʛ:��>��)<X��2(7��ڃ�ŕ&�vT�8��tw�W8��J���6$�m2����;pH6�mkq�� j�E#�A빘ĝ7����?xp���'1��n�R3��<	�l+?��Jmc���dD������-�k�� �܋8�.��<sQ�m%Ȩ*Hy�>��1ADG���i@$��x$ũrM�`��0.�(R��S�2��I'ƌQUJ�VZY����n�<X����6V��%*!q��'��!VW�9=Ҋ��X�n��=�C�qʀ�&#1�X_'{��/��$�vO��|ҷ1*'��뷵I�{�s�w��)�]@AjG�3�'��d�0���N�z��Q�:G���]L��\�'���X��,����
6��G�d�q�_w�;�B|_]-��#7���b_���D��gئ�,�v�M��M�1GQ=�t
��W��eO�ta�Qb�CG���ذ�X�BIB�y�B�.�1ņ6�H�;�:\�ӊ���j�i4�9���]���=����^~��'�Ᵽ��ON�ܸX��+UT�r��*��@��a!8��y�{#�4��>�� ��7���3㩾}"�*)���+p�,>B���j��FO�pcճ��$�4ޱӍ.�;ןN��cXn�F�6�Q�q�����k�k����i,7�o�1s��s�,4`?��]��}U���$����,6�/|<&�5���s<����w��=�o��Kmb4��6jaN��ׁU����"^�ƫ��{�Õ��ō�\��\�7�ݍmW���2\�+�)$-�>f����h��m* �fQ�x9No���^X&!פ>d���{ǝ���[�����g�>��x�Y��:�xq��m�seA�4�K!F�}�
g�u�^�}_l��yN!zv:�T�v�i�!A�d�L� �,&K,����m�ץ��:��^�/��5�K����;/d.�Ҡ�f���aF�խ�1�Y���q���t�����+?�C����t���w��,���Ԏ'�Iʄ�Yץ�n�s�o�ЕgJFp�����:�otz�+����Gp�uנ��(�%J{Ph/<��7���L.��k�.L�Ԯኗ_�i���[�w�x^=���O���?��Ç�/��,T|va<�H��S��<D'����q���0��i���ҟ:�?�һ~"�n�RM"'h��m���J�
�P�9c�]�huue̞X`���!�x��0PK�$�&l#�kӰ(mק�Rs���)�>L��@Ά�EF�⤝2�u��A.Ry؅�6<���fυ�s"��N�
L&��E��	#��3��e&�( �q���$����d2v�-�Z!^Cr�c�n�q����7����9NH{-
.���͔(O��8*�Q�1\X�h$�&�85:	�y�
1�W^c��[XYlN�b�MJֵ�N6��Qn�8p/���?2 ��6 xq�4i�c��'��<�S�������������| j 7�X>�oݣ8��43�G�9I2Ty�穴}t�m�Ζر�:LxG�ܹ�F򪒈��6�4����������j'R*蝟l��S&�ML&7���k+���(�b]�2�����0�2�q�<���f9��]��qa�Lzi�A��+|$�C{��ԟ�o+}�e^z)�.L�jvc�VwQ�\Ŧq��v^�{o��^r16�,U����᥷��CO���*e{C�����ڳ6f�&�����
�4[|I�����4d���@��i�$!L�
W�nD=;L����q��[��]_�ϴ͵:~3q�) Z��,d�����䃊�k@<�������l\����C�m#ՔT���!+^w�nH�����Fl�w}>�K6�� ��Q���ZC� ġ�?�����ߺ+���f �C����-h�XWQ�J�*l����xbaT>��zz���}W��W������g�|?~� z��~�|<b��D�N+��v�(*eM؝i�xw�%��vd-�i"�J�c�̋�6��ת�y�˓E�G]zrN�a�� ��~f��A��̎�yݐԯR8O:�	k(ݕ���)S��u!�k���rz�g���E� �5?�O3�ɡ8�P�[���8F�����.�	�hdu1�r���ҜL��8`b�І�rq�r�T�>}�8�z�C�ϼ�]�6�}�p�UW⪋.���e,,���Z�.�X�o)1ND�����d�d�N�������[�߫�X��u�U�q��W���^�?��O��/��'z���U����_9"M-��qI��,�����.nPo�C�`�g�����8��W�<�z>��˧_L;�yR�~ص���܌B0��tn���96n���g2��.����Sg��C�����s/�5H�d7�OJ�0�ϳP5��D\G/1X(0���'��7]��؅b��>��ׇ���/���ɕ]]��,M����3ya�b4�~!��n���{��~���8�&~��Sx��cxo������>�I; F�P7�	�Z���X�VsL�e�m��_��2{�S�x�i=@m��u�Z��2m�Q���_�����ӳ�'�jc2b:��9[Z[��Oۻɂ0��d�����զ�4�q>�d�ec�RV�m s�S���@hE�Xn�V���͞��3�C��l6�O֩���mIϱ��Vv�IZ*�B����9�#G���r�S�q����ݸ�mߊ�ˋX=y����~��<S�pr(����f%�5c�_H6#2��Z��Aj/iFDÊC"����M��� �>���e#8�� ��Ж&No�������s�����= H��i���*p�6�t1�V_�3z9pH�&�e�e���2�ߓ©�K�S^�&��vQ�'L:M��V��X���s��-=���(�ہv	Y�*2i(O+Y�J�̀�{�x��@�3�2�op���?b��s;?�\�@@�<<���QZOk%��i�^����\Q}�����u�������+wa��M��b���2�h;n�v��&��?�1����p\���z�i�ݫ)�0X�l�����uo���� C��1���.���aM�@��hSC>��k���NT#~D;f�yy�RG��� ��̉)�8%!Ag��wj����OUIQS�(�B�(-OJ�̝xBRp���>n�6	������^&
�٬�Pc��kmi���Gp��)��W��U�m�8�j�{��Ps2A���`�0@I
9qY&�T�%�0���/Ş�;�/~���x�#x���x�_�XŏO��^���;Z���f���f�eu�=i�� V�G�V���!�/���X-�x�(T�����y5΁.$�a�{^��Gm�ܤ��/���^A�SV{�X|I9j7)�� h�?��!��Ar�w��]��@�S9�j6�L{�˳ۮ�iCNNuY���75M�gk�̯�/�1�)��� =/��c�Z���6����NZ�f��TEav)Y�Ce��|�qR9K(�Uړ5�4ıJy�����܏�}?�=�\|���}{�k�Vl:w��[T�z�:�@��T�ZB�㇥�Pw�J/�j��Ԑ�q��P`4�JU�o�z���b���'��#GQ�,j�)+�I�B���1l���F�agz1�i�,��\�9������Dwo,�mE0-
���X��Z��v��r�eV|�4�L�]ƌU�/�v$���9�6}�IFq�>Q�th�.22t��NO�z���\�	�etb(�$���%?C݌c���b�qt0'3�x��)����)~��w��;G�}�:2�W'(����y�#�In�F��{/�|_�Vi-j'�8w�9���-�c�U��;n������ƃ/�����G��#��3�t�꿡:�SZYb�b٢��6؏�ۅ--�X��[�e�w ~1Irmǖ�Z\�Gd��<�H��eݘmw=%R�H��z8W�g��;�� �J>�:�Y�5�َ!�=�x�����b\���H���脗t���	�Z���
���Hf&Isl/�4�L��R��Z>�GVnj�@�ʳ�D+i<�<�5�E����X�P�k��jl���w�V|�����c�b��
D92W��-�{�E�����ko������C��Ɖ�����W�y�b�[S�MS�M�4/��_��pC"��y�v��)�������`����؄9��O�'�^(�9"�t�u0�w.!�K���=��h�7��.h�'J�;���$��>{��P��udR��ߎia���c��z���?$�X��C�,��o*)0��E�D2e�{9� ;�h�+��.4Ή��r��^DQV������E�����0;��r��W��Q-�&��<����k�R���m�q��������v��K(#�HVh��'�$^� a���7��:~������W1Rx�0�d&��-���	��ԤI���Q�F"��E�!���5�2��� oNYXOI���$Իt��,9��면�u)���i�%c@�t�I �gP��a'�I�Q�[�c���T����^E��_-@Es�2���a�y��&�+���Ȱ�Ot��0uz��
j0�I*�K����x�z����Ľ��Î��P���is���scw)�β��Z��J��h��a]�.�B�+�M�6U4]w�v\w�v�wߌ��|?x����z�]�w���� kb�X��/�^\��q������� a�����(���5�Zc�C��)r
�53$J�P\Z�e/6���3CE�G��Yl��Pr���A.���?3��-.���=�ˎ�H~��f���+���w'%��d���+]r��i,�f���3��Ԛb]�AD�&A���"����NY�va�O'#����?�e��=����Z�8��oT�q��})�A�3U.��SՓ�N��S?����p�y�q׾�����î;������fAsٙؗ���;7�� 	� Hp�f����%�d���c̈́aG�����Λ_a�<)�phfl),i�i������f���I�;�5	�	��������d��7�[��?	�:I�Uuo.'3O�-O��us�c��#����ib��%q�6�NB�1�Z&=p�Ϝ�U]�?�̧�c�+u�����c��Ng
[�d�k�%�x��D��yy�A �I/��F�=��`k*��$}a��=ᵚ�&[��$ТS��Y~�5����Ž�!��䧏&�Ʃ5�B>J/%!7��E�q�'�����)Q��a���<dw!m�����F�d���x����ev�"[����A��I��D�\M@t�4���?z�I��]w��k���hU��(M�'�9_���vS �	�A`�SĿ8>뿥�jR���r�݋�ˋ�q��s`7�]9����o<�z�u���;83�	+o#s�HPʍLQ��_�ex��D���ӕ����V��&�+�������9�63Q����z>�c�Ӵ̠�d�I轅���3���l]���,~!'i��]4�a��웰n��~����^�}ؕx�U�OJ��w?.*�7�vxFD!�L���=���I��3 ���4�ZF�@I���I|L��f|\4^�������E�5�5o�>���;p뾽����8��jl����P�3N�����w&�ݺ]W\���_�6��_���ջ�ZeT)�#���%�g�s��i��Xg�?8'R�d4�`\N�{0}$HnB��,�!�s���!��N�A}�ZG�:����5%t�q�:�@���M!��v�W^�m����4�*|nsb|%p����2�;��ʫ�")�\M
���c9`I&������1�A*k�1�����'B�\�����iƁ�ؠ���̄����b�|��N���l�U����f��}p6�8)���g�,��7	�o�9N���3K%hY��O'(�|�3�ZO�kRj�z`����ϙS���v�2>� ~��#�᚝�P+���x4^��s�ʁ�Ы��5h��n6C�6L*��mG�g^�ٺͱ)?�B�7&�"L��r��n�R�B���sy�>��d�yy(���<�g�����7`%Pk#�R�ӫ�R�n:Z�y�VZ�i��3����v�qM1f�����l�����B<��χv'3m�2�mDu��ꂵ��6G��c��Tl�������r�[�|�@D8�Ťi��{��Ҏ)�ۨ��v�BE��%Z��ap���F!2@��8aeq��>� o|�[�귿���zw9�}{��i� jR�S�N�Q8v{��ku���A{a�EA��>fkH������v�1J���C��j\������˯�
���1|���ĉx��y��E+t�A��Q]/,\��4E�ɺ;iL���n��G���i�0��'��!��7���4[W�>s��z8ڷȪ]ZӬ�O�6�~�ȝ��	�Қ.��^?��
���y��>����x�4Cc�O���z1����KE����#t'���*ݡ����9?}�N�-���=�1)�e�R<�_�Y�7�Bs��N��Kҭ��Ҭ���6����P"�%".3�q�$���&:%���o�.jFIS=TΡҮ���P�J`��{���������������-�q�޽�z�%����(�(�mQ�*T���~E�_���դ�5W]��/ނ�W&Ě�ZeNH�̡PS:�����|��Fo���X'	�+$��qpZF}R!*f.q>�e��r2w��N��|w!���Ly$9%�nGy��{��i�rxJ2�pm�F�Nd��B�����ǚطVМm���S��3��,3e��ڋ�k;�@Αk���:O��i"����t��;�t�]�k��ʄ	Mt"∤D|c?�U܌O�+,w���-'��s���S���]W�[n������yC����d�VA��A���M[����u����k=�Uѱ^Oܵ��M���#���!�wn���?�o=�$�}�Y�����P�fslb*��p��*a#3Y=��CF��E!d5���WS����r��;~gQ`�4� ��G��w�u�c�e�h�t��*V�B�?.��h�Q^7�Ie��Jj�\Ldg�f�f����c�N�Z�{Dc��&��y�ZR�|NI�bQV����=�I�^� �V�3��t�H8�"
�D��8�^���ό~�k�#��UP���n�k����N�{0����.�Rj��X�q��m���o�o>�]�32<�0�����V�ʍ=7�F����������<|��t�XF��(�09^�E&��lʛ)H��.Ю(� ����ۃ�:�#�4�*���o�;e}h�i]���Ы�}�(_w�������3��,3G�s���bų��kW�s=_׺��u<'�݁A��/u��	�"�m}B�0y�5	"�*��
ψ�IWn��&��hu��$F"y���΍BVmh/'�wN˜cɕ��Y 0P~��ؾ�1W� �SD(a�nz.1�U�C�`�4AՍ'm}V��)vF�*��P�_�z5.h�͌�ʕ	6�J���[p���y�zݽ�_�\+��Hi�P&T�%W6�p驨D��]�
֯�¡�.����x�ݳ���ݔ�6��(h���8��P�3����3��L�)9>#+��w) L`��rK�o����lj�� �O	˸0Ι�4���,��*[�d0�0��2u�� �y(:6��8}X�!���{c�s^Fkis4��}^�4�et8/����K��u�)	D��.M�D1�A�l��)�Sh�[�&^�Aa#a��P��
���մ���g��7��%?z 7�
�9�O�pvm�˅�7wQi=���Ѩ�6�@w6;�<�"<gM�6�k�w�(��F5�
ᦺ��W\��W߅?���x��������	Ϟ|XY^�Ф�iX(�g���d1p�]��><2]�BF�D6�*7��s�,�ʝ4�{53��G�I�s�$����<)u�M+S�Z�PR�ת(=���3u�o�tk�Z�3�+��I���S�	�r2�<�)}��}�jN��!.�Y��s����ƈ�q�����Y�4r�	P�{i��W� *�'��v���Ox�G�ʵP�Z����eN���?��
����F|��k�;�߄k�ځ��6b0Qދݞ�v|φ��T4�fB���F�p��x��)��Û"�0)y�Q
�	y���9��ŘǬ
�w�ߤ	:YP`����Ө �^IZi�PE�D�HX%�9-�R��)��q�D�sff� D�H����G�,Y�hԭί�P��t�`oE��ڥ���5$���I���:�Ӻ�M�v#�k�0��1Rʈ��#��2��В�h���U��I,0��\�y:�����XZ\`P�Z�#5DYӵ7�ͳ/��~	W}ㇸ�����ჸ��kp��M�)����	4Ԫ?���^6�����<�2[�Q5WbU�C��vT?�da�/ڇ���o����<�o>z��:N�fQ������I{x�]��6�l$B�ٚ��.U�}�뢒6 y��t�obه����j�*���TeĀ�b���C&�uHr3��� 3 ���s!��<z���=Ƥ��	�$�Y_���:]��}�e�gW�@��Z�
u�h�6W��ˌ*��7X��,� �v/�P�i�?�=���/�t'D�s�6�*�;؃R��zE�Q�2�f]`�e�qہ����w��mضi��7Ba���c{j��)����͚w�u�������܍�L�M�7���ƆH�kPhn�k��	_���oV�d�SG�	~,�8�f�x'�-�ub���\�f�阬-k�u�?o��I�os�uN�r���}U�X��	��`P⌯�k��9%?)���qm�y�TL�i3��l�dk�%�4X��r�C f�3U��*(��ӛ��fR�E�#��	5�E*�1CK�d��L+*��/����P�߹~:������&e���KK�}�|��!ٳ۷n��d�(��sRy~�{�7(��O%��O����".�~�／%�i�S$���(�q����u.G����� �#��Iu��Qx �5��~*��s-R�{��؄k����Ed�n�Ԕ�}�_w�	�*"�l|��猅��hΰ=�)a��oe[��r�5v�i�+�#hl�w�h�wDOϠ솬1�h~F?��&�25X^�x���k�������^�U��>�o~�֣�q�Nlۼ�.o�`�4�Ӿme���+S�`�B�'����M@�GK�**9u�Q�ԥKp������7�7���_x�}����x��9�7FօA[s=��3�9LG��wa��8{�
����x���ǝ֑�J��]���W�[�b�H��Īܳ�U��^ef�it~�#Y{�z������.�qeU�%2�I'��0if�|�m���Q�,��a����u�j;��^#�x�z9»|L��*�m���0�gQ(�����u(��U*�EP�>��ok�ưM��7)7�͸�zi����{�)����ĞK.�]���<�0��=b�����"���w���Iy�:�8x'��ՙ�
~u�=�m�K�T�Ǖ��T�IpM��ͳ��C��h�C'����0�D42H�H�!����:�/Y����:�s�l.�ɫ�����ۿǌI���� �a��O���*���H�����RqV:�_T&koTXˡ.�9$���I'��N!���c̃�C���iOZ�${R�Q
6���C���u�9ȳu3>�Lp��9<������o������K/�6 �p��Vhҳ����6f�d  ��IDATU:%lN'�V�t#�l~�E���3�]�D��P��˰���{�݁�_}?���������S�dy�AM�K��C�ѵ&��>��~7.D%Dt�*��1�./>΁~V8l�L��9��C��Z���̙r�M	�3M�Y������?��X;p��SZ�6�:m��g���	r�E��Z�@����ȸa%[R�|v5�Q'���C����L��9=��҃��xu"�v�Cw>UR&�r0���^�3�d��	�<;p��`*y��A[ꏽ[��S�w�#G���˱uÂ�v�k���>�
�'�v�3s�V62�K�a��e��Raѿ�b�x�]�5��@O�I��[�!w�wj�U`�x�U��A|_�ܢl*��|�A�	R�ϭ�M��~ �6�X�5����p���|�������u�8�6�x����3��ü��l�#}fj�������h�d�T�k�@뵱�B��;�~��/�iR:/ >56�u	%Ap�I��v$i���f�x��&bZ����R�1x�J@*_~��� k��Kwt��������V��5p�g���k�VP�ܷ���q�k�e�F�I]vR��ԅ��e�HwO4m:Y�S	$]�1�j �8�`4��]A9Z�B�/K�UИ�Ȭ�0c	 ���]�yI�.j($��
�;�7�-���p��l�5O�商��D� eO��{� !WG������M��TF��7��>��pS���t^���F��)l4`^�d��`�[.D�#�l:$
�7IZmR �}�~����g7��3�ֆ�-lwC�L�am�S^t�9Q��{s߃�zi�?z�}�]�q�UشhL���V��5��$�|�����
�����i�59zc����h��������uqWo������[�����ٱg�����>�
�Q--aiaC]Z#��72���1qW�s����7hy��$�!�X%FƖ�?�J6���*j��[u<�8sa���u�jM}e��i�+��\���JiT�Y���ׇ��{�	MU�,��/rc���'��b>e7f��7gq�ȭ�i�{MԽ���*}�:���H�Idc^�Bx�����W���F��jd���#sB�z�	s���붗��ti���5��,��������S�ߏ����p���K����o9�};.��`�'C�-���5���'P�'_<u���^��,3�VyG�舞���H�#i�;��O�F�sƲD��֮�aSYӟ�nJ�Y�x����v>�����ǥm+���3��^3�5�9&�	L�c3)���e27��[$�~!'q�&(3�:��{$�L1�ҌΣH x�u�h7�w|ٜUS�p��>6�A�U�Ӈ���#N���:"���8��壆�P����sy��z���x�[?Ŀ��đ���o�S��'n��[6�H��	�:���J��4z�vTr�lB�H��?����	9N(���ၳ�\�g7�ރ����8�Y<�������>�g�>���0Z^�B]����|������H{��9����t<Ǳ5?~�$9J+eGq|s�J�C�M��i:ϼT&) a��1��y�fH���Q&�hŁ���N��{�:�MmoN������A�G���&4
O)�fm{o�!�m�^�텤6W�B��U6�5rpG :�8B�a)Ϫ��@��p��HK��-I�1��!�r\�ϳ+��
Wlތ/�p��y5��a�D��v8��+���Hf�t�/'�|���M��zq��b`�2RTl����6r{0�z�O�N������"M��A�z��[�e�B�qsCrW^Y��W��R�|+��+���K��~k���3{�́�����jE^M�C7��m��7h�G��,��{����~�e���	��	DeF�`]�4ﱮr���Y�a���]*�UNsU�]� U/w��a��ӆ�Y���n�߈!�v8��A�	8��*�l�!&]��ڌ�PC.+�csb����p�H�ֽ{p��qǁkq��mXR��O}v�QBP�m��Q��0RW��~3�u��+�q��3x�ͷ1�S��6��B�E�#��c)�6;�B��c+�.��!N��u�|��+7MbR��v�Y����e`㿧��Ga�U�n�l�ԧ&Zv���x�S����%�JƷm�?N��\R�t&J��D*���u#����2<�7!�1k�q�!���,�$��@����8�*b��H���H���*��DOjū���
��r-�-\��Ɵ=�8���ppǥ�����٣����+�`���ʏ(��r�U!4v\o%�w(�hC���&S�*]/*G���ooٓf�umƾ;o���~�y����/�G�Ʊ�o���2&��5�*�1��վ�A=f����89�&��"'��/�3 �eE���Y�8���mVh�fL:��*Gܟ������c�_��~���>eg���܆?ۿ���6�n�D;$Sd�L��Gy��A���"����>ZKg���u�_������*��u��V�v�/�t!-��ه�<1i6���%3�:�w��*���n���dI�Eύ�S�/�mNl+k<%��89��X\��~����<��}�G����Wn>��:��;��%�]x��+�����pHnt.�`����o?�,VJ��%��`�F�(u� <�����+Ncd1����sE�,o��u.&�*���,�u55B=�^����_��6�h�j�B"L2�(�' *�MA�Mf�u�X{��M+AR�cM�{i������{�l1k��O���� g�#�q��]:\�l�>k?�n�4WN��9��,Շb��']#���u�7zN`���t偑�(�'���R(��怃�E�16�xQ�V����-6-���&���Y���o�Ͼ�Cܾw�p�F|��}�f���h��4�.x�zƨ�������*�3L�٠s�O�;v���p�s6�%��
ܵ�J|b����/}?�R��<�>�"ޜ�1^�`���f �#�_�aE�|h1*��v(Q9��GWOhx�tEݘF���4�G���8H�?��5��6�ߖo��k%�~�R*�:�����} ���v�)����̡-yAvo(��rz�4�#�/^'yn���`��Lk��C��}l�Ɉ4�pB<ۄI��wF�H�X��lU�78�\+
��U����V�ǉ�AΗX8w{6-�Gk��!�f'.ݰ��S���ՙ1
P;��M{0�����z/�J�pUn敷N��;�a��la(rz�N�1Rn쟛>ƣ�L:�v �)�Z�/3+)�fU�Mږ��(s�Q4��_���0m����u�C;��Qktȏ>������^i������D927OFQ�TT����3�u��\�J"�`A�N�����$R���t�1w"#LYwl�����5�U��x�S�k���>�����Z�t�ۜ=t��r�iH��Y8;T�@�u���Q��������:��4Di�Q���)���P�|�Xm�N�c���u�N�Mlh��F۸hy7^�w_����z�ٱ�5ß����B����^I�p"���*�������rʏ���_�����u�8P�K��sY�Xv3N�a�跬/�;v��&�%eViY)�J#����u9m`L���%a! �}����FL��r!7��6�R�-�E�F&@k�Z�W*��̌�=��W�F#�V�1�b2ur�]������Vlb1
��m�Ab=�~_ct����s�^-���L%!Ƒ�4J!$z�A��i�� �\����� �(��f��J�D�u��@��S~K9��"�2
�o�:�%�>p�� ��|P���x�{��� >y�����}8�k��~	5NN�[���R�x%Jn���#�+{��3h�hc�2�i6��ְݱs7nٹ���⾧�Ƿ�x�%N���ՙǋC�7��U�_�s�ve�6<���ʡ�֚\#�qU��^�U�i�+������FP���JY�s�W�(��%��6"r��Q0�2�>�����A�2iD�����C���\�+�!��:���"-�'�ͳ~��|�[����*����x7�X�X�7���踴m}C�Rs!�c�}�"��<�t���9-Ƕ�LA|�n��H{*-q��6���'O���+),i}A��I����E�߹�fj��Tv�˥ȷ9ϋ$�;������)�P�8����AEg��p��D�
��e�U�?ʪ���ܪr��;���g-�kqT�H��"^���������f���7��á�;��up~ŝ��TD�*�����ݟ?��>�(��6�ȁ��*:x��Q�x�3�D(9G�x�E_'w� }Sy������N����_1�Q��<j�m�^��<:D��'Χ�n�V�H�E��{RV�."�žY���:�y���}�\��j����ܜ�K�HZ�e�Ol*�s�e�!�b�ټF�R�g�(�Dnm��f������b�8!V-��U,��m�C�6���hۋ�͓�N6 ���z���9��')'33���$	���#������M�9��u�֏mh+�E�ᰦ���R�:o����g^�}Ͽ�]��=| G�ً=W^�K�n����ڥ�>@�����@�� ΦM=�:��X�9?ؕ�Y��6n�Λoo>��~�&��Գ�ޱ��o�s�0P.굠�`�����ZF4Wy�S�N�e=���A�`��GK�]���ݜDʗ����&Q���&��3$Qluk�V����֤�iy��M����>}\qk�Yi�ȡ�'�]u�!�`�"1GK��#h%���D��{r� �� ��\;�����<RbÎ��GT��O���=߇����hM�brQ���փ��|��@�X�T��tް�Y�(������6���Wlو[�݃{ހۮ�W^t	��C��w���+������������Sy9��]�)���/�tYa)��åj�;f���p�C�l�3�;9:MtߗRA?mo���5���Q9[~{9�0+��c�	�2n�꣼�c�i=HK���g�YU�|A�R��Z�M�{���+�v��$1�7�o[��[#�<}�h=g��Y� �0H7Sq5�O���Q��(HO�\��Ȉy�M#�G���y��ˉ����D�)�xx���r$�Q`|Q]���������Div�M�f�ƺ@FoM���N�w�;l����
x��1�e	=����y\��	���F|��[px��dN�����j�S�p�~�e�=�F�,�3Sf�!��yRTᙗ���\s�����Ļ�����?�l�S���TI�����Y^@bS��TOd0��M`���X�I�\JJ8������R_���6!En�党y����R��K��%��b�[/�*Z|�Uc���erF޶M�Y63�M��"���u�<��Țy��C�D+�����p�|hX@}�<l��),-%MرqG|��SsN�+բ^�i�)���h��I)!�x�Y��Q�{���_My�C�{~�����Gp��>{p/����+�v��n�WE�#�T�(��\v
�ח+�=�gןҞ0۾a	��!��'�����ӧ��7���2^zg��T�񢲡/+�2(�S�	a���m������~�Q�4�DI�ǖ�4�lM���Wź���Mf�i����A�ԛ��E?f����;bU���M'ǯ�_��Q!O�/Y�/�� � �"�jEj)�t���;ǿgI�#}�{�#G���n䚃?N�[�!4�ޤ�3G��?�\�ϙS�,�1�U4�{�W�C(�\�`$��px����I5ޒ���N����I58��*I�3Ft�em��#�:����D�r����&�k�t�\��?{ �����ឃ�p�M7`��Wa����`	�E�v�-|��G��C�VC{h�(H�ڡ��h�!���*>;}'��r�E�|y���Pt�P�.�:���%.k%f�z��(����i�v�4M�ONW�zb�4��Oo��yL�"庩P�y�8�I����W�Ա��Z-��,/Sr$��,�I��}F; :"@���=G�G�iUҶ"��{&�VG�_��'II�3_�*�To 
A�N�����+ep��K�w�=2Nsz`��4�H���_�I�o�����{X�����6᏾�)���|
���9�V���C�7pKA��{7�H7�s���ݞWe���):]���ف��+w�����w;��{����#�k��\l(+G��˚�
��:��u��^��lI��-H&�uC��]K,h�T���*��7�F�Es���[�wM���s��f;�1���D��׆�|���3�����Sc^W	�Z�PD�`rZ[��.t�*��9"�zB��A<�V4��h����PXY�,f#�6T��綹Wy��!�:	tքu�Ց�����i��w���d2��4�1�n��u�-������K122RY��]@]ѕ���)f����(�t(C'N����s65D�o굊G]v8ı��O<���e����dWun
\�6)�dl��,�A�j�{0�.�� �{WIv&��<�{H�؞���M9;}��H-P�ՓnS����5L|O�~���'�5�H-����M��÷%Dt�NI3L�Zn<����Z�X�a�9�I��{�����Ⓢ�&�f�v��X~�"9�����0��N�̛�v|��Z�/"S���� ��B�gi#�;W�ƒ3D����B	�0?�	E*<�+9��d�@Q�w��U�8{�\-4Lpp�E��'n����ciT�@&�Q��&cUz;�Cl��GUi9FVلu�0�d(:mZFo��������'�������1XX�
�;�Ob�@�ό�E
��~���@��HA�35#�&��.��҆PD+���l��r4�(� 9mP^�/=G�r����N"i^w���}�^��7�G_��T��B��`G�5��iF�;��e���<�+���xc�i�PU�7!������������j��h	#���N �H�}O����y�Bh�|xwCZ�ao`a+\wj]˨6�V�|���W��7���˶y�d�w2���E;�脯���>��*����QŦjSԼ��[�ώފ/�t+�8}
��
��������湺��F5���T�o:F�1쇢pTʝ@��[�WTUS6�
c�-d��&;W�\�>k�&}�I�
$CG|U�P��,���\���,���z�4j�$9N���F��+q�#�cE19�",�#�HYSH�C�|�1����ש"�޵Y�s��6.���i�KD�в�jR��&����S~��:05�Z�C���:
F���촖|�ˊ�S)WsY�2��]����"�3���j�]���Z�g��+�S�F���`�5O�����3��w�?���8|�v|��q�ݸ�-X,�x�������{�Μ�{���EХudw�/%VC�G=�H��G0�v1MyZ7��8{r���[M����-l�R����Գ��YxY�jVZ'�r����0�|[��F��� �S�:F�v��dL����]��4�T�W��{�M��̀J�6��F�A�<��!��r� 'l�����F�g�;�*3ݹ����X��dz��T$�!��6XAs�������8i���Ϋ!�]Y�O�{���&,oX��$����s�"ڥ��Xp\�h�Fa�*N%�a��ܷ��_��;v�_}�x��_���=�o?�4?q�b�Bݿ�FYTV�)e�:L20�5�!壷�1SL&C큏\�K�vD�ws3�i����[ZRЦ�3M
0cC��>)��a��I�t!�A@���%E}��ը"c/MT�SFYB�$f��>�BST�XS0������8���
#>��gx���Nʉ��`{0�pUE=�E�0N%ȁ�F�4qn��K�s|���Cܾ�
|��-���>�l�=eo�T������k�]�N���xh����;,>��a�v�xV*NJ�WM4ª��g_ğ��W�����89��m���u���c��p���YFA�FD�D�H5�1����ۃ	r��W�eVKo^�F�g���3��3�v!�.U��u�VX�N�Ma{;p({���+��CȜC�j*�=���ؖ�S'DT$$w��=���:�{
E(׶'�	����	H��$��!I_1�4~�i�J��2�$��{ ]�e 8�v{��� ��&LI�����.%3�F�/F�$�n� ��q�x�>Z�ty�r�����Ra�E��ȡø���q��+�}���arRؓbư���=jk��ǹ[ҟ���6e7"ᅇ `�1���y<y�5��7��{_~�j�pST�M?/�Q��q&2V�~��<)��p0W�`�{�����õ���CL]���YJ���.z�6��C��'3�U�JK���hR�T#ܖ⺘CQA��ra�c�?ׂ��U�y�N5R3K�y�{c#��$X#A��O�?�8��U�}*{��T�\ʓt�%��{FWN7���wD� 4R�ck���;q0@,��Z��E+�u~0'9��8�Պ�	WZ�x��_[F@
�D�����N�:\w/y��3����C�Iּ�fs�V�|�~���mؽ�b|��x����G��G�<�'�:�S��`�B�HnCM���
�N����9��n����M�ّ�6M.�IbH���yMC�P�[��)u�)ٓ�����eA��Ж�����'�+Vzz�h�
e�y�  !J�%٘�B�2��}htsc�Ys�c��F_>�Q%�8�h�H�'I}��E������kMg�D|(��	1�|mf�z�r�i�g�	OeJ[މ�/Qn��/4E�P^�yJ�]X�@W�"l �k�
����UU����!�P�f,��n��－�~�غ��͋�ش���＇�ϟ�V5*�PT�T�\�b��־j�{a��#95Q0#A4z����63@���!濳ˀd�A-�iN��8����׫���������~i�[8\�����i�n�����Bl� �s�Pd6x|��e0�|a�$�Ƀ^��:<Ka�9ZH{^;���)T��a�dF#�z�Z����02&RC}� ,�h;P�h�*c���i_�Oz��CEt�jȖ�d_(����6�8��J�K����Y��!��?'�Ղsb�=����w������p��9n0�G�&���-���b8'�Li�e�k�ti?5�[��y�8�k��sw������>����WϜ�����u��][i6�\Pw݌I��1e�eS�@�vJ���s�.�Ӭ`�e��^"fl��)�#!HR[�$�[�m�y�u~�ʰ�I�z�Z���Z�����ivIT�L/�[L,2��R#`L� ���s`�+ɧ�dz���t��D���c�jG�ͻj��Ѥ����_�7ݹw:��_��7.9�^zۗ�Vʪ�|;��`�N�P��=�<3�#��)����8螪��{~���ṳcT5��a�H>�Q�J���x�2V�u�oΣs{0��~5�p���y���N��L�#�wnr8 m#�Ć?�/����>�<��f���jI�8r�x%@Q��8 ��N�mz�\jx�
Th3Q��2V��[�-�V��=Q�lR񶝱���S���{�F���g7\J�}�1��V	v*]���^��#4�;;�޹��^3�\��)=K�57vٔ#�L�\M�,��/�k�|���oZG�!��!�@/G�/8��T^�g	Y� L_�q����� ��za�6�|���Yi6��RiN,O�
��X�L�si�>��쎛qx�lY^�'0q���ذJ+����p���s�K �L2��#jQ��������,ġ�G�~�^۳/�_��������Zh/�|=�"��	_M�k|���h�851��=�j��c��[J�8����Z�	"��{m����9"�d���~�3ϟ�7���R�a!�ɗ����=�6_�ְ�͗�ذ������� 
f16w�8�=�3ܩ [Fk���r�]9����d:ƹqL��L9?u����{X���3JR:dP�q��D{2h�Qrr�p��e��w�]Ckn2<�8���6�'����`���]haF��F^`6sJ�ScF60�>���X�h"X�\�_��7Mw�Ǳ%ΐ`e�/��te�q��8F��UA#�r'�4�lj��i8��˯��߽����x�W���wϜ~��mkeNA�ؠt�DZ����ܓm�T>J���Lόc��	�lI���6�!�H���Z��S���j�_MB�s< '���~�
O2��"�N�3��JhJ�yt���̲��u��q ����ʇ��z4����7��i:0�)i��mQQ�R�r�����a��(j�������˥����y�D�a̜�=r��1N�g�w-�:m�m���5L$��T�K:!�y#��/�;�=�'����(�U��a�ʺd�ś�/��T'y�l��9���eA���Ťe"��S��I�ߤː^O�Y���֤]36EΕ&�����Vت��w���8_�u�,���g�ߺZXƐ��b`�Щ9�������'���討	n>�t��������(sD	�l�c�Nj����v\"M��@m�����9��u7��ɏ��v��=Щ�(g�����;�Ta�X��D$��h<T����m��}wF7���F{ca������P�0�g�6���減I||ss���%�g�%x[���왽��E|!�T��y�Wȥ�'l͇i։x!�"�#8��LBV@�0,uj�{���ǵ,�q�~˘B��xbPx(�{{r�N601��D��a0W����
�fXu��[ᢿV����C��w"�B%!��TJ��~����ر�_>r�p��x�<|������/��WϽ�3������P�ڬܨz��0�|m�ϰ^��ɪMB�S���s�Lq�u��&s����N��JF��MZeR�@V�'���3�g"�ra[ҙ����o�ykP&�5)�F���:���P��	7ٓ �v��I���'�S�, r�6��G��t���r<�h�k�'��as�r��m�܍���w܂=���F��aXIY�/]��v\��N7�`�CtPP��-�x��X���h�u�:������=��=����O��7p~�T�Cw���66�v?&�4� sh���X�Mr"��
�'�t{�a&$�+x����N�䲄��{�p9�G*��T�t�;1ᱡ�ZSGHF��S�O(�l���c�Ƕ��4��r���#��=���i~�{��� ���
@F��c�[��4-E^S1La�JF�(Օ̚�����9��(�r3��|� (���5W}�k�A���׋Yi��p�\֜��5ɐ��a#,L0��;�(?c�gy��)ЩrB�( h�����p�S�8Ĳ����p:���T(��J��1����u��_�0n�.ٶ���6OQ�p���vJ�
׉z�����p��
��	�h_��F�8���5z�~��3�����؉7�I���=�62y-�'+8(x��9����e�MM�s؝HX�"����(q*R����I����J��P\y�Y�2�45Nsh�����F�gI����h���0�^"�d��ܚ;���gI�@�3X�xLjd�c���Q�Μ^+�}.W��K�+�ɍ@
J:���ǐD��k�	�"�R"�5"���t
߷���P��@pyp!��K�}���a]�v��dh�1f�t՞�2'�=!x�n�]�9`��T�lHw�+(ϯ�uUL���N>�gQ������;_(�L9qL�����yinٽ7����|	O��~��S��CO�Sj�8�qhY�1�.�~���X;ZoV�&�iΆ���Qp)DJ�*��l�� :��j}X�֓�)cy3՜����BY�V���"$��4r��,��z�&ϊT>p9ݢ���Y�cb^h���_.���-$MHY�4��s�!|%#��xY_��t�i�MwL��I$7)��*���-���O�/#*�4�}g��oN(z����[M�#�|<|�� �u�%�q��C�5�E!�ƖIf�a���Z�S{��I6چ��
W���N�w�9�Uao�Oi#*��3�v�Gz�ɱWǿ��}�'%��y�,��H��.��I�Ab�ȧ m\��G-И�Iv m[S�&2ۃ0	ќ����Hiz�s�V6��\�/FR�_��1K�Ă��m<���Б�18�pAy��T�m��5f��t�e���?�qn��CnXK�$DJ�=#�?ʡnq�'���&��S-��@�-a"T�7D{{t`��m���%�5�ky#q�>ZX�,n�)��(��`c���\���NQ��^5U�����b���!�_9��[j�f��x���g#��C��^�	s��Q���*LƐL�E�������_�m�8�_��F���i<�܋���<�K�yv���Œݑ�uy5��Mi�2�SӦt��~J��-)�j��"��䚓�{*��i�k�7�H�!�-.�i6��{oP~M�0V��(�DR�w�y1C��p&8�q�ӧ��3�b�3g�:�-�v�:ʫ����R|�K�!�T^�;��&U�W�J��bd*MeO�5��>���|5�W��l	����	�ܼ_��v��mp�5;�iy�;3)�V�s���b�j}By�pהs��r(�ݐ]S_8ok7t�𕧛E��s���+'^��籧����8�0�x��!�Ѡ�׍�A��Ydu\����D����Ӧl$��le�iET�UC�Ķʿq�2G�(����ƑXӉ-$wȨ��*�v]HG��2��쏕��฼�)uvL��}�2�m&�ذ'���̆	�[�6��0��fU[>�а��߾3�4J��������H[�N@.�$B�y7S�.��hX�H���ۀQ�g���-/R1�o����8�C��NXj�3���\��9��4��]�KΞ�U��ㆽ��p�u��K/��(�B��٨�Wڗs0h:�Mz&�@��k��xM�O�}c#���w����+o��_x��pO��6^}���y�Pa�|��D1�R?_59��trN�m/�"���8H��J2�)-g\�ᜎ��y��"ځ�}�.:�E�����ާ])'���BF)i���9���[�B�����-�L1	��65�-Uf����1Z{���(#P�(!�L^؏
	=�9��/-��&��S�/B�H5eVi���3Z�l���C���6=	�DcO	?㲆H�)T��:���Y_��C]��B9V��@k�ia3�O?<v��؁[�^�=[�bqah.۴��
���[��W�di8�H�E�2�6��	:��a��/*�y�nܶw'��=w���し^��_xϼy�&��y���;֕]8��G3^�o�F*T��*i��2�f��_�͓m_�N�����X]�n��������b�X�U��Yu�զ�GtZ�6j-|�
����]s#BNA�$ �;]nq�w����k��E=�o�X�mY���/HjТͦե J!�Yi*,� ��O�+7�}�z��e��"�Ll ���gR�Oe��8�w�|�tr,��Iu��d����-���s:$�.�]P@|������%���q��Gk;�+-jz��|;�k.[I���DM������ئC�Vj�KY㬼��./-E�v��9]���l�LӁ�or�h+��Z��3T�-S��^
��٦U��[��#��$A	��x�n.��x��g�SnX��S�E��������������G�h��Q�H�DFG=�5������T-1W�	֪��XJ��@}}��a�X�\�ֽ�G���mT��i��h�#ś_+�����85^�M��Ƒ�;p�ҲqH6@>P��Z>��6��F����Q����{�m���n��<���?��^�%x����Y�1/-b8(j^��`Y�Sׅuz�kc�𹙢�Q�~(H���G�i:ڤ�o��3�,B4%FZ�����?�D������Bq�I��|�Z�h�~2�M�Y;ja��ɜ�qt�\�F92��ζO'f��9IY:� "��y����aOD;gk�R��濳+XOp�֍���|��8�w7.ݲ#��S�Y�0(�`�3��xZ���~��287%���<����{�'�_ᢜ��w�����'𳧟Ń���c'���&����:�+=:����"�I�������[��X�ژa9(�M��,��Qf��4I42�ڙ>2����mK%��H��C�Uݯ�kmk�%;����E�fK�������_T!���y� ��Ͱ�=d�猉k��z�`4��>�Sʸ �SJ��JAh�y�C{��g��Q:��u\ ]-d�)��gLM"��Ĩ ���wA�`
m�t�<и�d^Aj��p�8���W��70k��ho$��&t
��wR�kL&�uܸ�V���
����^�];�c�4U(�6����xb�/	L*%�q��^e��FC�0�`Y���7ޛ><��|�'^z?x��Z9}��� ,�M����n�MGSv�o[�+S"����bk�e�v�x���R\�\��jC vB��>ޟ�ƺ�Qi�cȤg9ťO�F�ӥ%6G��8�S������ÙG:3�t
��R��$����Б����x׷t��H�?F��e���ˁW�^����4�(��)��zH��Qw�ƕjv$:����R_���fg��?���?���z��#����V$Gu��'��/��Ν�)��t+>}pn���v'vl܀��:\��������pB�Ɲ�y�́[�����,p��6\y˭��������{�<��_zO��6JsB�8�ؠN%&����+�4R���ν��F�rk����V�$�?SR�Y�7�{��V��������:on���n%�����8����UNaF�ˍ~zy5u�L�K��}�Ԣ;j�ju����ϖ�\��/'v �G���������@�Zi�o�,%{�﹪5��牱��0��h�灝0/�E���[��ְ��G�i�I��iNuZ/������x]H{`�*��6'�ͩn����P����_�?C��qt��Q�Ƌ`�Ǿه�P:�v���QF�0JL��C�T*Xࣃ�,�+��ҍE�9�S�8�<�+����� Yb�I����S���vWW����
���ef��c��"Ȓ��>�5��mZJ����[�T���ԫ����a&9*F�#�A�0��cr3#keHVe?S2�߷�_�����4��*�M@��p��IΕ�J>2��������8n���9��Q��4����%��=��}��7�'~��F��{���_�[\��W��������v�����ߦE,�ȓp�t*�p��6�V�6�]�����}Y�Փ���O��x��:�:7��F��UEv�.���蹂vx*���)>g���Ȕ�*y3G
H��|$Z�Y��ܧ%������K\׺�R�.�5�XG����Y!��� ��MZ� ��^�L�U�ޘ���b����&G��f�\l[{ص���h��+�Ǖ�2��-p��}���q��{q�֭�4�	�r&B��U�=��*=�+=�_�mN�t��`?�ǆV.
��b����k�ٺ�W�~?��w�cx�_��<�.-BGXX�]nxd��8����YBڅo�S�����^x�r�8W9BY��RD��߀&H�4�s-� ��;:��S��~��H#�����nF���r�����w�V�L�Q�O;k��C���d���5y1#�.�Ye�ɜ��0������Re�I>՚R$5ݩ�Q�x-�Ծt���h
rH�+����b�.$4=V*4j~�(�Br�8���WX*NP��f�7�F�ih��(�&+�g�a��u�m�|����M7Yb�V0�
�XG
wTم��zb۶�.]�����&�c�a���[���ԅ������3+x��q��O�;�?�O��r�T-,[0Ԧ��>S��
tГ6�lD6'�����D�[gh��1��C�8i�J,6tJϕK����/$ I��3�[�釡�u�TXS�d(�1�͞R&�Z"�uC�F�m�`���I5��<L�g�W�1C<��+�x�1fHǮ-��[��I^k���2!�A�D!�G��k��d������3�Q�jF@�Fu�Ȉ�I��K�\!��X{��p`9�u�.,�nn
��:,{��?Ŧ<��l�
Fū���Mx����pߩ����E?}Wn^�]7\�/�r�v^�K7-;b"i�+��چ��"\�(���V�2�G�#I�Q(p0�\u%c�[|��5����8������O�~�<|�$&F�ȍ��l�M,�B�G�'v��C'����8���)R&e����w��X�ʏ�����,tl�7Kɻ�R���^�����j�5��R�x�pжx0sxUܹ�ã��<-��5��|8oj�܈�s��!�;뙘����)/��! iC�WA�I��5E�h��/43�|�����*nxJ�L�`W�t�h�F|�5-ДDřu�x}F�;�5�yŹ�8�._��~�R�N��h�i�cv� ��l8��I��}�t��1�yɾ���ΉP*�a�#�_<�(��g-�ջ�@�,`ԭk1�B�C�TY�#4iP�B�|�]5�غ�$~�B��Z�&a��k�fg�QwD,��tM�ͰD]$��G�/�k� �$c�N��_�u��Д��ܵ�)JI|a
'�����"��Eׂ>�?5�N:\y�������H/c0(J�u��x0ęb���>�x�ث���/��oߋ�.���;w:�k.�K�T5N&_ ?���O�c\������R�P�gKmd��}���o�:��|��{�G��k��cP�e�Z��\�� ]��͉�:-F/���τ�߈����ԧ%1��I���l2��ء~�d����9��e��#Ol!G:��Юbj:��v��Lv���t.�����(։P���AC�ױ�"�:��=o�r[�\$m��n�؃���V�_��_i2Ξ��5G��}���܍ۯ߇�M�'��=���0S[i�ڈ�^>�H~�Й(v���vQ�w�֙���^/��`
U�|���S����W��'~�;�7�ش�jð�3��(���G`h�pYl��"�"�/T�H� Gy��S��?M|i �ͮD��=Í��e&���3�I���t�!a�J�ϭ#�@�B�8�U45�h�O~p7J�^ǬQ��
+I�eN8+&�4m�2�����a�p��-���E&�R:�A�@~�FE�ӯ�S���I�FjZO�S��䴱�6���&g�0 �����q6�a���9?��ꆁ��T�T��A�$� r��E���>��>1�C^��h�#��`JD �l|��߭fE��1t��>ӘԊ�d\3�I��F�n�_��v�uc�lnߎM��%�r��P�HQ:�h�Ϭ�aT;����Ai���Z�2%z�r&&�1S�ȝJ=7����o�g^Ń��S'^�Kg>�;f��J�`��z�K���?T��=q�ô���2���	���{e��L��ϥ��I��5�w��n��t���mr�U��g[�:�}}��#̷��$�}O�F�M��7(�9GϕeGB��f�h�r'x�ǶyW�&i�D?S1X�j��-{_�n+wC�"��r�0s��s�a>~����)�y�m>�pGr���a"�e��Ȁ��+���I!<�+��5��	��N���`�R6��C_Rۦ��a�����邮)��Zz�ǂ��ǒ��p�������N*G�]Z`��G��߇�a��-����s��=��=�,vmX�����g��];qqM���o�-�!&����!�H	KK���0�T�Im��%������|��-x������&x��-/@/PV+KUz�D�#d�]c���ȃt�;]��w ���d#ջ���� ��ݿ\�Φ���і;������|�a�,���Br�q�r�[I'�${]f@ۮr� ѵ@<��?�[]�ɯi)E�E4`T"���S�S�I�?[yN�c�븆S���w���ݧ޴o�lG���ۺ���k�R��������{ZG�r���O�|��Z����ؿ��� �%�hQi:Aѵ� 僴]��$��#^��'�k�����b&H(o�<�4�ٳ�"�Xe$�MAϋ�JS"#�´'"J�MԢ�U~a��]c�ސ�����K�L������}7��--���m�ܜx4 ��Q�ӐE�)�P�/l����=b�+�#�&���=�lܭ�8F����ԐI0Q	ncǠO����M�v(����cD�T�:�8P�5#�h�G���R`I�*N�_\ܑ�a����'�/�X:0���Ʊn³�m���䉓/t�,�y��9�*��n*�c�-^0:N
A�Qt]+��(9�6?���΂ZayT`8py�[��\���O�<�G�{��{�Ám[�#�����a畗�eFP�1ܪ`�J�1�C6֩ni�1��h	���񊉐8ā������œ��O~��t�����3P[7�cS�,�>'�z '7"�]�g��������!si��	Skx���6L���]����St�U������x�����f�������/<5�e�	���<��R��ͦ�}U-'}���q ��x*�sz�~P�4����	S�Ɛͫ`zE����]*�+�����Qf/�
�I�r2�*'�jy	��ډ/��] �o݂偑�VP���6#{m�ۿ��+�F��:h���*���W���6tѝN������ƣǎ㑗^��o����Vp�d.b��`+�B֞a��Z��F�J�B�=?����Ld�`��-wh��_}8�D#��Ҝi��ο��1H^�6�~��"���.�Q��)�����]�=��ʰ����~��?�D�a�n�4�*A�:�U�(�k�H�b鴞�"!�LT�&,V�F��DP|��r�j#/�6C��F�{M�>��Uyb�f0M4~�����A  ;s�7\���53��7*.�� 4h979���d����K't������q��2��+�5r��(�%Թ1���_~%�n?>�:ص�mخZ����2������	-�J1׿SA/Lc�+$�Fa�j�具O�O������pc�_�\�J��{�Z�`�&�6O����n|+/))��ݜL��a�Z�C�79��������Wr����h!���`mD�! AND�=�k�v�5�1�>���Q�"j8�֑ G��x�ާP)61q-'��} l�f�|Å��Qy-�Z9Kr��p\X���4>R"�N4�|G� �~t�׺xd�ׄ�U(��S�6�#�*���R��9˲,��S6[�5�ʒ�m��:j^��0`C���tz���W��:�/ά౟�����W\���܀���n��jz�5O��K��w�>��w�f������1�'�\/Yڄ��z�_-���c��o��x�L��k�WbX��#\�Z�tM�9I'.S�c|�hV�[��f�_"�/���i�������1ՠ����+)���F{]��.6Cl	k��[c|�m���kkk%/_�:�0�`+�/�\;^�Ż���/l8����*
�<�=r��}�+��g�ʬ�;+⟺���;5��]�9�N�R#k�u��}~��p���yb
K�:�_OC�H�<2���c.Er��;Eb�
�)]�� ��ul�����N�ޛ5�B�٪��R�m���2F�K�Kl'ʄ:����ͫ�Q��Ѫ��2�4GB� �mb&�D�L3~�by������M�ND9��CCFg�Ô�,Ǉƿ	[Q�ae˶J���j�Ǽ�^�����	s�E�����h�u� Yd3��g��G��e����T9Th �k�3�Р���ø��!�6��OE�&F�4�y}����lN�ͪ��y��IJNGXp͙������x�$~����M?�M{w�˷��ݻ�F�Ȝ�^�g��Ig�eB� M�����.{���g�s<����˶����o�+����[���}�--�,���U�0�VQ���o��r45�]�e��'l�˼�����zNn�������ks~^��	�BI|��|����_$Xɋ�F��dF��k�1�Nc�4Ѡ��d�G�(�eF�� '(=7l�k��(2���$&��+�T�g��j��_�sUr�ʫ��`Vp���x�^|��~�s�Z\}�%X��&5��&>����d"��òDy�~��'ssF Ǟ��7h�w�Z�^���q�s��O��<��i�S�rfR��Q��D���Ljn5�N�pN���[���yN�o�\(a|�I��G�'d�A��u/.ä����Tx�x�������ӄ70���m�����\W�t
���������˱��!��#MU�V!;`6��Ҝ.GE�l !��T(�(�L�ӑ*���7Q��D�~����K!���*>F����C�y��*bj��¯���ڗ�^|eE�|�ҁ�Bʄ�Ԁ����6hi.�F������a?=����Y����(� a�kY�h%g��P��#��w>�	ݿ[LXǲ����ia�xQ�BT��Q`�����~�rkBQ�S���C�0�:P.���t5ޜO��*��cO�M�Q,��М,R&f� �QZ�X>ܫ��^�d4���iLīT�w��7\V�a�Pɹ���	Z��##|�n�g̠� �;����w"I��%��\���g��(�(\o9���N��o��#��W��|�u�ie.�,�yn-Rf�|��K܏�,z���A��{�� �s��LЧj�ha�O�&�&z����<�1�q*A�8��e���`�jN
FX
l�(���x`Lt���W��d4��(6��Xa81a{{ô=�U(�nJM�W��6m��5������7���������?u+�\�K�8����Oʇ=�纬���P�z��l(��ꛊњlޢ���D�����]���{�����~��..Z=��ŷ��]��[8��Ȯ��"a�9���Y׼̚��Υ�n�4"q������k��9���t��5�8th�//��
�R��x*g�pyBԗ5N윽�*A A���K�~���������1�����\2��ܙ�4���سn~���V|ڕiTcM� ���;;�A���f���9�|���\=�#��	+T��G�����Үc �t��D�`���茎H���Fb/[�u-F�E%I�_"�W�4/����q��!=m��i���T�(*�!��AHh��殝�����,mv�Y�W=�I܌%
.��j�ym�u���#�
��6�-�B�qV	L�q#G�p�m��(�	�����s3��&kТс�G�b6�8������HE�%�"n�s�,6B�t��UC�%��d��'����k[W��0R�i�>O�М�#�Br��y��1��~9������7�^�򲱏�������j��}	����Ƌ���>q_��&\q�Ez�w��9�;��C�h�F�<��N�]�8����E�umc����������/qS������'�=ΩQ�~��Q������e�u�anR��E�6����.�0^�$Zv� g���ʯ9�a-�|\�3���̯ט�p��\��`��#�������6�3�HР|,2�J�Y5�#\(-us�X��<���:����EN�?K�1�C���k��߹1��c\�e���[���o�uW��������^�/�x��Ю���E׈{0n��`���ޛ(�����t�'s �p]M����z���+�l\�`a�baU���1z}*F�3{0���d�e�(�e48&g���Nq�y��F���/6`�ў#����$��}!��쁤�ے��d�%��`80�b��ɣ�q��ruRl�>�lB���Dv>.��d�Unt7z�ƻ/�DאDD�\�tI���ӱ�
�x�J�.��6Z��o��<�j7�s�ɓ2���WYw�T�t00��_=���G5�sA�$��|�q/m�/0�~s�����I	m���&ôu	=�p���p���������;nő]W`ۆ%��`a$�Ii�؊�VP�g���w^�����W���ҝ��V;,m~7H%W�ӹ��}�EҀs�lY�명�Iݟ�
ơa1�@W�Z ��R���������T�8�$��s7Z⺥�*���{��!�|�b��uN�D\�n3�7~���C�!��E5�3���(S�[9�iU���8&}��/
ea���I��Fݜ �0\�3̣}F�	�/a��p���|v�`�
��HkA�I�m��v�v��;}ï�Đ����P���4r���fE���MN]Қy�2S(w��y�R,RPͧ�^�B
g���~Z��7(��Q9�l7���9�),,nD�P�T��=�
�����-������m��=Wca�5^A5V6�����X�_�~�N��b�i�㟥�>:�W2)���'nϮ��;��������>��[�۱�W�a�6�gK��P��D�\���$:�x�K*�>1H�α���	�$��M+��K��\�Y7��q�H�4�M��ː(����W/b��!]�޾��XƟ],i33�]s��1�'�cؚ�{p�q:
�f&<$��Ϥ�!&����K"O�aÇ������V���O��N�O���Mۓ������Ia#�O�ݽ�yԬ@��_s��(�5��@q+����s��UL9BTEJ�!x�@&?%��Y��ڎ��T��J�O��"�M�K�<:7�T_���-o��/��q�/�X��L'��fN������<����X+��$:'�Vҿ 4�Y�4F]@v𳩇��[zm�|)�����XIh�����&�a�E 8�@�?�!B�`�J:�!A<�љ=��)�:O
��&"׮��#i6�����u,`�xJ�%��z3��<*>�ktNv�wByG3emm�K({�����.eq���� R���Z@�T������i�d�u&��U�ް4������B �MH-�h(i4�0B�#��#�����1a����̏�C1��+<�4�F����Abmh,����F��߫�7}3�̓y�޺U�����Uս���s�s�d�_�!��o��]����f|�[���=(�	`O"���r��R��:A����q���ǴV�@�4��y2�HM��kj�߼�.|ಋ�?�?�
�{zm�h�vX+�늈v�/�����<��RN�w=�ΩTئ� ���Ct��S�W�f�S�{%��#��K0���s�!�`�CN4g�䜡���o;����^��$�K�Qȣ8�(o_8�߰��6Ɇg�?y��&:��2dZ51�'��>���/į���q�����/��1J��Q�3����B�fST�8xV�)�lmv|B�rr��m)l]y=�&�oBr�G6{�wS-s,���:h���ܑͦ��5��ty�KIǽl#Ow�7��T@bl���[�����6)��ΝL9�מ��]�3��������c|R��-��f�	h�A�wnA��X�0a;O�����.�1�:ڜ㼘�a*�.-�(�v���
[��T���ò6��w�g�=:]��A����zW;�掫�Q�����w"or�u]rLBӮV���bL�v����(cfhy��+�}k�ܴ���Y���N���g�8�4��� (��Kxx�S��_�Ib;��z44t����8��7\|1���_ħo�	W_�k�.���mŋ���O��:oh��,=<k�.f*�4Z����9�B�I:j��.;1n�yG���
��������+�*�K�F5��va�Q�N� /Nj�U+�72�B ��H�d�~�c���J�8$XC'`A��#��;ז��*D�7�&$+�X8��B�2e�:�|�yo6hv�3@���B)�{��؊�.i׽kT�xL��u -��I<,�K���������읇�"�9S���b;�r�7�
��Z���8AXs��_�Ƥ�>�R:��s��"rΩ�_����<���T���4�F��F�yhͱI�rE�g��H��O��O�I_sơ��i�ܕ�{��7�I4;����2��Z�D�,~�Փ�������0n�d?�� >q�8�|��X�c�����&��/��ф���Vi�F>	� ��� ���N��?�|��ev�?}�!L�)��Ry�Bz�G�6`2�(eNk�wR^LI9ٖ�uC�Ui#��,�1jp�s)o�x�a�k!mhX�o����v�r�����fw�5���
�S����N�-Rt$�o�'��N��/�V�΢F|^��
��m�[�r���S<�Փ:�Z��O��tҚ�-��ZłT���O	�"�-��9�Sn�|���\<�8A�=��tVfe�	���
qZѿ�wr����R��*��,mUF�1n��B�He;@ќ��}�U~n�^+�6�x�[� ������zI��-ؽ�S��Od�p,�L�x~~	�#;����i��z��r��u*�Qvx�1;l�S�G�x�n�Xċ�-���oeu{%x���#�{�Q�I��Z|w48���y,-�8@�<���9]�K���������1橭��vs�\k%y�=ԛ�����!�.iK��A�z�]���6��訌Mr�v�<����㿥L'����cp��)�7HI��[��]��{��U)��nc��9���U�6�qӹj
=2l+8>����G��O߃���>y����mW]���v;z��&͊ŉE0LE،����9�H@%i��͕��u�U��_���O�����Tui�p��YH=1�5�Z��}�0�����wG.)�6���w��#Ǔr��`��M���C,[V�wA�0������{2b,
,6�C�D{�*!�8^'�B�I�m7�5��]���ε]�p'��S��f�h�����铧�6&�7㎫�����惸��s12�3vފ��[K�ڜ:��X�	<D��mb��J�la�@hmr���L��E2�;y{�T�]��0.������;I��olvf.�aNfb��:��9_�Gʨ���jq�YĦz�I1�4��{�ñR�q(3������n�R��ɔ4l��)�Npx8Qل�$SI޶�:��:�x9!�m_`���X~6u��좔e"�r0$cI��Q�x&��fzJf�0;���MAx��{.����������&�C���]Tf̲��h��Y���jA�@���V��gR��?ʣ�T�3x����B�]�R�?���ʜ�1i�L&�4���Q��\-~��7݀��לS��ìu᣹����42h�Q��qc�`��]�:�a)wN��]�c�8q��Dh���P�+��C�M�=�~��.0�[xQ�;�P�R̱L<=��h�I:�CPAs��D�mz���?>m�j�T�^I[$܈f�W	a��<�B��h~38"����$M ��ɢ�g�D�_I�G�M�J�6r�ϕMN鎌g��E�̈́��4;�ȱ���O�[Rd��l�j}�t�N
����̫4Eo��$�R�r���#���r�|�刎肋+��oU�J6N{V����e�H��:L#�H`���,"�����+x���^�x�y\��U|���q�M���c��]�d&3}׌bYW�������	=x^D@�*���-&IM�)�s�r��o�|�<�����8�iڢ�p~q�U����|�ӢXt�<>����g7O��|�!�:H�Xw�>�ٵ��^0�_/�G�He:��))}�}�4�_:��N�_Ð�,>��w�:���0�)c���XfK*�N|=T�3�������3Kn��]~���\�e� �J�{B���D�t�ʼˣ��A�������+�����,�;��N�9��nc.S�:���Y�>6Y��z�PV�χ-@G�Q������iD� ��MW�TTI��ktD_N�e$A:ԅ<D%E�Tԡ �������9$�ʯ�O�Ә�1�JY'�G,�u��dC['���_ؒj1wd:a�(��
��;�I-G�+���.�CѼ�2���7��(�1[S�I�.z��Ds��V^�ȡ��Bg�,!
��kBM��s� Y�a�g�t�cܑ�9]����g�te�U��Dm�G!��g���ZY���y^7	�]#L�1~|�£?>����qǁKp����7_�+�]����&n���
;L��UU~���Y&u���)�@U�+����Ĩ����G����~����'X7���G�����Ƨ��F��D2S�ɚЂ�Q�Ǡ�1w�<F%�b&���|z^g��b��Y��@���~��eW� z�L^r��P��R�2�mYC`+�
̷x�f���q���K�o�HN�+_N�����`�U)����.�ք�j��ͯ�)�M%Ӎ	���t����;���W^��k#g{�&�`[y����	������R~�����
:sV���4���4*�
�ע�������K7�F���ܵ`�Ȯ1�ψ�K)4;P��A}�=^d鷃��	��n:�A�@"����
���k0�J�F~'s��}��Àvn�G���϶�ϱ^�rzqO�;E�Oi�ߌΖ0�4�mD\�b��8t���� �t���;����wK�
�h�`f"�eOl�JZ;�`D�gw�͕��l���3��^ �CG�	� �L=�����΃]�O�`�T��t��?33��������9<�Uue���}Ԥ��O0j��ţ|��kq�Gn�Go����e��[��.���;U`�Ӱ����-���|�8wM�3���7&�K2��:)�1���_e�x��)���q|��}ػ{l�Z����s)�Rk��H�Q�Ž��)r�|�H���NG�j����3��!���0P��i�G��e�*��4�4�*א�IE�7E��w��D{�<�Ӽ��<�7o%g ��������Nws�W�2^r=�1vz�1�
gFy�M�.kiU�JGO�Qp�О�Ўw���r0_+}*����j0HV1�t�x#��C&˞�C��PN�Ԑ�*
�+�RY;�w�gQ2pw;�J�U�2�&�)�[M��3 �,o�ԍl3W)5��Z݅�֧�ѽ?���0�_YÕ{w��}��5������"�4�NkQWSO�!�tDFGV4\'��YF�S�(r兗�W�l��Q�G#w+5ŗ����ᏄV�ǘ���Z�1�k�h?C ��S���5�(�4��z܎Gs���9�8O�����EF �W�H�qF�T���wq,50����# �_��L5G�v9�Z<M���Z��'�"Gn��<s%Շ���t�������RB3�>����}��>�f�3��![o̓�cM�_�DF��Q+;�	KE��OR�#���>���a`6��I��^ͳ!7�￼㝟�6�{b�?�8(� y���&�o<h���0`,��}i��:�I�-��M���ݎ�TIw��lH�.WD�8˚��������MJ��}$���h�{}�p�F�$���V�Y�D��Cy�<r��q��'�IƼ�ԁX�W���[�Ikůu�`�h�U��s�0:�y_zLJ�U}�
�o��1*�A����И�����n��3��+O����\�s�6��U�q����O;�#�OZ:e�ӳw*�+���:ו]�s'1��7�r���a�X��F�1� �����e��Lq��C��K�avD�c��̄<=�&/
R�y�̚��b���FW�r�{7�OlG�R��]R=��lR� r�g��[F�4�\�T��]�9�ʦ��;t�jw�,v�sX��k1��ڮ��+tui⦧6�6�q�9���7݈_�譸�+p��qv�]�b�`�ɜ�]W�e�+���������\{ٝ������)�8��F��cbqr2��o���GO�c�\E_Tn�/�U���nP`d��P���;)��z�iϯ�8��{�EZ�T��\��.�Mg��9z�4��/�� �k04�@,�����.89�9�ِúg��ьC�0��!��dX�6�=����U �C��ᡵK9	��%��"Gr���J5�������z,
��3F��)Qނ��r"BGoB=��&��ʂb 윔�K�= � <�PA�lX��:x}N���F�Z�$�7J�g����a�u�u���s0���P���ף`.O��ך�s�ב@�c�
R�
��U����/{f��
uS���|?z�9��w·�Z����~�z�5(M��X���WBxZwǓ�;d<2��j{���Ĩ '�;��/Ի=�Z|���I�0��㺤!@'i�rR�ϣy�d/I>(�:���e�@�������΃�Y�L-�%[�c�.ݮ�ӄ�jԷ�o������A�iYɩ���id�)��E�#���{2O��I�~, s�]a����b+T�JX5�6iw��Bc�kDa���c��,�>}+Hf�ᑿs%��^�#�^7�7�r���X�_ǋ����'�����n�ꢋ�4K �F��)����_���
�R�Ȟq�o�Q�	ŗ��������-��}+�^��EGa�},���4H1�1neB��AP�IS�,�-!�-����?}�Gp>]F��-,C�JC��˧�m-g��]! �(Pg>3*ogH�ˢsyu}�qB}�Nm��B^�K�w,�ۭ�+���!����:����S5D��5@�ɀ��)Ʃn�}uҊ0�̉O���1�k:J���@���G�����q�[~�1�ڔȃi}�@t� �: �3��0f�B���]<����2fY��"^����l;	?{���͂�#�^�Ea'I�"p�J>����͈�<������e���)��c>��8&��HG�J�HgQ���ı���E8�4���}��� �@�|ǉz��F5��j�~��y������>����+OŶ+1����D���%Nq��Hc\��1��ǵ�����Wx��EA�ې�r�ѳny�:�g
��
��	1����:�=�`�,
��1��O�4��υ��B9u>U�x^W�ڍ��Osi����\��*@o��B�v:��i��Չ����z�_��V�r��8o��LLcG�8�2���O`lI�n�w!_�SɌ��s�+NW�)r�r(�(Gv�\㵡���k������|�\�?���8�w7��]Q��s�o�����e�����PvS��fk&Y����b�}����ZT�2�E�[*	�I�V��=�F杜�A0��f���3���3X�i�N�.-B-6Tg00����v6!8>�?�^�"8��f)��η@p**���� �Z�-���n�L�9'��Se?��.h`��ȭqa�`���ıy
�u$���d����7V� ��:��̴k�;�N�0}�u��iv��8%�ۏO~�F|��7���.Ď�U8���}������t���W1fw��ߒR���us�\m��7��ۓ<*��S�i��W^�=�?�{y��r�N��s�\���d��=����X)���Ôi Bi�Xä��w�t�LN�s�ʌ�(>,D򋸆m0� ��:���LnD�����I[iS�b*8M{�U�+�	]<�|�9���t�B����:�d�PlS��җ�2ٱ��I|����o����߻���^D�D2�C��ē�ҽj�Z�b�)$�����p<�F�d0��M-!���>�VyQj%wع y��Þ�N�a4+�<дˌ�l���]Y\W+v�p��w$�N�hs\��t��n��D]�ؽK���|��+��w]{.9o����R_k>�@.*Z9c���B��ꃲW����[x����w��q��R���,��������o�`բ7p�@{GwF�$��-rH����u �{���aO����jG�y��KTY��9����dx`��v��<b��a��;ev ���˗��$�Y��[f�A__�
9*ɥ��l���"T2#�nwy)7�ɧ黎a��d��P�X�kU9��T����4��Z�iJ��e�(#)����j�2D�a�I:�=��������qp�؀)ː��Ų*6�Fo@
eR3��4��v�r�ǈ�J]wq�O��|~���A�霒GA��RE�S�ۧ�3���݇�E9�g���~3��C��	��>ך�����D����'�X����	�M���� ��,�g�
��g;��A̴�������٧̩Nh�A1�8{D�Q�t��Y��<%C�kZ��#��w���"{�=a����ٻո��;-�����k������?��p�^�nt���/���/�=W���D�uྗ�ս;|��9�ѹ����maZc:�DyB=�?�AOH��>��mLC�~�n�����{��%���/t���H���C>a?;��s?:��+e-q��yd�a\n�(�4X����]L��o`�x/��|�-���kp��0�NV�4~��0�Y���H�:v�#�jsz���J�����k�b�vT�S�u�v�U<~������{�����c8V�����Q���4�S�A�b�:�֡��&Ş���M�Mж1�]."�Q�&�����2�k��C��T�*�|�F��#���)6�y<�k�Ǫ[�:��~V���.4�P_�<v<3�ѻ.D�����Ya�+T�c|����b��W�6��?�f�ºhiJ�f-?�\Y�T�S�1H��`���$�3�wy����j��(	:�c�4�r����&���1M\95*�g� �
u*B,���S�7w���*�	vV���݀/�s����cǸ��'ا�;^
M�Cs��4�O��*�)��x~a�k��1�M̑��o��O?� ���'�ĳ�k�*V�Fc�睃]ʵq��Ǝ&~� ���_��i��)��
+�xH;-\ �%��8�t+�D��8����<bM�cW�EԤ.I>�����C�;Zw2�C�v����)�٭�5�s�Ӯ�!����!��~l�QZЏ�����\�t`�f�E��{@OJ�}a�|������+�>G�y�W+�V�ҧ*���D���&ߧ���� ���;�!� 9�f�F�Zf�R�O�|�s0��6�@*�������,	r-�6�i�ʓ�(���"�b0N�r���/JwW9j���x[�;!�QS�x�
~�����w݆k/��y;i��N�ú~(r�����x�"�Q5�K%��� ���t���Cx��c�Y�&�vDDXD�3~��0F������Ek$�U	#�<A:�u��e*���R�3D��	���;�ؿ��=�&��XR�:�r�Tʛ�5}r�SH�s���s��g�/�;t�ۓ�w���m��_�G�d��c�y#4��:%�ڔ�����	�~	<#�S%N'��q�3��o�O�;��U&2��/|�;�2g8�#8xG<QI�&?���/[@4���*z�8��x�#5IG�\�'��Mu�A����S���8M~���#ʗcc$Xċef���9�E�u����ɛ�}d]g�	r%!����%/����8����W:�w�������dv�˚5��C*ӻޥ��4����#�#�=���a��%u�eڇ�q�qFd'�2���D�/��(�7�GV��ko�4�E�cd±:�R��QE�o�/l���Z�:�3b�� ��5ptM���iU�E\f���g0T	sI���fW�Ğ\8�X�`��P�..N����o�����o���?U�X?M��"�Oi/x{�r;�˂�{�K�tS�i��NO�g��>�v�]&�u��;)�3���yt��\�
B��HG3�{.���[nR�!�o���Jp1|L�s�Q��W����ш)�E�g�O���έ�N�2�V�o�Z�����/�fJ_t�"1h<u�S�<b�`
QOr}h��C�IN
��?�#�=Ѯ�Q5��0�v�O���K���ӟ��K�o�����{-�F��`�����uZ�K���'P�*<� ���٥
+9��˯㾧�o����K�Y]bZ��j�}�a�ɷ�g{FƖV5�X'=됡�L̇]�Fʭ�����M�`+m����rc+�P�:��:I�s�"]�k�ە�qt�Wѥ�i�Zf<��^��%Oۡژt�y�2�ԯ����F�F��E|����I�	H-�d=
_h�},p�B<{�����
JGR�3=�oP:�#��e��m���(7ӏ]uT����5���o�R�aI0!9�*��s~X��`��*�f>T5��'��+����_�b��8lL\>�Ҵ�� �0s<�=�3�K���q\������]q��ԩx�ȋ���O�����׏�&���
�ݥ��Ss�q�0�F�"X�3�j�U��g����W�Q<��qb��A�^
�d?�sFJ]�PRE7Ԑ���:^iL�&"~�D�ʏ-�gJg�6C���8Me���19�y����m/����%���u_y���uZG�
�"�彨��|<��b����61&�њ��w��Ɨg� �����t�0d��.k�[�"�+kC��v@�)J��J����X���6�r�Nͨ��U#�����_�dx��\�5��_7��-��b���i����O�p���������U���6Nc�d���*[S��N�<bÇ��)��FI.�\�^�Ͼ����� �=�Q�j�R(��i�1�~sg�����A�4d|P@+99 ,�l��[�H�u-�owT��p:L'o>�K��2fk���S��`QmR�W�ܔ�Ŀa@<��]�{��>��%i��ƃZ����0�G}�.'-��[zhïV�3~�I��4�B��W7��qző*LR����:z������V��5����2)_c���A�y+s�N�>bsSS�ٕ��{��I�ߓ2�@�uO����p��]�6�G.te�2yx���]���8-�/�!c�
`f7qL���u�3D�gu��a��:��L������U �g��y��+���r�)�@���1CʈO��7;fkZ�WE��iQ�Rn7uM'g����-hմzQ�.��Mq��p�כ�&�J���e����6:�篺���|��p����K7tzS��g��V�q�&5UA?aTdu��m�����v�V�z�}�綾1�9r���Z�|�������h�#�pbT�~�S����y�D��C��&v�Ї]�����N:�#.�l��1/�gsp,I�jLc}a�Щ&��=���2@e��bZ2S�'��4RX����Gk%���"�vq7�i��
��	�p������8p�~��	�1yۯ�[,i�E�D�|�������!uVō&�k0�����`G���<�o?�$x�Y���:N�
�;��(��W��O�$��UsBH���qa�f<}8x�ye�U�,7��GX��Ow�]�Gr�>I"�;E����u6f?���a4�Ä�m}��W�=/zE���)����	�^�G�Ak?����V�֗%��u��3�ρ#A\Ë��oY#d,��Y,P�ƺ�-�-3��l;��N 13d�T�I��p0Ⴘx_'�r^b�
�g��|]+�j$�/��!�7��p��s܉�*B%�:�<[�;j8!�CA�
]�mSt�J{�#{�WP9~��:�z������_|	o�7���Ş�&V���=!SksO���`=�m�8/FKT��'���}Mʦ��sat�p�-� �9�CG�#&y.Fp�z�,"P��)�	i⃡��~"���8�lGl��.��bD7�X�ȕW�U�.�X{oauL�b.ϥ*�/��<uy4 �|�k����q�J�D_���S@t��_L������L:�)��B�<j�x�Y[t��hkQbʏ��M���^�Ν\�9/f����U]��e��.F{����2��Vpn�K#쮳�������G�j����X95�%�U|��K��ⶃW��}{1^idʹv'Ni�l��<�2X��n�*[�D��Is�ٴ��ulNL7�/��x�՗�v�ݎ����
٥��*�g�@_D�˥.����@���d2�nSV��ǯ��),��A�CQ���`�ت�W�`}���1�2[���\�x+��1;�8@��m�6-gM��\7M�ﺐ햄����xZx�����Ϯg]U�}�ҕ��������t�S̖ӓ���KƢK����O�9��!;���<��5��踀�au1)���(���
��0r*ա_��@�ccin�����<����i�e�Y���1K"З܌VaPRc������!�ECn1�ka�o@���Eu����e�x�S�"!N�<��7����h~��Ļ<>�Y��GzJ�0i��^. �p�ͬ��,�)�"^�u,M�d��s~�pN|[d��od[k��L��t]�it����VO��3��j��f�>F�o�F�9x�n|�kpǵW�+?��{�4�J�6k����^���Nn�	�o��j�^��"�_�r=~��s�?��8^N�ڔm>lT(�Wط��Is'��YG.ZLW[	ս|�����b��[0�FA�`g��5�ދ�����h��S���O�	S|�*�R���#��{Ry¯�X~�v���iC�%.h"���W��,vZ^�aj�ܜ3 �t�,xǍPs��N�t��h�^��d(����ͣ����|�>�"~��3���ԫo�1��C���IZb���UWٍ�e�Z�i�E�T��l�:O�������^9&�L�6H,��3�eë.�K��ZbeD�� �3��*舲.����d,�S)g[��iY!�5x�-�Y�.k�	��>u�8��|�.���F�tA-ʆ��2��j-<����T�����5Q�q��J*b�;�[�ґ����P�4�����]A:����ӂ��P Y
hr�Фdڻ����0m����>p���|����t���'��:o�n�sj���60Su�Cv���h�Q�x�)�gG_Ƿ��	����x⍣8ڔ9]݁Q1�hWa�FQ��,{�
�n!�ɷ.jR�Fͳ�(�t�=���BG:����"5G���)�=1UP�z�2�����dM��u���7+�*~���=u�E��}�=Ӄs���4ﱅA�C��T1����$���>����]]ёt��]09cg.��1��e	 s��_M� ��[)q�/��Yx�����Gz��5đ�\v�J� '�T!�tBd!�O� �w�qX���.|�@J�KPjw�FU��"%�>�t�h�������y�0_�2������?t>y�5�b���^��jd�ޘ6)�NX�WO��ۢ������=s�6���j��Փ���z�?��7�7�<
�f�79�E��pEQz���6��@i���a	�8w,dןAuQ��xvN~Ĳ��:���hg�S^]w�>^���T��3�ۛv-M�҅�m��{Ƥ����F�j��2�Lr����ai9C��6�K_-җ��w4Vq��]q�,dH�~�֣�����~����S�������j�k�����f�I=����E���l�re+eT��Z�jA��)%Ҵ��_k��o���w���ፂR����ċ:jS�/>��6fɜ�ۿCr�ʹΧ^^]���[	Z�'�X�a�!!���.9G���٤뼼��C���[%�y�����Q�(�,Ҟ�����Niq�#�{�}.nK�s���,Ԝpy23��*I�i��Cm�/�F��'���S�������~e������n5���L:�^cMU8�sw^}9����q�����@�4:W���Yf�p��4�X�X2T�5��
j�_(�����߅˷Qm�{�-��?�S<w�ݩmlvE�x�Ka�p�ٺp�	���-)�����:ɫ[�j�(�}�`�j 6�Ut�<gʩ�l�Fm��=A�<,z&�vw� (�C9������f�H0$b�v�ߚ7�j�icR��L�۟�~���b�Y��1�5Xg�v'��.-���'���_Ouz��Üq
|kcϽ�2�r�}����q��q���
=^�J�Y�F��O�5��#7�����z�m�	�r��&�����tM�����0��\iM��Q�w]�D�n������vN���{��"N�h��tt��>��Q9z�Էǆ�H������t���Ė:$,���=8��`2�x*L�;��}�>K����Z�w=�(�� �Tj�"%��"LHeʜ�.��];�6���l,؊��p!���Uې��~�����"�!�,��m��j#pm��]��_�Ư�µ��G;��})�~0c*�]���1C}T^���Y�����ko��g��_��|�e�5�1m@�:�|���P�BY��E�(
H�Ѡ)�p�+v�Diߛ���LEZ*y�V�l�T�^xk+y:|�传�d|�H�[��"*r!�.]On�AT2Oj�U:�p��L#J^�D�u�{D�����ѮE�e�T��������y�|�fsM-�1#��{�?��e��!c�ت����
�&jb$L�{WHw��[f�ϼa~Pڡ�qV�~X���Y8OR�e��!?�� x�AΣ�5ϩ1�iߊ\kU����Jzd_���V��UVAIQ�����i�=-I��P�;(�8{��8�N�l�[��ȢF9]m�}+n��B�}˵���ᢽ���(�rj4w�u8��ޯX8y	*r�r��,�;��+�� �Q���t�0)<.�±����7����Vw�1Sy@�
y�t0j�����4�@*aX�?%��0���iNo�d�/���ɐGF�e���s�bV�dO�0ӷ#�+�v���M�[(��������x'�?Bվ+|¸B�q�������$x��&mb6�D<�Q_W���2K.q^]�}�u��&g�^t���]�3ڳ�����8�PhL�ϖ��u��@Z�y$���s��2�d^��"��w��� jU�Z�_}���&�[T,ο�E�K�$�n\��w��̌#ys�O$.�XN��V䥻��#�r���c�0K�t���ej������J�{rm��_��r�w�.3tٮf:Gt�~�_ϏG���{�4��w�edq�����8�g
�Q����z�v��(���<��)AfI��ⷌ٢����fʠv���@u�	ML��<�$������멵y�6:�nt��U��jA�eӊS���̕�����^�_��&�t�*��k�=��8�[����;��u�ͨ�#�z>�f������;J>��}�
����yt�#����?ǡ7�b����R�~�_
�/"=*��q�C~�F�$~C��9��˽'��!� �̜�?��dt���ŧ�l+g�Bܒ�!)ҝ�E{���g��D�>	��r�
��S�P栈�3���A���Z?ؿ�D�i�ВU�Օ���>����;/���W>����O��,���'�lcO�GI��B2L{ݖuߨ\�ju�L��^y�>��������o��Z����Ź������O�)��v5��Wd�RΡ��Æ]��q�ܧ2�T��k��	UV�٬�cI�Z�JY�G^��D']�kik�zJx�9,��5���3�s��⾉�_�.�/BE�!�ȴ�Ղ!8*�%gm`%��8�[AN�e^��t�)�8�N���omUM�F�ɽ�M��Z%,3�yI�D0���/���8�-�aH\��Lps͠t|f���Ӄ�ɜ^(|���L[k��n�qq���g?�[������vi����pP����g�3�禲��)%�qi�:�*���w�j�~�~�E<�������x6n�ٝ��d/�j2��Q^^(��i �=��&ÎU�"JR�4)�O\g��6o�	��2��K���=2�*+��X*y��C|"�;O�\V���i� ����t x"蕍��Rы@)6/y���.�)c��'�+�EX��c�6��O�CRX|��=�X%߻�H#��J˂�G�X�l�~�̸nf�R'�κ��q��d���h�(?D�����[%�&��sF�hR��rrH>W�)�r$ʐ������ǚ��n�-)�1=��Ē�;l�t������i��椦jZ7
�`�w���������ڃ�g�Nw����t(t��v�e��I�nv�@b4�fU2�5�UF�a���������{q�շP��jd[����'`GȐe��ܐy�E]::f��)2]w��eF��_R[Z�,>O�oE����?��n�.�t�H�Z��E�Er���(��[}�¼���#�ݮOp�`)�#��atU_���ʥ!}��Ya�ƍ:Sn!���lڙ��`�!�>�2�(���zBN.�,��"��+N.�YT0$~F���C��?�{�h��>�8=8SP\°��f~aL2c$F�v˂���y��^�J���l��Dɾ��R��i�0`�63�$����]���fF�,^B�ͦuz�����gخ
����͇Y����y�>]��:J2���\窷���D���|n2���/�m*v��-&��'����u�&ha ��|[�7(���8K:b�L�9M��S��b:�Z+]m��9}GMn�bG������U�+?�;n��^xVƫ��`7LjET�zVp#��GnN��KŖ>�)ґ���C�2�.J���x��g��}_y��8fv���Z�wM� ��_*÷s�'ә��å`�dw=l���V!��9`c���\������B*s	��h�CI����p[⸘֥�o�a�f'���e%�v��.�)�5m%9�`c ZS1q�{�*�_�U�]]s��SҩpZ��6��
N���xɕ�5r���7������;O?�o<y���:^=5qW��<�IVaŞ���zYړ��N�7���1��c�NL�S�k��ݵ=Eל�ad�H�j�Rt��Nu�f1X�� �7w��A6ĺ��H]'��12���P"���� %CC�Iz�ׂ�I�̮����.�v����+�![���uL�n=�r�	�����R��������7�͵�mVټV@�\a�8t_�*�$ $%N:sp�q���"�'@No���	�΄��E"�2R���N�����](W*9iD�]n˅3oLN��
~�cj��r�_2rе�!+�_k:�Ko���ʕmyfyk�(i'�~��1�����z�=����B�(�%NclO�XAY9enj��d=�(�*8p*�0s��8qh��N!�� ��r�
��J���U+�+V�"��S`]9@�WW������љ��j�9��R�/��JE�&�0�*��c��R>S�ݵ�t�N�y�r�Gş���c�/���A�e�"�k�»}g���^��^�$Z�r�H0��8Y�T������t����D%D�CḂb!�����?Pq��I��~�+s�H���\��wɲ��2K�5H��U��c�A����Ȗ�oNų��c:��n�|/>s�A�q�q�ҋq�ڎ&��-��h��k�u�+����W���)Ghe� ��7p��ra>Gc�^[���j<�ܫ���?~G��	4�*v�vw�*j�=A*�F��wh���1}��|�D����c���$k�t��y����h�)&�P�1�@T}p��gC�u�(_�Ԛ��xBH��2��1��t���/�B�-Vv-V�ʣ�i/�b�۞�ٲ�w��q3�����E����>T�J��8s��{`f)��IЮwi>���|Ҷ�  ��b⦸<��qʹ����Ҥh�8K�岶�w�H���uX��"g�6�ԅ,�j���t!�N񡌖�b�	/����wVzMNQ������J��l���a�����ǃ����!8��E���G�������)����~�U��n=��O�yK��sR�sRX�\N�_E��!�J���˼c|�������*��1b�H����c����l��'����p�ff�`��Fߩp|�B�|���mb^�kw]w	>u���������Z�6��U(t�'�O�5��
@UU��ti�u�׊;� "&Y��G�!�8�L�?{��{�0�~����O�&�h�N�����f�1O�%�N��T}D�qC�ts�nJ�2C����� IS	���!�D̻t�)����N>���VH��__GXX��lYP� p�ҠŽ3����UO�!D]=�gu��
'O��n�n��
���d�~U:Ȑ�O�Mu@.�1R���F1�����O=��>��}�Uz�$N�Ͳ#�N��X�S7�4�ז��dY�ڝ�dN�(�Ƽ��kZ/p�t�T���Xr�:;_��h�sG.d�Y�V�����	f�ai�My��W^g�Z�*>�#=mD�#�an0�ېs"�j�ҿ.�Hs���9Ǖ��R�/;ؖiD|f�$�f��ŮP"ْ�R�v`SG��=b�N^ϳ33�ɿ�`3�U_�"�i�e�`ĉe"�J�Ha	:��@BF�&f^k9汢酦��A��|=\�zc���Mrޠy�j����t�����;|��#8� �S��W�(V��7q���F�_��Y3L���a
�{ܬ�J��bE���Z���-ܗZ{E��RP`E�bA�"U�8�~��NS���sy�o�Cd������|hQ$���xt�:Ǖu ��`���"6������u�Hw�mg��e����J�p��gRNtA�0�hz½�b.�W1��� >̠����Z*m�d�lIN�!�"io�DQ���4(�����&ч��^�t|wj��*0�*�QK鍬�� $]���V�:a��W����������K�W_qv���4&T��zb��gZW�:�K�u;R��d�͂�ty�j-��1���/��?��w�>���x宝���|��č�:m��hVΕ�e��uWI��dDt)4����,֣Ӕ�Ms�L6�����SW����aV	s�Y;jg�1kw�<a֮0�Y�i���ǲ4�Ep��I��KԶ�u����o���\�㒎Qθ����~����~i#�¤H�);冹8�]�k̄*��R_���|��w"]Ĥ�&1�l��J)u���c��Z�Ї�%�uɧ�e��������e�2Qb!/_����z��yS��xٸyY<0���]�@ �,Hix���Լ�b��Ƭ0Ϧ�����x�nwY��Q�:�""t�������e�܌��ꀫ}5<��H��T0m\� �(�ݷ�c�s�[rҋl?�)�K�Rʯ��ª�7�?��GV�݂[��/���Ō���O����=�t���w߁;o<��^��9��KH:&NE1��hg5/�l���F#��\
ј��7$#5����a��R��;���G�¿������O�X�xe��r���ȶ��S����sQ$�"�k����[�8Rs���WΊ����UR�T���ʋ�X<�l���{V�J�mGm��zO%lTyv.@��z��8ō���F���/��;d����(�e��n�	;v� �S��r�0�k�k��S���fָ�·AW�I��x���
|���ULVV��V��]Z�;	Ğ�Q�6�7��`,��[�WS�G�����r���������տ*
�}Xx@!%oG8K�>�:�=���Ap��S��jl��MF޺k�H�h$G�*�K�ZˮcE29]��ğ�6�����?�C�3We����)�������|��(����fp��M�u��ۑp��� `i	*��}�G���e�D|B�N֥��1�o�=�-�h��ѷ�:��P/��Y�hR+R"ͼ����d%�4࡮�������G��=8uJ�u`:]7j%�c��]�Qcd=9��QdmR$�d'�O��� �U�m�j^L���cظZ�~���2��D�q��� io�Ҿ�b�:�"��3��&�iI�b��sT�x�K'p��mP��L{�O5����+}�҅��Ux��U:v����N��]+�}�H���p��3�(��<S,���"�D�݆�`�
F�D9�x�q1����f�Pk�'�K�B��Վ)�O�s��gBM��dMʩ�A��8/�2�S^)Y]ݨ��������;���/:����=��*0'^T��K���H�D%�}��5�Z=�ħ�?��q��s�9�?s�GaT�1NL�x��+x�����c���_��N����;�����ɳ��5�nhe����V�,�_�"����yVKNDs��[:�u�B5$�Â(��+SQ6M:�D%��k���'��3
�y���J:y�NԹ@��]�x�f�\�;6��</�~�m��npd�Z�߬���0����i��~Y�\/�l@ogeԦO��ZD��[�������=�U�Y��J�ϛ&�*+nA�B$?M��ȅׄҳj���[�}��JY���"��	T����\�Į.A����+�Y���8qU��(�d�
�:Ғ~��oj!icc�!��v�. ��#���T:o�N���H�e'5���JL	�4`��)=�C����j�i<@������Oq�B:�I��׵�����X�Zċ�J�y5��c�i�w,��5�+����=�C�lY6;c)CM4~�����ވ�?x9n��b��cG��T���z25�e�|W�0:�_���`��xgt���N�[]�����g����)�s�	z����W�ى]����|-��*E۫��w�Q+w�[���1�����aA�E���q�A�3c�RRu��6@m���Y�l��<?���0hs�����RX%@+�,����YǴbH���4��P��Qvjv7g���+ㆧNjg�U5^u�DQN�Sպ��y>���ȩ�u����M��ؿw6NǦu��\�[�WP6<�0k0���]'k뭂\t�k5���E)��q�&�@�j�IkYO�7uٍTf�F1Z��i�l�&��^~�k�s�RV�r}X�m��q|5��>�HB~Q�����?�
�Ê?�v��=t6�!��'Ah:8^��� �1����,���L�98�P�$��zt[��U�C:����ls�'XY���!�jH�vJ1���W�I��Y�`����?y��r �Szһ�sy��N��^8#Q6����������M`�P�Fd�/I˒��
�t�u����}+�`�[���;�B}MY%����Α���Fi۵��;?z+�t]gG�9�'^~��I<�܋x���pl2�iK�#���9b4���&����&v�pW�h�4[�pFS�t��A���F��F�>
zv�
�|����"í��������Ex�/B2��k����B�R%g�<��:2�����("w:y�&��9��h杵�(2|֊��L&���]��鍈��lj�+��a0 �*5vn����H�i�0_BuD�TqK��|/0
"�ϝ ��B�ߑ��
�z(��
s`��DY��S�C�� �2��J�v�_,f>��\uؕ�N� �:�9y (���W&��_���>��TNvd�tR``��#l���`�;�KDΡ��s��UfO7�깗_�w=����Cx�ŗqr2A5.0�5F�g��
{ea��q��N�R���,�w/!�p4��������;���A�
Ɋ�x�;�xHCؽ�/lr�ό�i�#~���=�#^�I�l�9Y~ʻ�vIM+=^ʰ��J<��kl���eA>&ߦB(�q+��������4���\����9�c��W�?m�u��c��'iW>_�m1���.}&YӢ�;�ŘL��꧒O?}�����q�%t�x	RE��
��D-�Hteg)XR�����Q#��,O��a�<xa�����A�u�d�Ho��ʶ�O�O��y0�T�V�5/s��.'���sv�vv�j$�⹦��Q'ɹ!y��s6K�P~4&Z!۟��6�@d��8��Vԥ���i?瞷C��>g�V���u�D�<���2&�����'���@<��-蠝�.���q��6��y߂�i=[�x��=֦g��%/J��֬�h�:r��"����`����_��e���vk��ݕ(�кyހ�zZ^�٬ί��}���-����/���:�L(����6g��'7��sO�k?��=��r�9S�Q��9�J�����������y%&�制��O�~�Sz֊�$�N�[gCD�h�RG�m�d�}Aθ���)f���fa��]�r|)�H�y�8O%����ͫ�a�P=�RM�Y��P�x6`o4�"b K�f,����ر�5��}�yV8[Pm�A�f�/�=	Ý˸+4KJ�rTb����K_�<~���~���_x�}�	z�U<s�M�Z�����r�R5��J�
�I��!��մY��WٵZ/4����q|]'�-m��O�:����aKd�D��8G��=8�(���Fί�z}���짶���Y��v���f�SŲB���x��ٵw���I���Y����(̲e���"0a>5���2F�gnRo6��7�G�{�9��&���z�N�������U(R#�	mEa��ő�d�L�	��F/�L0�`� ��O������Q� �G�z���{���X����HD��o�*�8�|�H�*�1٘�{.��G6�E{w�}��۷_���z�~���/�g�OA�c�f����a�����[�v�`�&�&%�9o�S8*�j��W�E�s��<pV���H�v��a!d��w��.��� g� .K͈骜(����j`݂_�?Lҳ�G��9��"���,#�"�&U����F�\$��IG�D�G[���!�� �.�5t��(�����~��
��ۭ6��t˨�0���L��Y�������.ҀnΡ!8BT5?��B]y���,�k�u��µ��g�8a�v"X����zb���Zз��3f:\USk_4�uV��*��U�v�XӸ�Cv���G;�0���ϊ����3;ފF��n��ȑ���_����#8r�$F{�`׹�z�5��ԶS 1Jqȷ�M�kɂ*'��IW%:�>�j���\��8#,89U�o���c؞R4�ٸ�Z����Wu6D������x4*�g��KN�#��bl��f���Pq?l�Ldd~��ק��cMN�:��ۏ2n*���I�mVi������m����4W��<3�)�I�t���-*�]�*!ec�� )����UO�\���J�Qg���1	6�s���"2]1�����vr�0�$����V�.Z�c1��t���4�v%�<��o��-��
]�~�n��'��dW�?�G���ط=f:�kȦ�9Rʟ��t�N���>g����A�7�������)d>!�g����(�EL�dz��!�(^p6KǢ�4��+
$��N�V��H�m�F�	|Ė�"fR�Q_�������Y�0γ�~`�e�Vx�Čͽ�n��\Y��;Q�v]}l��-l9.v-6�����CoCA��)V��t,w�~�7Om�p��7��������au�������2��>���}��XGu�'��aI{^��^�	wP$�e~/
z�M��!'�f�����Md{�U��P>Ky�<v�~{�{4hwj�����,[)��CA:�߭x���eWD��Y��$^T��ȇ�^$����yd�u�0v���o㗮��]}���[>�$k֪�'d��hP-xz��QM����v4�F��q�������?���x���p�cO���0|�ޜ�&"V�i#cL�#Wk]�Öh%��Ew��+�����0���sX�.Ҟ'�/E�ͦ/tX��VQ	٫�o:B�qm˖xԒ���LUZ�M�3Xz��vG�!�GѓLK9+����KR��#�A�>�iYFHu�`u��Ha�nO���V0�iyI���Z�
�����{v ��f�vBt\F瓌,Vf�!�=gl\�@�H��6��"2n�=h��ڽ���B7WI���	�g~O��C	%�CX�g�����  �����N����VVw����m4I�����4��Rީ�H,�� �]���m~�$��2w�U)PMK�
�F;�n�go�	�}?x����O^;��Nk�v��X]�'Ԗ�_9P�m�6JmMDowq7���%�.�s7~v�Q�}{��&3L�wE� ;ohG8�o�Ɉv�B}�z�aE�� T�4}��Y��
9Wa�Pa.�:
����Xq�|��#�����o��7d$���a!��2�ſ�d[%��_t���rx��ZvH�:
PӜ���]9��q޿���:�Z	Yo����������S^�%�R��i�"6�ʹ���_Y�t���=��9�i<4)�������i��tWy��&�'�Ze#SLE+T�kj�ʟ�b�[�B;-/��V�Y_(�	6M팙娑/
G�uϏ�_}�A<���X+Q�\����Xyd����u�QI��I�2��r �)݁�ϝ�R=#���G�i�������ӫ�9�g�"�f	����z�s�ع��Hd���m�\�/0�y:��G	5a,��bX�Ț濕����fޙ�/�0�"��;�ݵ�d#BVf�n��w^XT"�Y�Y����ʙ�Lq��k�O�����/,Ҟ��m-�IlK����w}u��l)A�QV���ܫ\��|O�À�Y��� i�*����˜|�3F0��|��ds����y@�c<&���*P�&� /;�f�����,�[��N��)�!2�k�ɼ���Cv�
^_�>[x�����٢Eu-&u<��y�+�������2��[ES;�~h�&'N@>���eGv��9���ȃ��b��YBj�\����:E�w,yV���T;+��at����m��V�+'NM~T���3j�&ݿ�"o}*\��j��X�vx:�B����+�~j���t6hY/�&�Q�S�^��g��+�{��x��ۘ����/.,�D_[�Q|��^��*<6���Ց���k���z���V$o����xp�;H����_21�	������*���{�^���<��)vT ���ލ!] ��VW&g��[w<S�w:�����DZ��9*�;�)��b��-V�ܩS������������@al`�!o�Lrd�-(c�S+��B���K�4�|��8e��n��n^\u��8��;��Ͼ����G�7?y��~��K�v6��+V���S{J.��9�\U\U�K��(���uZ��H�OO�q���d�[�)Y?����k^G���s�|�.�l����#��h���a���`���#�_dx�Ux�,�t�����]�lBڊ��4T��o'X��3�������ʵ^h�l���)!�m]���Ṽ�^�A�����!��"x|���)�־/����I��y0 �+'>OQ��+j[`��e��r��	����x�-��ݟ���k��Vwo������	MW�0đ���8A��v
�U�j�X��y~��q�/~�c���7��?~�z����5``��+���j ����C��P�Q�f�L�t�������:(C,�L�E��M���ى�-P��0E�q�� ��ؿ�O�6����<ʚ�F>�R#�9��b�ѐ/0��vR���ѝ��"�1�@dj:�a΅�ECw��RU�`<{�<��d/�%�M�q�nS�<��G{Q4t�z~n��I�n"�AYaCfj%�S9�(��#Y�QZ��d�Q�h��:��P�"�@s�+{���T)�n��'O6�e��8_	�3Ue�3��n�h���7�ǝ����A
Ti�#��j+�\o޾�����|�z�q���K������
�F���[[�6\��8IAg�/-8;��h\��~��h�?z�ʜWDUx�e&/f�c̘�!��jd@����d��UA"2���Є2��L�
�8t����s,��/Z�Mw)�L��&|bh�m�s^/�ℱ��+}����2���D���s�yUA+LT��.W�������6��>!~��gOViHE��uH�ѻ�g�qe��*N��@�λ����׎��RwJ��tѐ��%���c:D�9d�2!m�f�<ա���;$h�K<I�����~�qr���]6���+^:�v��S[`Hi��%��__���YD�O%�O��_�5>�¸�\^h�
�[yiAܚuM4FVߡ�΁�-���Kt�P�{�	4����	*��������}9f!������*��o����)�i�)�����^��g����?}����c����ثo�mw�!��F�)Kg"l��4A���W���-D�'��{26��Ⓥ丅�M���(\����Jd���7X9�ueP/��~[|�vn�u�_�ξ9[Iz�y"B��m���:�[e�����0�+�=/�|�x(�����ߎ/����;qh�4�������:��G>���O�(@�3���Cu	�Ij�"l�R��-�Oo�̴¹������������}�<�2�����Ρ����wp����+��^�U���{�*	�Z���p<��Aс9}ϊO��]��v���̿%-Hz�u��
!��IdB�����"qd�H�M���Y�>��5���=	 փZt�ڝ���H�'Oi1���"��:��殡�ۓ�~hN���z��Ovt���dϜ�e{nq��V	U�W�YnPK,��͗yʝ'��b[Jd�P�uI����2�^�B�lc�X��}��4EF�<	e��!���~�Ɉ	1�4�i\�(�T���|¹��+Q�nK�9�2²��F<:^ſ�����K��~�7q������t%mk�<љ.E�W�  ��Itȿ����~��O�T�����.�|�.�t��{G��7=��<�<��Q�z�M��( �v7�����d%��dT����w �^�i_��Wb�y'�o�g���o�Ҁj�Pj�r3y��)����u ���"m�Nu�=�0NH���U<���9���)?C�oFP�:�)y]H)��H��H�U��\�D���������U��%ElV�F>�M��R�銓�C����dDRu�~�A�i1�0OB*�3�c���X���S~����R��jP��U%�:Q�g*��j�9sOs����7
�b�7
ei/���u�������2w:�]�Żgx��Q|�q� �\{��9�\g�jA�u@�V�?sb�yoN�P�nh�Z�N�@7������?��>��v�Cx��F�^�'D�w�Uv*:"X�S:���;[#f8�� K�3`�.\��Aq"��f�&�+�r�M�E��d�;?�:��uh�,�d��~,�7���Ӈ[g.��.�y؋�+���=1m�2���:�N��&�FŃNm�T�.L��q���ܳ`P��ѫ?�Ӥ��g2�����g��t�q#����Rg�8�,5�Q�|�;0�9�����ɧ��b�m�����(��N�&��^ӂ|��B ]J�f���M���*��}*�,-sz2W=�lL�A���� r��9ӧu��ח�J;�� ���R�\n�m�G;|Ȑ'�b������C��O���q�}�nl��]���H3Hş!N��{�IŦ�Tg�"ZT	,@La7k��/W^T��aB�	�v�X9le�[���)�9�X���hV��
#�S�x{��o��+c���m�6�:*3�w�O�u:hA��xa������4V*�o���XG��9rL�����;��S��?���Y7ִ;0ڹ�5�S�����*�3�wM�q^/#;K�S�}-�8�Y���$rFG�y���!�® ��bHm�l�%�B�9'�l��w�Ҿ'�U;
1��\�������q���)�6ٵ�kI����/��b�04b8�V�b�q�^�92������rNo��ʢ���T�C�
���+~�9�ޯ�
���9��Y�1�RY�YtZ��������e��(���V�Ӛ
:aS�W₵s����'n��_y������~��o�[M�r�ݬd��7�X[TpR4Y5u���@�f���7��X�rT(6����r��7��lM1(JD�q������#.�Eb'��W~\|[}�k^~��J�3:���\Z<7e�.}�_?Y��x��ġ�i�N8Ӣ�޶�Eq��
���Ya�8,C��@"du�5��x`Z��ZX���ٙc3�0ǎ�����$p���*�����?dѶ;Ϙ��a#g��=����;�U�!m���w �7	3V��͜R�S���j�,��V��5�'矏�z���g��t���O~����6�ݴV0�R�Mw;��'<�� S=��v}�ݛi�I�p鹻��O}_��Gp��#���'��š7�Ɖ�T�Ȗ5m����i�6*s=��vs�^�^+x��O�;fh�ΐ�#��F���D�挖R!c�sP�����29GV�㪑b�C��бb#,1�-�ʰ<��BP�U�W���ŉ�e��E�]n~����F�Ἠ�8���>3�7��0�x�p���=i?��뭬�o��F�#�	�W������E���
��a��[<H�ٿ��?����x��ny��E��i��"H�N����$��$W��&(��]���[�3�/gCBu�M�/ߜ�Q���4�iH��9�ᎃW��č�_���ۉ���X�z�U7u�#�$e+0�y�ҵ%d,��)��5��:�+��1���S|���q�O��7���&�hu�=;�}��wL�V~f�Y�
��Ap�����h��VI'�\Zi����������?�+zLN�L�%�C�8�\8ˠ����$8��:$̋ks�*ó"���56y=4���3P�[��B�Ⱦ�:�kH.�7�]����c��z�-���i6U.�GM%�!Z�pm�� �s�d1]�%$<m���{��4�mL׭҉���t$@��D -�ӳ#��zJ^'YG��ߢNQ�AJJy��X\������o.R�m���M�����<��.^Ԗ��sdG�ɣ�.^B>�!s��wCd�B�:�v/�At9Ut韹���u겁�����>��D�Q7�<Z>IUJ^��9��vLhWC�\��nU�S�z����h*C�%���Yv��v�l��EM���g�ا%���^K�V��j�_t!��Z�p�%���}ص�bo��S�د:k�������)&$7�Y�ƽ0����q{%��Z�}��KG_�w�)������_�k'7P7z�xǊ�w�m��]/i=GF(iVQ���l�i��7�G/�K�ܡ�@�c�����M25R=�;��p@`�˱���٤����<������� E��1y�4�C��ɫב�5��S�����ݜ��r��N���B��	�,Au_#�Н8����:�sv������X5ܕRE#'�'Gw����������w>�i|��Ǟ��6��	��Ef����Q�Si-�q�����~,�	6O� h�`��Ss����{�`���L��SUw�B�H�� ��I��-�"*4ɚk��-v��~�w���G�~�x���xF3����[d��4@	b!H$�~�:�˟�g�<�Nխ�?�[U�������ވ�����?x��~�_������/��jgDA7z�2�D����e^�li��\�YG��9ͯ0W���b�F�|����ˑn�MF{��� g
bDB\�лO�/�J7�&�jv9��J$/���q�pLg?">2�a��Ѹ9>!�MQ�B��4K���/�� ���>�!��q���>s�����	��ʰ��/��6�5Ѐn�����V<�ߥ������J� Ԭ��s��V3��H7���'<Q28KX��hmu[ /���(��g^��c�h����'��;6b��n
����(j�(-�9O����#2�2oVX�^L�1���������b�ݛ��/��}�>î������/�ƅ�.G�j!/��Y偣'᜕IO��ᑄ��a>�������G����ޕ�+��7Bm>�X L"��,a��W�,DPO�jR
;:p�;\+Kk���3�^��=p�V	/���_Q��6�v�ʆ�q���=!�����V� 2�䫹9����TUsӔ�s��H�2:�c	d)N�H_ϧG�F�_�0�r� U	��i~�O�c� ii0�Xs;��,���l6�{u;L�ɬgqlK��Ư]dWsl����w܊���oل����S�01��R����� í��:#�{3��D$\��<�h�C'��ڵ��]T-��9�.�$^ݻ����oN��455q�*����Up�a�:�x����6fAK��eB���8c�#P>�z AO�� �4����l�Dk�+4+8�dhʏ�yu�j!��QX��U�)#�qѕ���NƲ��/jq�x�T�.D5�mR�b�<��OF��4�u� gk��9lܢ�h/�UA���v4��h�,��F؉%�P�#`VBށ�I� "�]�yp���E��3�J����B�R3djޢf�*H��t%:�����.��'*d�kB��.�蹉Ƕ�<p\e��Z:���Ѽ	���a� ��e�7>�~�E�%��{�I�J�"��@��!Nr���/�C��I�<�/���뎒#����J�g�Z�U���09l�i5��<qϝxx�]�ㆵ��L�gH�E*󄊴�4�n�=0�C-la�F�R�P���g]����C��JR�9����Ρx������1��|����	-�e��;��y��7�Of�m䁃Lx��7�O
'�}�����ey4)Kpy�L�Rrz5��@L��c <T�?��ǵ��I�d�"��?���,�9tb^Hsk�>��=�.&QrdM�Di/5��c�
&�T��}�z[�K�+�jK�p��I�yy��Un�!�f�g/������v��K�>��?��q:�rS�k��ϫX���F�]���D:?�=g����V������6������;��?��Y���8�:�	v�)>;w�9�$+ooNW�y��\�*�<�:�@8]�����p悴c����g�ϩ�>g0�k��`ܹQ��MS0:��,Z�ku�LG�/�'��UX�p9��c���Iv"�`������d@׫Z�����]���{���#=?9(d���/mT&����8&X,Ҝ�m鏙1Y8T��ì�}�7��nE8+�Xw�Y�3����M�*f��A��	�?6�0��Z�Zb���}b5��06��ѹ����ދ?ݽ?z�!<�v�w3n]5�v��B*�S֨�2ȷ�A�an�vE���.�f�g���u�i����x���8�
�}z��ُw?:�ç��̬(�Uԗ/��y+ ;y����r�*����������x>A&F�+Xe��0� �Ĺ�o���V�2x�"�\�[7�*�ϔs˟�k'����択p��~7�x�V�1E�0�`)��n9\}���q���l�:�=ܵ�3Yw�-�u_	�}���vO�|WX;��vՇ�m�Vh����:���iOJ]d�sX[s�ܴO>r^ع�u;֮^���0�-�6p>W���a����=� Q�k��,s�z�5��*MG����S+å�Y��K��������f�t��6��)]��qbp[�m��Ȝ�d����:1,��
�%�1�@��6M���𹌩Q ��=��5ޛ u�3!��&���n3�p��4�K9<���-�!3T# ��_K�䪆�,�׏K]=}��FQ���3H�I��ˣ(
�5��DM=Mڰ� ��E:�ʸxl�T��&/�[|4���&fN�rC����
©La��k-��n�<ſ��]�b���[D8Cz����@t�V�{H|��83e ���ɵ|�ұc��f�*��kޚҙ��
��(��OG��E���o�p�gʨ!�wt\~�#2��P�L��9�<ؿ&R�9���\��Ɯ#�&�J&j�Ϣ=��-��mx��-x���ؼ�ft:@w^봤l����x[̜��V��m����H���De$e���5U�鋗p��c��;�����p���d��Ě)��e��,3O�iOV��q�ՓJ����`�i��k@фma����p�V5�E-v�2��W;
p^ڨ�#(�)n��n��x�����gY�# �cq�8`��+'"�c#԰ a����ۙ�S�#}`LT%�d(�Js�437���t{�U�Ο�ޟ�������;���۱�;����ϯȹ�~(��,���W!��4��������-G�j�sX�K��<�E�]�n�]O��o=���to4��|���O����8�w�V���E̘�v��u���X&27�����É&첓�yσ��o�.��#a�%.бl�t�p?�"m�sД��M�?�	��dgC�K�N�dG��ϊ��¸tX�AY�*���e{>eppO����-�{��#.���Dk��3��U���8I���
{,�:��l�}N铫n,��u�~���2�p��@�	~ȡpd�]R�%��~N�a,�ɓ��=���]��Uz=�&f'é"��ڃ����y�j���6���G��΍�P���4-��9���0��'$��+s�F.�<�AR=g�|���i!����xa�f|w�}8�vr��~|��7�e��#D I v֎��I(�#Ҽ� �~�3�f�G�C�.�K�l��L�lIϴ�^�-���A%b���ޕ�3���S]zE����x�ï����9c��G
�+����{{<P��j$���0Z�+�Dy9&�a����=��k�U.p�)\Ey͚e�O.BP8Kͫ
���f�ϗpq�)�xxA,�����}�dR`p�ɭ߻��qbnq��t�$&�9�9��3~~q�N<��nܴa�ư�ƙru�L�"��s+ڻQn�p71,핆 ᎖��8�j<�[�:}ϸ���['��
��{/�~��>���EI�@|ӌ~#��yLE�RZ~�4>/����A��-V\r@�)bn���Bv�|�7B��yՖ�e-�r��pOP�ږ�Je��u=�aE�mU��*�(@�l��kOx�4�+5Z��WS0K֯�R�@��E�Y���|�	��&<KI������5�C?��	Ȋ��GS��$Sg"m�2��_v �O�Ӝ���q<�Bۖ*�i����LIB.��@�Nq�b��<a��K��U�ɍ�����w� �4ܵ�DA��&j�ߓҵ/�'d-ni����aX�<0E%Z-}�jӿ���"+�1 �ӏ��c\J�t���{`��2D,����o�����M�<N��}e�!V�?1�Mf��oF6�C)����[������Ƕ���Ç�3�m�ֻo��L[?���j�ǖ�u!r�>׆!n��T�J]�1G7���#��PS� =�e��/k�!����9|��Q�������O���,�f&u|k�}�E��=�b���<��j�����	���wB��O<*��z���W95K�l����&�9gN뚁��.T�j����m��[5�Zu櫌C�ð���ډ������.s���=�o�ߊ���k��)���jԪ�lK=q%����l@���3�Nv����x���~�*�p#~�����m�v�F�^���S��V�΂�r8Q��3��6�~ņ����tvs]�
��qr
������'és����}��)��*�(��E�Z��[�fHm�OVn�)c.��������>�%�Tċ�F�
0�G��)�mo4���8�b�,��x��['�t���$Ƞ=%��"y�J(m KO[�"�vwɎi<��B�oF�k��j<p�u��l/t^3�P���21��S�е��$�[nX��R���Q�rV;K�m�h���n���i��OI��|@#Д"$6� �*����DT���KYz�,�қ�3�������ޮ�2�̼�W���������r����c��G�_�w�Z�Gn��`&������u7���vgs�ń�-��$p��KU���c4�Q�5�H�,Vw&���;�k;���Й�ׂ����2s��\�)AW�hf!�¹��rmц j�2a�X�ZK�@[��@�9Ei����'�JԐ���pO� R6De��H>�6��r���{�)�s�"�����P�p��V��i/U8��xl\J�j�Q�����\Ii{z�E���Eb�FH	�:s7}��p��
�!�>��~,JM���)6��M+��q�չ�1�r�3ܡ��Tʻ�Ȅ��qI�/|��`�@X	{��ɭw"�R){:u����.n���s;���؎-�py��U��Z���Eϔ`�ڢm�p�
xd�����1c����	W�ݤ7d��������l��:�W?���~q
g�s�N� �Lb"��f�.��P�F��]���c�ī�v���C���x���[�������\�����,���Z�"c�n;z�x���Ã�l�Ɛ��D;(��b���/�)oL�x��!�(qX]9�N��6���鱅�]�ϣ��Bק�����Ѡm��9�Ӗ��ҎC�:LknPh���˖Y��`2�EF��mH�EZC�|��|U���5�6�A���#��D0%B�N�wj[ܒ��h>��$y�Q-�X��Á�*�lsąF�',�ξ�tɵ�١׍���=��6�zb���e���#�/+�����Ų��pbJ��x֊}�2.K�h��#Z��E0)u���Q�'��T���\��&�|Ff5T��L��I�]�dS�%Ӷ�9��q�Vѳ�>�����7�g'%<p0^�.�8�x6�� .��pP^CѼp� ��+�i�6D{ހ1�0�=��cK������Hs߆u�����Ԗ{q��7a��$ښϔ[�"�<G����m뜼���]��=\�a^7@�~�#��^�#R��Wן���]��w���;�=�?����R��o�]�<3�L����2B�� ��iV�1�'��K��|�	��7��H�l����h����`F�r�6UQ�%.u����p��Bw5�����K���`�E�BR�*!w�� ��hNr�����y�r�R��p��Q\��D8�v<����g�������)I���I��z�"�Ŝ/��xUh�+C<+4g����-7b^v�^>������]�o�Z|g�&����vםX7=��g/U�J�a�i�;�t9ֵ���_:X��W�d��h��y���5k���?���}gϝ��SӺ�:.�tE�	-pۼ�lRm9sEJh=j�i'� 2>��$�֝�[�O;A4q��N!4�����3L����/!E$#Lvⱥ�[�h-�h��{$^/�s�꾰���w�{��]�у�KΙ��i{u����5�q>c<@�s����7�:�X���<X���8d�I�dqB[~�)pE�Ҷ��\�J��'P��p��U�L���C��\���>�B�ʩ0����$�\�u��$,3f�0�T|;��ڵ�|�����~��{�Z<�u3��cP��''�iM��	p�&�ҌSB>��02`O������r~���[���U7�;n�P��$�#�c��+��}���k��%��if9��2:�l�2\i��?��-hN8����a�+KT�b�9s�h�DL�0����;��^�)i��`׹hV M)��x��@;�0�A�)�X.4�ס7�X	�΃���c��cň�j-4������q"9zNnbPR(���I��8�&�(�Zpn_�h# �T�X�K-p��.�g��l!H���<�<��C�r�-�I*��	�+�$e��3�b)cu���3,X������o� c0��gF�?�_��g/bס��7�>���é+]d�S�}�VA'Z�y���c�F�(�@U�Kb/�������C����9�,�;6c�d��%�:��R���F�ٛ�!^Z?>�C�l�:<8�K�I`��0�	^�!�:��
��H>
�2~s�"���$�dU��Y>O\��~s�v�s6����8����6(T��+��Q�啃u��V�W4�l�9`J�K�}�'�ou=� ����Q�>�"�G%�jJ���x:��p!�`P��f&�%y}1��'�*#�$�a���c�Օ:�w����B� 6��ȌCJ���'�3t�������ٜ��VS�+�>���psCӪ���y����=UuGt�F��!O��2�?�i"��� ������렴O�X������]J6�����\��&f�X3?���ی��y
߳	���`��w���l��w�e�n�`u;�~��L�Ȥ6��7��FG�gd�T��*�FW��ã_��߾�N�ť"Egj�&>�<�b&+7�Y��V�E�n�@2�p�!�&Ô�hmE�&�jT ݇�q1�N��kL4ْvˮܪ8y28����<�pX/*��|ӌ��G���Ey�	p�B:/�k�+'���h�(d�q3�k=+��%�m�Rs��И��p?���+f��Uŧ�,�ّU8�>���l+�[f<�_*����v���׮�x��x���x��m�r�-X#:E:u3Wdn%Ƌ�_&�U	
2�齾t�%�b&ka����{�:[Q���G�
���g0� �_�@IM������"�o�G�r2�:�!�t�{�V�F�%��賤���@�sq�������	Y�`^E0&$}��,�Y9ǃe�G�I�3fD9��x�F�v�\1����1|5_#��Yַ׃p��3̈�E/���X.����7$&����T~L�G6!}	KD��Jw��-.T�´1�tl��r�.��̚��\��ŏV�HU��99��g/a����'��½ko��݃��cضi#�D��W���]`Y��ۑ��JI���&)��T�Ɣ����[�\z � ,3�L������i���T�.%�������qƵ�p�x���u�����{�_
�N7j㽼,�B%���Zt�a��iL���Z�y�c큵�+wR��ܣ�XЉ����n�_.�r�f|`�8���V�3jhr;���t8DKx�W��-gMJAw�)�$<�ɃA�e�&MY����"żD�I҆¼���om
�����ww��/����#�b��5�R��GZ+|��=�scag�_[ᅌ�F؈�g���"D��q��BT��y'/^�{ū{���r\��=�
�'h��ί���:��2���f��݀�'݁�+&�
KC��̈́�IQ���s�׌�G� &�
��AD��Z�.�TQ"���� ��j"���V^L}�?F�3�1�D�OI,ހ�a�i?��t*P��XZ�Z�$�2��4�5��w�q4�_J$�`�u�(�X��bm0Uq���To�Wv]��A4ci��he⻬��P�B��V4��>ur�WLq��sY>�>��+o�5y��Ks�nq��Q ^eus3�4��M�K)��l���g���a�~���s[�r�ESPŇ�Cc�8��a9����#�l����q,��.M��(,�8� ��5�r���ΨB]\R��U�(�en^�n�ܵ�ۿ�n���"�,0?o��[C���g�&֪-�l$5�iĄ�72�w8�La��rF�-�[%�(��(G�q��Ƈ'������wｏ_}���0u�j�Z�����Z /ܫ� =i�.�.D2%�<��i)o��MU	m�B�pc�<�R��\Bx>̍�����w��2_�)g0,Y��g,@�1���旧���iC��>�%���~�y�o�Ǧ�ä��"�!�W�ks>ʅ=s�ѽ��ʱF+7�X������r���E������׾����q�M7㥇�ǋ��ĝ�ܨ�5ѐ�3�.��0i�ZX8�@F��aiqrn��J�t��%�\ҥ,O_��*�TE=]��]�Q���E1m�Q���t�I7�<��^vx؟c��V�FP!>\�r���2��Wu�.֎�nV
]p#9#(����E���{P��|X�+�x���y]{V**]l`�[��k�{�@̈��(�gK��>�J��8���A-��ZyP�S��B�q���|`��Zup�2Q
�^9!Q?�B+wi��J^I�1ׇe:���gDr"m�%w��\a���+]���䝏��m7�lŋ�<�{�߈i�C�!Z��qf�_��;R��~:�[��p�cy���4V��r�s��/k�C��Y%��xo޸�V�r�c�7sM���q�y�`�'<=��R;$��'����mf 1L�2b<<c7��BX�Ҏ֛�̇�/=;½�8F��Y�T7z+��6B���C4Y�eD2��������H���o�!���ܬ�Q�o����y��.��_�x�7�%b��������^DP��A#��c�P���\�
'x��7Ӧ�f��������o㉭[�a�B�*��Lk����F������`��]��`;���{�zJjw�+
;}�
vt?�������t���m��E	��ѱ�)3������9t�ºq��S�9R/���9fA�9����,�"�+P�FlNf��pu�܄���ĴV����V�S}�ˋ�C����./��CU�J3����x�j���bky<�\�q#R>+)8DX��]\�3ゅ�g��˃�A�l���O��2oc_��5Y�>�/�l0oXM������j�j@Rm�	b��^`|�Z9��v)߲�q|P��1�]F������y;�G]��YHi��G���VŢҦ��H��Z�pZ��`��f��fo+���b@Y��#oD�$ӳ���	��xw�)Yz&�>[��d��������8�tXAt�_��e?.^���;*"7�U.�o�����|��o�7NNh��J_d�g�ͭ��[��\0=Íl���!�Gh��o�jo�B�i�PkW�$>9�^{?^���?y
���v�H��o���yc�n&�<��������.�c�$C�g��e��s��IKn.d��<��������C�O���NF}�ښ�o֠�	�1pM�a0�F��k���tH��1�)ƛǥZ`�b��;{���[�@
�zz�Oe.�.KyZ���A�y��Q��AA�22�*}��.�~��%���^���؇�6݊��>���^��z�^�,��"|�ݴ���elsG�p��^��3��sv���7z2��4�.6�:��Pg0hO@_�U��U�9"V_s�I�G�~��n&�XKw�b��3�cge�������x>�.��h�e�+�[�L/�iJ�y.n��ɮ'�~lV*��=�Kp��Z6��I`��0��P��Fi+��5��e_'̍�T4�J�� �o�p @z��ect�f�v��*$��`��!9"<�ڒ�T���e�[��Q�7�2wp�R֡ړE�l�Up����W������/~�Om����><�i#�m�'�چD�<�+sd����8)��2]�@�4mW�ʲ̰%���[׮�œgqU��B6�DK��4���P1	�F�t�=�∭RJ�
�-)N�U y[_\�dy��z_ $�Aʊ�8e��s7�������s\0N�_���g;�m �~M��>��j�o�v�$�4��o��i����6�9�
�2K��R��vM��T��Sq�|}!a�R��R�%@彮���m=��?�]ܷ�VdJ�ʥ�Di�B�cxY���^�tkH�����b�un^�BO( ��^���G�]{���g8=߅�������p�6�3a���F<��X8������l��[j�W$Mё�>��p�9d��6�!�?����Ek1�E� ߔqO����r0�X�C�&��q	n��e�j�l��U	�\W��n5�� �|��saQ\J�z��k[]{��-9���~/�am�,6��q���WV%����@H="U�>�R���]Nm�qU����rU=n���ŝ2O�Bb��%�Xl�u:����Y!�ў��,���t �͐1���ZY��m�g���D�����"��w�(#$��g\�����)	��]t"��4	s-�����t����٧�?��m�5���E���hC�;)���kH���\B8K�@�4p��'�jko�������s���{�w��s��b��33��vGi��.e��3m�njˬQG o��H�6e�m<\�����&0���Y����D��*�F����++R�H5Tl��7����E��	n��#=GM��Z�0vS�KP�A�/�����s��kzO���I�����5|S�Ln�r�Ѳk�gyu�2��6��`"�|��k���?>���[o�%�������6�v�:L�Z��C�@c���<��8*���{:r�.F+�Qg0��T&�iu�e�������U�s���iiOX�zAM�����LJ��?�0s�i�t���b"�~�E��N��K,]���\��u�g�"F(�	_/϶�3�𲉿����%����e|me��1�g�pUz���ܙ�RY2Qb�^����)F��*�����Fl�<�C�o({$Z� ^6Hc>CET͘�b���'��{��O��$Wj�,��s#���������;��&�1����4�L§G���������M�+�3[7a�M7�ӵ��Ue��Y��h���e�E��?I߽���L����խ���߆����C�)��7Ğc�����;������ԑ�7�r�uZJ0���b�M�g\�ms'���FX6��q�<	�9�?���,�=�Z.	5�����Y�!q3��u�Ƙc��pKэ���nr����sp?�}#�|1C1I�+2&e��. F��#�77�fe�U�?� �g!r7����/���pC�c˩��a檉;�~�L<"�ۖ����ζ;XpJ+�l��+�Y�<��K�{&.�{g�~X���̭��^�䅧���[t��J��Ld�AS-l����m�CϓP]ƍ�n���tR�Zt���q��x�����w��7g�Z;�|rkV�B7�o;��B�����/TB����	�j��h�>X*&A2AN����O��f�n��$�5O�#�a��w��)j~5ZC��M��'UE/C�V����ڋ������K�_��_y�;�Ah�g�q/<����D��.��,�D�������-Ś���~<����b1�a�&q�����c���I�Eعo\]�eڏqz��8�w����`*o�yY��[�6Cͦ	�i?���i���4���hm���^crx���:��=e�FQ��!�MK|�KS��vݪ��؁�d
|�Ï.,?"�(�c5p\����_��2!��RE/Hf!C�����S��n�?7���M\L_.*�ȹ5�哖I�~7�f�܊^3�4��֛����n�,��n�xސV��}m��ō�X�!����Ӧ�z΄yVRݶV��^��݇���~����l��f��KT��_ZZ��0Z���ӿ2�w���~[��p���"B��.p����lIN3�$_��X��*��YUq"�QCb
��T4��.��/[jc��~�Q[��ɌMjM����5���]�����(����a�,&�E��LJM� ��x�r���{RU�p׆l�sN��_��*��]{f�L?�"��_�b�~���ӗj1=��U9�]�����_�ƽ�o��۷⇏>�G�܈W�B�k���������M��ђ�G��g�4���E�6���^�c�������C�w�s��:9Qз����)c�[G���``u�n�O�u����yr��=?�扟;��$��暭��B���>-�,V�8�a�kw�x����<V0M}!��&Ϳ�����؀���`{w�t�zYQ�(aIl�y6E�,9�.p0�ˇ��-�:"u*aJL�jDC����7�*��E��H&Z p�ē�r�t�Jo�VO�p�S�{��br}0&�A\f�os��˴��̐��D[��@���.�rg���� ��
���?�_���.�w߽��>���k&� f�`6zf&]�n<�u���3�0��ֽ���yf%ӆ&y>�������-��Ĺ٫x��a���;x�ȧ8U�s���V���U��VDK�T-�⋴o��1�2fE�F�f��ݥQ7�pϻ��}I��qZ��A	9��� ��-����<��;R��.�r`���"\��P��MZ� �Ȭ��z����\�<��<������Y�"U�����Κ3�1&���⨲��+h]��3��h�:�K0��ȃe�	+���.6ݴ޳b��]�ְ�+^�Nn�4Nύ��`�D�'T/��UtDt2\)�t�^{�=����8r�".v��B�s����گo1��;���S�eNy��g�����u4����=���&�+�pG��;0��qw�d��%�P�����/Un���@k��$µ;Ȅ���F��Q��9:?��0.Y��#�pC���V�(�RH��à���Q���r�V�XꐸI>"U���IY���dW��	�-hZ���6���~ف?���2Y �x��Z�<�j�V��)�e���w-��Nk=��J���ל����"N�$�<����ԋ&��W,�>��n"�~sh���RBQ3��9� ��t���M���g�JpTjl9��7�O���!�i[KI2^�O&�s����a��$0ge�,��|�x �!��[�'2ŬɆ�쩧M�.ڭy;ÙKW���!�ힽx��O��AMv�Z�A�sH�[yǴ�e˦���gt�����8��1\�H�1K_w>I"1]\z�W?���yM��u�iow���"�6LD;ݒ�r_��"�-{���к#��  ��IDAT)7!��vfА�Q���!����}��W���2kh�t�=��2��H���i�9D[��Z����a� Y�v� -�&����.�{� ���Ŧ�~���x�����0��MQg0�=��0Km]�n���,�iN��wҭ�˾-s+����|�(p[6������_��o����}?��.�}�%.+C�N3�!�+��If�F��̘v���ɾ��Eܺ��
��o�H� ��@�&�K̭�]	�dLN����6�<bGR�%�f'������>�A�J=�yu���g/��X,AVx�iPt0�P�"/�[�0�D�R!Q�:$�:<�Ց��q���0ӘA�xyӽ�(���z9�h(�E��$&����"1-i�s�u�b :��P�6����~����׭�ގ_߹�n�7��M]����<��tH#�
{�����Z�)w��M�ZL��eSb*2t��M��2�49��{�lۆ��<�7|������O�R�H������dݞ�p��1l���r��ѴQ;%#��̛K��wh�����vh$�sO+T7W�p^��-]�lb-���>� �zM ���:�mU|�8u�qteiaN�_����&������t���4})�NTE�8H�IBG���j��I����a�m�`�k�}4��c8a�	�GSo�\R8*!M���|����������Cq��I�����T�̤~�Syx��\�����9�-�߅�it7��]0��;��%%0^��3����zN���4��p��bqza����W	�화�[�}�P�V�!W����U����Z����7/�1OQ��P�y`s!�$�f8�>��p��w�a�	xBDh��d�H�7�
*p��UJ�d�Y�-k���@��qgm�<-N�7I��AY#����X� ��%Zlc�����p=����ߺ������y��%���_{�	���n��!��Y̶�����h��F۸*�g�_H������ �L�$�w�/���9�*b�D߂A0���WG͟У�tߵ�Ti�VSm<��n�څܠ��a9U��0x��Sc��#ݺN>�2���\���9�w�K�v�(���0>����<�`r
���Nu#��]5��rr��7A���C@2��މ���P�0��K��p���P�i��{���?�K���:���iX�fr�аQ5��K���v�����8�/�;��b��B�ҟ������0ސ��e:�1�θX�[�a��ҭ\td�h�|:Ֆ���Ǆ0/k3���60�府<�ć���o�_�ًGnۀ�|l�|`;6�|f�9�PN9�)u桌$`/풎�8j���z�����,���Ïҩ؄�'�z:y�n\�����Ǐ?�C'������!��$�33Ȧ� ���p��\�ܢO�����x+���f	0�ę�H ~�M#��P�J�t%��� ��b]��E��>�O�r�m��0U�CXN���֨�[�~�Y߸ad�	(�Zo��⃋oC=���:��m�Q+��������������ID�C��&��b
Ú"`wC�J���B81��"��T2�0LY��C_f(�:�J� ��2�H<�RӸ��{�
�}u��7��7�G;��;l���b��tQj�֭*�.ʭ�/��H�z� H.���p�ߐٷԺ&]�����6��t'�ز	����������;����Wz�4oޛS�Ɣp�V5��_����M-<���8Y�Q�@]ɉ��Y�\V񬔇g��`�,D����/=#�2C�_��Ǡr;�PAu�?�c1ZŎ�㡸bbp���[6�3H`�
O��d�l��s�b��K��{��%D�3��iC�2op#�T�2��6m��R���&�-����H�s.�t��B����ؤ�<�PT�������.��x{�|���w��'/�Bc��v��n	�75���^=�[�`�̇Q��HF �a�|$����Q�2�8��\D9��^[�0�]Q���%1H������� �CT��0�;�V��B?�ZK7G�g�v�{��M�eؽ5������4Q�� nfrWzV�W�`�.%�Kz$^��>�5PX�8^����v��.��I�`��\��Փ��fbظ�@�XE�zEڽ!"Y�>H�`O����aI.�+�NBK�H�	p�Thp)X\TF�.7�U�E�*؟���al6�$_	�~xC�B�24��'&�E`��ȓw'�u!~	i����@R����`Sݨ�Ze��E������8>Ўؒ��S�X����������g���پ�x�Mh�D�t��e(a��n����U=��~��x��!<�.t%Zt�;hi�v2�p��2׏,�e4�$�L^2�Ab-x!�j0��}�/�T� �R��������}"*(�X��'C
HԬ�������b��%�-�*��E��]�����'��G&���� 	.)��c�V[w��p����Jd��yS�u�2�#��}ސ��gmM{�Q�D�{��<�����D[=S�
g{�|q�8�*���^|gӝ��G���{nǆ���(*(h����7ܙ�`{N�tqf�r�^r\mi�δ��yӇ9�N&q��46>��?pN��,����v���S_᫹fa��g�L�Bo	��ʲ�.S�sC����ӿ�s�����T��	�J'}��䂪1��`8���+v0�8�A�)nm��
[6a���M:k�� �&.���P�11*q�N� �}��6��=������Ĳ�P �w��OFZ���Ԃ<,>��!D�T���dA��7�&J�`��|��T�0O�h�sR��������=o݁�B�����mo��7�Fw��Ӆh�����a��z��}w�~�1<��Vܰz�f 0��VY ��#�,���]jO?�b;g�(�-si�]P�<3F!�eH��iV��s�X7��<�(~m���K����a����x���/��)ni�4D�X��U�Z^xn����}/"��"S��h.�ZeK"5�NOsH��(�)%y�:��Z�Nψy��������@L'w:u�Q�����Tށ,�Cq���]��'DPW&i�T�	 �|��YE��a��7f���_<A9U�<"�ʖ�+1�u� 9�pe���wBI����Q[l)������ ��n����c-L�����}�mA����S�r~me�9}�N�购�aSe��\Yٛ�Ut�u��S��� �z^N���9�:x��n���I|���QF�X��m���,o�	��I%���n�26��3�/����"����j?G>޻k�0j��H�]B��n�/�)����H�7�DЛ@�ļ�(yMT�2��h�H��}�r����S���^�B�#Ѐ���� ��%��R7Nj�d{,􁨐�aUM��˰�@�?�5
�?"
/�U �9���7�ҧ���u��{icV���7�ŭ�I<�r�Y���Q���p�BZm�$�c������8���od5��A�a)��,jG)K�+���p�&�Cڜ��������f��˴f�L~8�$��Y��Ӗ����t[��ɣ��{AD���~���/+4_7w���=���݊�()���B�hD@�JU�dz�=R2�#N�c�o���1�Vxᮐ`\={6��0~���m�eW���1��_)o�����{=����FW�M��w�Q�(du�G{�h�J���<���ރW���O�=��\$&�hϬ�Lw�E�Jf�8��f8|�[�����OKI.�F�M��ʍC���&���t!��|���k���G�
'��h��L�y�,���%>D~KiQ+m��㑔L�܌�V�����ܭ�:HqH췢etV����D�+��q ��m���X��sW,���W!����lO��������2BCQ�H���`\��������l�w�)���hm}&�k��\;ȩIt�t���8~x?���{��n�G;��?��Ǳc������q����i��>��g�kni���Ȥ
scڜYv<����|��YY��v�ƍ7܂۟�?x�9�<�^}�=�����_�R�V�'VO�S{�W�RF��B��.��=΄v��m�~�������˷�-�f4$���8�a2y/!��y�/%+Xz�c��1�Œq_�'и�=�R���X�������;�^���ߞ*n�����7�)��D�`(�ņ�n�V*��_��0�P�۝*����D�2���� �8T3>M! L��xR\�( 9�B�!Ldl	!\~��;g6�����3<��2��U�n�*`��?���9��O�ƫ����߀�7o��;���ĺ�3�\��t��,%�
�P�.�|ft[B�G����4%:������i����|�!tu��''��c;�G�ǉ3g�g���� v=�ogV�|��w:E�]=6z,z=-x;%�[P^�`�1_D��N�glyw`Wq��3���Ħ��� .Ǧ%�Q>�a"�Ok��� 0���/i�SHr���`�
�C,B}��t9�8h?:a*ȯ��T���9���<s�,�m<��NN��� ,~��ݾr�P�pWsš��������.�}v�>���߲���ڶ�ΔZ�ai���F���a���8so<�W>8�]�~�3�g��[�Z-����Y�����X���8��VDc`=r�)�ݸ����y9�N�7���������=��B$N�CA*@о+4����!��b�%�����fL��:������6V$X��gE�������s蟎��0U�[�M�&u��A�wʈՑ:�j$����
��)�$C_"�C(.�dq\��T�t�D:�L��qôa�v�lVZ�Qǂ>���(n��h�n$�y�DJ�3��
�o�Ca�A�����ފ4���W�F�A?u�ޕXb2ވE��>��u�0�$��yU���*Q����}��L9�L^�4ۈ�!��b�^63����5֗�7��$�%�*I�M�N��B�Q�Go����,���ٓ��T��}�H�)䖎���y|x�K���=���Oq�s�+�U�[�;�VKZW�"�0�L��n�Az��	�!��`����EH�v}�DH��(����>��\�a���)��0�$ԍ�����$Q�1O3E2j`h�U�:T��������cj�<2��Կ�:�u9����j?�IO|;s�м�~�z%�Ҁ@ӝ\�g+:@�e�o::���e�-N�OfJ#�m8�jk��FE��>�Q%�m��*�m�]*�gm|6���;�?��(vl܀g�m��m�����dA����d��X��k�t���k'1��$~Yw�ԇ�nn.�Ҡ��eћ�,�zqlӍ7�?�����?�#'���w�c��C���Ϭ�ż��N�N���|��ԗW2�ˏ������!��!kׅ�-'09T���+N�Z��y\�_4ǡ\�P;�k�.my�!o����g8�V@&�sd 0r��b������pI����0�+�	��V-z�<,��,m��R�YB�7me��%#X"����V!�\�a���Po�ك~-�*�^�K��]�^�UF��<cH\.PŮ3������O����
�᙭[��=w��-��nz�\ g��P���l�#yK�&�����V�ne�O�8����)����7c�_����3x��O�o�څ�=�/��ou0��/�A�Zpn�bFѷ��1�Ϳ���a\r���]���Q�J9�~�`�@��0&���a�8�@sp��+l��:3V�Y�-Z����и.T�v�:����u�~���0�� 
��Z�)�bUTy�%Tm�#�S:�f�~��|7���}�-/��	eաp��mi���y�Y�]��;��q��9���>�1^/�}��y�Nt �m��LiA��QX'b�4�����7l4,CѪtX��7u�,HZ�� S����!dI}`(N��D�Ym�M���/��{ѐ�"�15�*6����qxվ^z�tp(�0����1�AvS{�m����<��P�VBc���u[�D2�_�>�8�N�w���1G����*�TƩ]Z����m�r��9���A�H���c�:�S�S��������cF��x1i<�,�$K�(x"��,�x%_�6�=!�c�G��ł��X�i#X�%2�	� hq�B����>����0e)�L��j�U�=�H��5�g�c.͛��JK}�˯��ק���wZ-�5РL��)�[��v~�?��N��������z~��	d3t�ɤ�5BdW��~H�r��6C�H<e4.�1X�a0�W��Q8I/�H��q��сWB��/��oo�|Tj�.a�����[���cL�n
�ǟ޼�����%s�-�M��J�CGI/�K����T���f��(��0bYQ���9���Ɲ�3n`��h?��_�K�-a.U��6�P4&Wg�<O�<U(/�LF=?��3��E��-h�/O|�?���x��Mxz��x�������y��I{��0���5ԓ����R�SY�gvA:GMrs��H��[|_�j��-��Ė{�/�^���l�^�~�\�;�e-L�'b2�_gȽ��p����s����zꕦ|��$+��%����EW�K��Rz��3TTW)l�PA�J�}-������^���>�z�&�,8dz�]��@��fQ���^҂a8�R��4�_�P0y�"��.�k�d&�;0�� !$���j�V�<3�kb��uM���Km�=C*��
��z�-�����<���8s��Ov��u���v�;۶��4#��NvU�r#�*�Z[y�cb���K��#�V�Ϸ��#P�����\�1S��g�ߎ�ށW�}�?��W���S��O��Y��W�%�����[J���Zb��s;
�@~�����
S���!�2��"Y`Ȕ�ۊ��Bm�y�+��Ze�dl��:wG;-�˹K���P��B5�� S�	�wHa%E�e�eGX _*NQɒ��V��E��4�?�!�pB	�[5��\����G���;����[d�{��u%ĩ[j�<�s��9�����k?�;��EX�.�.
Y5��2��t #�êAm�*�g��m�q�}���-�J�MC"+J�BL�=q�������'�O�9�[��@ɵ�)��A(�R�j{;��X���B�A��3u�-e ��h��������o��j�Vc��'�d���u���N��M`�4)$��!P商�d��.Vu�5P��P�1>�q��bq�>%�D".U&*��'n��-4���M�&n�2��"��K�~�:6�xk�E����ıpN��
r�ۋ��|{R���vTX�4p���,[���P�)�:I��JI�w��72�zez���K��ÀH� �ts�t�DV�_K���XA8�2��p����tQy>#�����u���&�kc�d��y��DE��g`�;��	���A��� N�=�n���BΙV�8
�G��WB���y2�[8S���[��>NP�\��l�e���G�����J�B���E��U��'>�ee�%��o+	^#F�R�'�X��Kt,W2�&����[i��b�Kk�:�8H�0�fX�xź�@�>1A��K���2��A��Yw#��1�\j�N���V����<�b���C��(�SY�����TQ�O>9��#l��£w߆��܉�6o����bB}^��B��O97�<E�d���)nҕ��>{���{/�4W��S����o<�����=��[o���+����d�^�<�"\	�"q�|)kG���Ks*���y8/�.D9/�&=��3�.��3�T�W�%'➜�X,�&k=�L�B�f��0�7l�!����8�o���P�"=�	�A �k}��z*�܁��E�g9�ʽ�./�z��Dw�gV.C�I���"1C��2�"�S�=5���Ast�ͨ��lfgz��>�7����z;n]�y ���AܹvV�Y����/���|�q�X{:KEa���~��,a�k/�M��y����Ý`�ݷ��������#�:0��W��Oΰr�(P��YL�=�X��v��؜U��k�-S}|\�OF�q	����oL��P�v��ᤗ�Q��>�y�/]7�(A��f���N���G�7�4��=6��7*V�QҪ���H0��[�H�֏���?r[���B�Z�|:��_����O?�w�[��U��5�ƕ�s������]{��q��%\m�����v�s��%�74�~���B3oWZ/L\���BH�b�k��y��#�@\�D�Y!�D��I���p�@��2����J%�ŗZB�� 6�ǘԢ�r_j��`�6�l��B���d�ɫ�F��`��+vʹ�h%&xA�C��b+,�ճ2�s�`'"xv)�Ζ��¹���L��Ϫ�2�ꌾ;�(Àd\*_M=u�j�*Q��|8F��յ!��4�B��8l��STU�	X�&n�2���[O��<�ZW�LO�u����r��1.��غ�ey��=e����A�
�T�2�%��b�֪��p��$�G��-����T}y�]p���m���5	+W~`lת?H�:����!\��6�-���ɓ��������{n��kV�35�n�Ź������a��8��iO`��i}xղ�Yn���mh>��^ҏ#�'c���LU�Ee �T���j��|�67����S&n����/������B��+6RET\Ҡ�-ƕ|o��1��+�,&b+g+_�*G�i${�Iʔ`HE�� X�"���q0���4�.��~A����3�ڤ�QO��rjn�]���������t��jeȧ�p���3����89�'6mď�x��{n��Ag�40{���m�}
C_��J���2�܃���g0^ ����� ,�b]ч�����M���O���o�	{Ƒ�������H��*�TS��e�3���Z��)�����`X~��v�5����7GP��`�t�.#�ϴA�򁄨T���a�$�z6��R�}J�[4n���B��DlS�C�eډ�����G�H0��JA��*l�(P/'�M<k�H}a��	P�ޔ�?e?+�i�
i�Aa�}Ҿ㖳|y��Y�3Hdj���ճg���_����ģ�o�w�߆gvnÝk�ajrr^	Ѧ�,c�Q$��\:C$�&�ל���b���N�]���5k����E�y�8>��0�)�B�c�I�<sHUVj��-�iG2��!/׃���q,%����vz�C�A�/�@����:Nn����� C��:�<��-��6��W���0��Q���)�݃�S��D~�<p����v3?1sF�i�<����:ד�4<,�~d�!M;�C&����o0�$-Yx>Vr�'m���W��f�>l�a�N�Ҋ�o/]��㬜�\'C�z5�s�	I��e�X�-�W�e����i�:���&t	�))��~�>���"�.��*�$�|��g�z��I/���MlLl�SQ�=nBMq䅀��h�~����0_|�4�p�?G%�1A���s���ǖm��d*���7���D����,Z�4G%��Y�]�`:��dߪ׮���k V�ǟ�y�\�ƽq�$Q�$��!ΏDKW�q�	�5ť�Ԯt� �ד�{��M�̠m�̘�"UX\��I�d�� +6&[!x�(e9�uP���\�~W��A8�l#ˁ�r���*\���t����c�z��9��R�^�Ҟߚ��e��pW0�T�v�S
_X�<O|�]+��c~4�KƇg�}"�o?ɥ�4�XΓ��͍�S�ͼ>ֆ�j�m^�/⏑��wưB��+s�(�n�y�Xk���z�~����k�aݪ5X=3��٫�����r�ZŪ����h�â��LW�4gVF��,�1�p��.İ�_���3j�2�1���ب!�&�W�gB�
�V�au�����y���̊�;�XΑ��>9K��RI��)����J�w-59���`c�p�˖��dVĲ�b���kz(~zxfc���ƀ��D�Ϯ�!�st"���R��x�	ſ��τ���0���Ҝ��s���ʵ��i/h��O?��>=�ۧ����;�������͸e�jd�6D�h�Ձ���e:dڪ/�ڱ!/�a% �V���̖ԓh_�ã���?~�I��ӟ o����p�3�^?Rs�Zs�\��Kr �W`�,<��X���d�B�:1o ��t�nX)������N2E�^C�iy�W79�2L?h׸M�[�¯{:��*�|���
��a(�`�'����e,�ߤ�@؇�L���B�J��Z���(�s��+'܂?0� !���"鬐��U�槅q�%�Q�����s%���
���i��ȗ���o��ލ��|;�7�]����e�ߊ����N�.���\x�)<��
{ѝ�ݷo��wߎ�>>�|hB��(2'��f6PnDCϥc���q���*F��+pp�T�}!S�w��ir@X�h:���Z���c+A�a�:I� �:�A|X���R�ʙpS(J����pJ.�;d�t�+��0�<|
������ޑԸR�`,��\�������{8y�"��+�~"�)Gȳ���w�6� ��L�m�aL(�y|��N��Y�4IG9.e�)
�ǲ:��"�?��Xz��F���x��Rg���t������ʱ��Q�?0� ���QC�@.eTR�fPZ�mL@��ϫ���ס8��P]z�/?�Z��(,j����l,�of�E��Ұ|IY��q���N�/�����g\�C��)$��Sް�K�0�_	J�{��+�&q<>�/.��Me���� .�T	N�6�Ğ�TL�*�g�,�4).������4���R� _�0J<��^:� eE8��f%+��2��n��$��8��u���K�O#_o�@��M���McUh���0?����4����<�-p�|!��0��dK�9JVR}Բ}f�mDlytn�J����<8�MK��Q¥�$E�R�Oz����ӧ�
H!������I�sTLzL�m��{4ѽ�F�!_�2ܭJs����_f|������g���qC��k���a���v�F���Zɑ��1�6k�k:���*o��웴s�e��xiKP�g[�\B��ף��nu0[����G�O�߼w��[��?|�al�p��L!�u�K���:pu���C����@��h�vP{��M��c/����íkWᤢ���)"����V�L���"u��� ��`�^Jzʢ\��C��d�a�R�!���r=�T����ts|8}�"�5��=��߃��7�P�|���mٵC���(M<�45{�n�:�6b����\�X@�����9�*�a�����f��FP��"w�W��!^��В��#/0K�e�өB������;�m7��v܏�~�Ql��VLL�!�v�oio�hF@�$�f0#�
�|�%�-��_��uk���S�DK�ړY����J���VTWr����� pi%[#v~=#HJ��E4�![Ԁ@�kW8M	��=�'�/��Gk�z\�c:4��>=$��Sγ���%Q���6��H��1oM�`��f��y�����yb�X2젼%�����9	�ְ�¨	�6�0���被���;E�c�����ں����z�����xK|�#�:�	q��;��C���H��s��r�Av���X��=�*�ų$�W*K���`s ��n�1�1լJh(��u9��J���J�ʩm.d��g���n��<pT�Y��0�Dz(;6�)'�}`p9�Y�����b�nq�x���`'��\�*@�=-qu������(�B�##�8I/;ьE�J�2P�B`��UA�ϲ&�����>TO}L]yXeM�`�S�H΃�K/����<�d�&;'�ae��3�m�X	l���0��.�_�fT�\I�I�)/ӗw]�-�
.���L��lͰ�R�#N��ס2.��柔�9���cU��c�c��D/�abR�;=�_p�,3���-#Gi\�9<�z�et	���!�Ld�1`|]�q��8��4T'�Pzy�~�S��?�&LV*�}�XŻ��q�UH��^!�tP�$ؔ���_6x%��;�aHɦ�R���N�D�q�kWñ+y�H�(e��ĸit�j>�+�t��3�Tχe�����EO��3����4�ä��ZQ^y;��(�<<ˎD��ӗj\����܍��_��7��v�GO�ĭ7�A��A>��Њ6ʞ>��JA��X�ͻ*=�A��t&��,�]�D;ǆ��q�m2TM�{A��Y�boRz�j��x�-~>�2Oj?E|��ý)H'PKƻ��5M.2.G�SE����*�rA��U0L{l�1�A�[/��N�0K!-�\�jX�����FQlL�R�H9����3^��~;f�)�$	��6ι�D�<?a�3��㐣i	�C��T�v���w���\�Ǒ7���z{?�o�O�{���V��m��x�+��'u��95�(�昺�%Nk�j[xn~Vj�k��
�&>�~x�w� ��|Ț�b�s�
�,����\Y�V} -\�������\� ���y������@4H��v��c`��P0�6H�=y0������&K\J�H�oR0��g9.�w��)K��ؗu�űn�ፆ7Ab|��V���.2�Sb��.fh)�Id�(%�b�0���kn��@i�o�1�LTY�G�D�(#M��Z�L��y�5߫r�F_�Նd�\T%>㘄}���f��~)Y���C(���U��K���f,%r�2�;�ʦ����x�k˻����Uk-� $�{���1�Jc#��I]�~���|{"�yW��qM�0hۑ�ǡ__��]פ}����DPU���S��5������	�{Y�G�{������@�bq��A{KP|{ LJӐ>��Y�JŁ���]���ķ�@�L\Cs�T�� ���9���@�1�Dr�dV7�7��"�h�dYx�b�����#!S����Gr���n��ܒ��FW���.#	9�J�L?��a<j�gR��>P�e�������ƥ�
�e����YY.Z�I\0�+"<����\�1"2�:�T�`g`!�)~{���X��C�%��r���)�?���Őc{�D��2��C]�����nE���i&=�j�~���W�K���e�,�7,$C�
扱LJχ+#���q�\�����-��	\��}o��*�٫����M��m������k�:L䙱�D�b[L[� �^�v���������..�� X�I4����M<��[�ܮ�2?>
�%��YE��D�*T��!8O�8����+n+����eq�Cu�� 0(���@
�Ad��� fY�42�b��X�Xx�` od��/i-�GV����,ǅ෬�d���哦}� w�RB�C���+B��0 %e��
*��qG�M�������#\��+Ȳ6���M��&���YZ����&Zci)���(ra�(��ŧ��oNyۭ"^�o�q��������G�����<��v���<���q�:L�7Z�>�>H_�C���Wf-?33��8p�K�'ۦ�txH����
umW����)����m#�z�32^ ��m�N�!�'Fl΃>��$�5��:�r���.������D�<���k�<�A0o����1�MW�1�7���^	G�R�g����H�E>g�)A��$�B�J�"�.�����*��Ȑ� W���t�S��}N'$6�d(]�Ud:a����+�m�k3o_2馊�>	�%�K���r���G<����WI�6[.��r1��J�jЏ�|�_J����h����=̌b:�)�����u��0Q�r��)��!Or
��n�n�s4�j��0X���`p�6R�;Fy��C`����==������*)m#������cuE�1p��}�8�Ck�(��WM����!㚔�d����؏�Ɋ��]�δ~̾Π�ё��d\��i�
��P�;�e�ulI��p9ђj��N�_}�e��h��w��,g�fD\��S�G�<��W°6���T���N�q��y��W�1282��|�>�J���=С;Xx�S�?�^�o8�����ᶡ�c�@�8�v
���.�l(��1!����]��ȑ���C�g��H�f��WL\�7b��%���:������&���1��n��#�e�g)d�ʘ�Ą����妚0(��$	Z�rh���?d��L���B!��a����@UU�z��M��C�����c���`Ba�?E�*	Z�LX/���𺷖0��Z�W�Px�6F�<�����`���i��|G}�����[�|��-��'�c۶`�̌>�t�;�>��|ݱ� ƞ�����p웳8q�[�;3�<�Ww�r�S�������~�?>?�g0��ὣ���'�ҍL�QC�c�{�	�(_�&WV���uQ�N��TP�Y��R����Vк����Ԃ��7 ၣ���� �h�b����:[	�	Z�bF����tݍ�P�o�	�t�QB�����j��I�v3��IdV��u>>/Ff���dv@h�TƜ��G+�	#��CŖV2�;E��I|[��_��O��1�����?�~����ޛvYvb�����Fh� �6b#@ � IQ�%J#ڒF�3����3g��_}��O�����y���gt|,�3�%�"Ep� �5�F��Kc_������%2#"#�o��W�@׽���Œ�9��e��yN)�򚜱�5Ӵ�/\���|�JN"�u�G3���zN�|6�G]ШH�v�	C���6�!� ��uy�鉌B2���v`S~r�,��yF�-Ђ���@������w���̯�D�ګH6�$g9n��	���f��B�.�'ZT�R���ͱ,�2�D��n��g�rs*M�j=]�1����H��.���w��8G�[�:�]�c�n�18�c��<��󱱕,��¹AO�f�LJ�Hc�>����$F.#jʏ���� (l*�G�J����hs(/��Gi�%�������hN�6��csL[���EV����^�<E�G0�mi3/[dV�>�DpAܬ
�C:�����]ٌC+9���w��TO����h���K"8��҂��RސoL������9�\FؼЗ~�p�ܲƶ�7%m4�|���A#yD��^���3)��&�ߦr�,E�g��=�a1��2��^L�Ͻ��
��k�f�� 0�R|/�8/����ҷ�>�(���������r�<���$�YxK1�es��W�i�FQ2M�F�A�hm4(w9�έ{�D޻{����+2�Q����:-�p�5���2lB��S�X����eDC�i��Nj`�Qr��Q���S'�8R����ӈAFPd2 ��s����g�U�� q�,��?/����6�t��7��s�"_ɩ8��B�N��߶�	�@¦�ҫi���)Ly��#��]m8��`E���4q��qO��(�mm�����M�wq�?/v��cO¿}�a�̑K��~���w���u����wb�I`�ݿQ#4�P�ak��q�<y�LlpeoPꅞ���ʲȨY;Ӿ��VJ�(��]�6%l.�:�CYt�S�k�;1�KO��=9�1-2����^y�c⚳�ĺ��K�"���/T���n!���UX�
��4g��T-�,�#��d��&D,a"����N��e������j���a��ax 4��&�d�ܘ��3"��͇m�om�N�h�?υ���c��rJ�Z���0�8 Ϸ[�?~�~��<������?_����c��y������4\$�MG��k���_��oÖ�h��B3֍�{�{	[,�3}"�@��˛����I��,p��{� �����zIN�)��Y͆ ��<�ds������= �,
���(=ÄR��c]\�CW�YN�f�
N6Ǧ�L,I3?�a���H�-)"�I����&;������^)s9���/��G����N@4�Pc�3�B�Ka�&M4h�?�����֬�U��!Շ���і��e��ɷD�EJG+�M��
N�{�h�C���r�а|Ÿ�iC@����ª��b{����a)i��9���˹�F�@6���Ѥ��;&K��
*L%��%�'A5�I���*�rb}3�V���V�O%�,`���/ϡ�T�l�����foH�h<V�0�d�hl��!6sB����Et���J�HI�����'\u�vJ1+��߀�&�Ad���3,�[)���H�%","�:��b�����`��k�x5�Eό���I�Mם��r3���7񴤅�mT���G�C'�أ�3ҵ��h$��bl�3�D�D^��Y�{<B���M5[+��q"�FVb@�'��!(3�ZɀQS0~=G��" u�\;=��u���%��!ɩ���K�uu@걚��n@Mט	����𘱺}$hV�d�]6�{0�xÖORh�!$�6d�gQ.�"2�"^SQ0ً��wm6|D/ �]�쎰Fwh�.|ܬy#H�O7�+������;�����\�7?���\���O��?~���hl��<��M�zJo��������>�(�mplF&�'���5��؁w?����e��NuV�{0�x5�Z��m�1xyH���V�`�c�G����>������a�a����zD�
���9P����jn�Ei����)kB��J�|`gzcHE�)Ku5����n0������c����n�h	���sC�o��f�YE���]�b�]�����O�~��_���|����k����f��c�����8-��r�M�ޛ��Ǟ:��7�	G�<	��ۂ����Y�G�F��CT�>����}�l?*\X��E6VQ�SwEP<K �yt��N�lgـ�n -p���W���L����Ѐ�j�)]��q��@q�aZ�#�D�)U�l̴T[l���'�"
[X������[�-��Jk�z6�6'�7�_s�wkN{#��)��_ݚu%,�%3��0b�Rg� �5�� %�S[VɠG�g�Fɲf���e�sMy�(2�N�֊}	��@���n�<p�+/򂛉^F�m�:�և��S����xg+N;~�R����\3�����h�(GY v��y�Sg�Oā֋:��ʩ�兺���FÇ��3O�B셤�8�ƒS9Df���Ee���N
�zZ�g&|����6d���^{�5��$tW��:��^U�ۇP��d��<��y�)��x�h���njЮ�H L߉����&�Y�ƺ@`�m"�AGq��� R]�z/m��L`�u���K�I4�q��n�Mh�Q8-l�a�m�,�ϗ�ۤ1�����Ӿ)�I;��t���9�H'q٩�'�OI#�fQ�4k�j��"Ә7�6߳@�Ͳ�w���ҧ�aM�	ݶv�����0�lm,:SzCh�z@���)� C6u�o)�(��'|W�d���=��m6X����?q���6v���0��	؂�{�s�8\��_����O�
���:��G>�yO�[�w�Z�o~���G������
Y��u<$={0�k�xK�T���@tL�W�pvm�GU$�9�@����8/����j�(�������9��dMfT���0���Z[��� 'y3�?)���%�Q�4�e=$������	��)�)B_�pa�20S0'd���%F_�'���fA�	�C<�B@�b��F����m�p��tj���l�o_|�u�>����g�\�����7]�]x���L �}��?������f�������t
���6�t��� *�T`�Y��[��Җ�	���0z�Ao'$+�/ܓ�����Y����׭�ف��N*h(|�z-8�As?\;ŏ�<�2��y�'�z�A��
�D�5`H�1�X�J�s�r~J\����
a�����-�$�w�D���.&�Nyz�|��:|�O�;�/�y�?���)N0>��#"��M�L����&��<'�f+��@A�AS��r�d�5TF�4MJ&9mѲ<N�i�m`H��ƍT-�L���������(���F[ä>����{��-�t��m����N���cVhA1�kl�}Ft�(��:$������r�@��J��';��1#B2A�N#����|��_���
���J�(-�OZ���#�(�4�����ŵ=a���q�����2�<R�8b�0�"N�h�=���wE���d�bE�5j����4#��ޤ��`� �:&rv^S&0��8��ٛ�6PĘ1��J���`]�$�쁃�R�s�Џ4<��T�])Y� ���Jr�J�`���1�Q�&��PF�?7`&-��ia��)���7���ϼ�2�5�>\? ��:�ǭ&�&�Dv�c�k�U*W������	sr� b�_v̺�+m]I�+P�Ɗ�J�Ƴr�! ����Ԉ���e�O� �SF}�F�8S�f�i_�],��yX�sv{�s��XZ�	��_)#J������������d�6��2�³�^����M���^�E�t�9C�>n�= �ك�G�"^M���7
Wc8��|����-����h�1�8c��'^��|�i���u���7�����r�ep���N�لx�W�?�<p�xˌ���FWv�/�&����mcۤqG�d�Z'W[9����|5����ڛ��$�F�4�.���d�g�>�����ק�Ҁ_�Bt1a=3X6:A�����ɀ#(����VL�g:b�fāw,�g�2�����d ���J��jч$�S¤b���`d!��7�����˅��
�tO����^9�7������q�ݱ���eG�ٶN�uJ�F�\_���z�e���
.9� \v�a���!���������ih�G0Z�����]��14I��:$i)��u~L�gh{���7�}��,���6�^.����O�=6~��g�ib����'J��g��C�3 ��i�e@2F�2�N��l ���w��F�&~�
Mȧ̟)Qq�P:�s5-Ȓ���nR�ӚF����p�{����bT��)tW��k��f��`�����G�~~�λ�ȥ��;q���S��+���>�y�q8�֛�ƩN�:���wY��@{7�
����L��na����A���2�jI�A�u��1���F����w6�� P��oI��O[F/P��v&g�3ϡi���D3EK����F����R����Z6d<��Ƌ��SRJ��oһ���)\���7��u�ᚤ�u�m�&hw�rw;�4�l����l��C7}�E&{�]�SÀ|#y���}�����?����yF�O��4,)��eoW:;�[_�i�y�u�r���ʫT�^dJ�O�c�h���	�!&���OyY=<���Ǹ�������8)�_�� ����i����y?꫞'��/A����F&8��~j��s	��R�:(��M�/J�IO��9
Ƀ�k��WT��OS�$�#����\/�t����u(�TqP<`��!�p����>��/��>y���ѥ���7ބ�_|���G��c�����������[�B��3v�)706Ȋ�;w�dԃ�Ϳ]{�Yzn�*A���f�{�o
�-��)�ǐH@%��75Z浴�MI���S����G����s�`��`a��Qd˞<gS�S�����k:�'�z���Z
}�2N���:���B�q����FG
㽲z��Ct}���e?�5����y ���(����[�Ǭ�sn0�&xŰ&x������/�&8N���L߸C`��d/<y���#p����.�؀�_N��&���;�X�`��z��s�X���-�,�>�A�O-��(8���p�z�����$�����6�������rJ����A�d��ɹ3P:P�'�-`I�5�>�������=�]k�f��=p��vl�V�+�P��� 1[�5ba2Ai*��* �6MX�qB8a�j�z���Ǳ�\�(�ǔ;��!��ov�����et���ND������ҷ����ϸ����~��w �?w}@���ڃ��Jq�M����4���d��T5��E�A����Z4 ��O��mG7[��b�!����<L�%K�UQ|J()���Fv�t����R}zO3&��yL:�A*A��>.Σ@N�P��mv+��pZ�+~Kڬ�t���ozwJ��h���&�q�G�_��o�=��#G �e܄C������7^�������x���SO�/�	o9�㵎���V��#?�B����6S-�1L6  t�fښ� 6m��;s��'�\M_�|�yk��T֠O��*UW�W�����2��ˣ��"��?�`��1�к��H��;�}any��Plq//^Q� ����D�P�4V	S���}
�8�ᧆ�t�(��d�8�����H:����P�����S˳����`���t,d	C�q˔yD���MD���E���
R>9o^���Q*zAn[	I�9�d)?�-���0��Γ���b��I�2�l���3���Hw*��y�8A^��u���<xM���i
׭�d���x3��'g��w|
����M��С�j�C_��/9�^���O�
'^x~��;?;����g��wOé.�f}=� ��^sF7΅|c��6o�Z2ҳe!���gSM�Y�q��E�/��S��&�&�٩��l�аű~,���`�8tC��,	���y��C��>y��17Hat�̆�ȴ�>t�S�;9�|���b툕"�.eE�5�hc�=�3D�Z(W��mb���fs܃i����5�;�	�G�Sp<���k�&�ux��^8�F(���9oF�:��M���Qܓ�H�U=F�SĐ��=���$(P��HW�PU��v����|m�!ed�⁣�0���T�I�:���v�u:��rAfA�	k���ֹ+T���;˄�TlY&S�����ڊ\_6z<�Ż���_��ć��T��^�2�FK�D^9B�fJ���,*}�QU>�|\�s��xn��v���_��8�Pӹ�-aA�Yu�}���##랍M̭��)<�4��	Ĳ����С����df
Ub]&��w��Hd������.��e/en.�Xk9P��
�P�\�ۊ�1�x�6p��~MT�H}��!	Yr����@�n��'�oTX�M�Hc�cČ+���[n���ƹ"l7ᮋ·��?����U`�&�xZ�|�NJ�:>�~!|��;�7��~�=x�ċ��?�<�ƻp���f�+il��0=�ү�@�&��0Q�s�7�&�<��*9��iN0'H��s�&�P���@y�dP�U`&T��[LH؀M�z�DQ[��U��_��Q��]LdQ��P�ڙ{���
����n�xWO�����EeA|�0n�`��P1I3Hy�'��ƿ�g�41���ʅ-���[-�$�K�E{ю����iq��ޗͳF��v�I'�S�æt�s&�،���6�M���A,٨E�-]��Hᙆ�U��7��EVKGYb��9���ư�?3�[���bW��7�F���Ѵ��T���琄�@��
�r���*'�+`)j#�8ǝ���{�h��H�i[��y�-�'w��������3�b�����_�m7^q�x�u�'��/����ѣ��ǎ��O�'ϴ!��.�QXSZ7A��^!g4�r}�Ը���1��<n�K�������dL�fi�	�f���B�Q���^�+�] ����ri�M�>Ho��46��gh�\H�d.�5yH>v�(J��<	ɖ��Y�d�=��2�FK(8.�QHFoIyޥK�C��|���w�l�<��/�m��t��l$��Ϯ�5o]�8O�q��{�G<��=��
�&~��,��"����)�z��Isv��yS�T�4���`�!��jjG�#��5�-�⟑��EhM�IzcCf;a�P�y\
�p�J����bx�i�t�ʐ�@ʒ��T������j�4!B~&> p��4�ixm8�pd�h|@���f�c�'eq��{5���6o������vV���[�=Se}��!����m>B��X�G������F�Pn���̩�E-l�P!�#-\�pU ̓J2eʨ�"LS�T2LiÁ�쓁Lc�)�=���|2+�F��@��y쵖[]0�|��O��'
�&�{����,�3�s�ҞǸ��1U<��)��^6�&�T�|&߯�0O�w�V�`{���|�+�L�d!��Dt��ѽu(�{�s���1|��k�K7_�m~�{���C��c'�w߁Fk0q��z�I>U�&�9�;_k�*6(5���ăh�blb��'�e���2/�W�a$�N�4BBF��J�H��NK�x��u���t h�+�jQ��1Gy%�������`� _�*GA��5ݠ�ql[N��9գ�>FY�q� ��K�O�^*r���LW� �r�������O�p��7+.C�������i�L�S�`E:���F	�W���A�恲�1���ܰ���T<Cp�NQ���V-�Qe����TG��0DZA���sms��~�Q�N`𔪁>�I��6aӅ�x1���N[���O�~y���1Q,�e�������$�lmn�'.�����p��-m�I�/PAi㷭�^�C�qW��/<��W�?��x��w��?��c�ȫ��+��85���Fm��Q&�ƙ����x5�_���߀�<����bC.|"�Է
�΃��H�9���ڠ�既�}WPQ���{�H8#҅��d˄���=�6���1^E8��N9�t�d =�a(���P=a�Ls�P	Sҡ,�r����y�%�cf�eN�gs�L���U-*)SaeTpC�Ә�H�vJ9�]���zH�����49�������7ΰ�C�Z�1������Κ��2�̇(��A[�}L�t�t(��=f����&�w/�8�J��>�c�G@M�y��g�:Fz�!;��!�Y�y6?��s}�@�8���}�Aڜ1�T��K �5�4!���P��$Tk����L�}�z *�ѽO�oy���DF�x;uٕ����BJ�lX] ��QA$����f����&�n���;�ºF��ʔ)�V��b�Gl?�kS��A*��	,���U���hh��|Hڒj�T���9,�Xˁm-ۈ� �G����]@Aj�b�tM�D�
q).*q8�&�m�zT.���ߣ�����z�[�eFrPK��P��H6�H4���!��6�,H��{2y`ÐP��'�m�"�֩-����p�UW�Sh-!ʉ7�\1_D�Q�d�=�·/�r�}�M�ƩS�c���=
?y��x�}8լu٨Sʺ���{㰑�{��Nikڸ9��S�)G�J�I	j����i���uS_!̠�:��4s��cb&���Q� ��ٴRj�7M&j�拶�2��(�&� �mg�M޽6.
4
j`�@z_(�]���Ӥ�ca��0�e�Y�!��&�F6�z��W �k |�h1�3i!̖ϔ���D�J�H�&U�0
���9m��S�����Bo$�j�s0T2?%~-�Z�<�I�2�<��
�q/�����SQ��:T�{���Hy3��¤=\p@FN�f&���*��ռ�q^`������J��~Q,�����@�R�ţ|�t��^�����a�+0�s�e�ڭ��ѹ�)`;X�[�Wo"z��B�E_$H~3��5x:�a��#�M����N�/������Fg6᫷����+��O)[�6m��ώ-�pcW���{/�?����7ނ?~�{�Ix���f�㬭C�)<k#�>~�%306�8�-��K�(�1�=�rŁ�ZțwzK_�0_e�T5_�"OB�U �L�d�:�,ܕ�0�ݎ�Z)��,�zHO	�@c�n�=�.�^��M�#���~��`�����M5��f�.�΢'DM������Ho��>�8S��4�GJj�>�iH�L������%�| W�$d��Q�1�D�!��$_eE�2��nN�d*�CM�������|e#M�Y����!��B��g��N�<	N{?L}�E��e<r��J�(�'�}&Bˠ����T����A�C��J��&��q�{ku�����
mԶ���sW�,�H��N����E�w7(���E��F�.P-UĞ�
Ȱ).���&�@�,�'�ߥ�
9��2��Z+j���F�'�*�)�,��io��G?�^K�.;�XL��#�\�yI���=�^?'r�R;K�!����R`��Iޏ�=J�����Eب�-�Oh5�j����g��m ��GNt�M��ʂЂ��9X��d'5q���w:_1�����8.����q���i�����o˅~���Q ����:u�C����p���puJ�y�-l<h�h�1��&�w��8t���6��O�
/����i���£��������c�UVc߶���x#�D�b�4(��Q)2�p�^i�A�D62�[S�P#',3���L�/(|&�Ӹ��� 5vVӸ8��&��%e:�9�jhݼ��r���ɲSP�kD��&~O�˕RI){vS���� �ђT^�i��՚2�0 zʭ���Nha?���aw��+u�?
��H���������'�Mx*�hZ��mZ���a�F���J~0�̙2�U�mG)ھ��,-�a-Ɂ	{�>�s�o�~a�%��L��W+c�8�����ٸ������WT93�R3��h��#穗�E~�.��mR}�^"3�|�^�r�,ǹ�Z�4�jʡ����uи�_���T��)b.r�f�/���n��b�ĕ_�?��g��/�wz~��������Z��4an��sFn������#�9�<��(�X6r��6��E�����j�;7xV5~0�]2�$jW�8ߜL��Qz�;�,�D��<��	�a�kWay4A�o���DA��G-O�oj�;�R���3�Uu~P<�f?�X��	K��r6�x)�[���p���7�}�dih���J���Z��+���}�R.�J>oX�YL;"e&y��{0O��QF����̗fad�HŨg?R�����e�����7=�%��}m ��:���q�Ua��D��ζ�ꠧ��pL�z�Nh-�i������;��8��,��^��l�!U1�~�T!��,���{ix5ip�V�E#�\Q�̧J��Mэ3�%v�E��	���WƇ!MV�Mb��B�$��ʲID�c�-NE��G�a� ���-�����1LTh+����7SX�yX�V5+.CF�p�N:[4�YQ!���жq
l3����(�y�Z��@�գ:�XЖ
���J�{3e�~�p 4 <i*`��Bx$xc�j�J��\;��h� حhЖN������T:�N`��s�G/��r%��W��?s���;�v�|�=x�#��	����}iFAlwf$���h��L�݄EM�5�$��­�~��T1�����0B�и���iq�7����DV�K]��Sc��V��k@=p�S�;��F�ي>�I&�Ʌec���L��{jC�,���dW�YԘ�,�Z���a*F	?�^ e4��d[�ւ|�z)�k�Y�<$eg�T��zk�<}j�
��/���E��o�!qlabL�J�V �l�y���9M���~=$��^�uU|�ϡ�)��-�7�(o�[�Z�!�f����}Q=xV��~/1������+,�y��A��)��C8Ocz��B��e��ܲ����C뗣�Z︲�Fk�>q�� ��U�L-~L9��M]g���1�kC� ��	��5��7�go���o�Ϟ<
�}�(��9x��>�Ю;O(���3��x͆+ۘw�kdO���%�7K�O&X���:h�LՍ76J�α%�5��Lŉ�O�����)�Ѹ��c;�p�X^��Z ��� ���T\�)g�Q�Ƒ~�,�Xض�3�N�W�B�Ѹ� �өцeznM�Yơ�*��4�	/�b�6>l�D�O1�����y�MJ��ܺ��0�E?ܿI�r��Vz˝��|h�X@�&�A���r{1���TNB�'U+�#��Q�#ڨ��|E�y*��7#ޓ�:���嶙�ڠ�s�`��'Z}C|6�%��[
�ݖQ4�����O�f��� �1W�KI1�g�T��օĭ� �g~��)j	�@�,�|�M�۠�N.�}s������W�]�b���e�H�*�n/� �ax\Z�"���K�-Q�!���S��� -u���^s�yC��`�c���Y`�.3@�&��T��4���^��1���Ѥ�X�M92��m�%�".XF2jȽ힓H.���L3�g�N�:�m8H鴲�U7�m�H����Mo�q��k��]��_�g^{>~�{�q�ѓ����::��{�:Z�e'�?cg�ն��0�@�`��+WB��>��' 8vh�c;� L� ���hu��������*B=�,M%l@iEv{��;�N.̕��_�5�r%H�m������vΰ�h@��b�2Y��L�
��+�ԩ֫E��_K[5,����٧��}Ӗ�L�!�B��.%�!�Wu�8���p6�)(B��#�b�|s��K
#r�l�i�"/��:�4���d�Va^NWn��4���H<�o/}����,Ǘ��"C�Y��s>Y��E}Ӓxa�u��D���g��MU&�E0�|�>zQ�Յ$�:q���xw����5���L�gN��n�84[1g����zD�Z�?d�I����7�7�����~����އ'^|����ۿz���.l��8�+(M���t��xM��CQ����%zh���8��}�6�2��٨�(LN>Հ]����i�d�~SD�")��1�
�y&8S �iҾ���X��Ac��?�5=�س�ś���Ȉ>m\+'�YGR0��Pܩ,��L�J�I�㓮��`� �+��%�/�2��_"�/H=��V�yL��7ܾQ��c��p�om���9��a�d��4���s""�h�H���@�f�e��e�6L�'��^}$�����G� �|� ��2��Y�8�%,[��4��y�`Z�w˚R�ci�CT|+��V=��P
V�Vb��A�{��M0j�P�M٧��,�`�6z�h��/�\!.�#�v��DܴM�B����a�kC�<��{�	TI`h@�Tf�@�q��D��%�����v���{�b�z*���!;Y�D����r���F�`��x��)
#}&\A�g�oA������Ã[��Af�#�O��
|���}�^ ���n!Q�|ԍb�\�M�!�jf�FþN@� |dc>{�ep�՗��u���'����/���_�7&[����[���<��N���k�[��.	�lX`�/!\q�7�S��U�G�;�gh����sZfo�ц�&m�����Z����Iˠ�5��Km�$=7�w
f	���'�LR���B�!<ʈ0��Q�3�%>R&���bb5
~�,�Gۍ��4�4��7l(~P	��iXɳ/lV�eY�,k�6�X6���'�q+��=W}���p#H�6{i�|R{������Lm��~S�N]w�}�xxA����9�S�ԌU�F�ث�~�Hj��|7}��Mx%�4���I�D�*�C��f�!�P޷Q��4:b����NiؚL���~��p�E���"�;��}�Nz�I�i�'�
^F�|7��5�χk.� �z��������_���~�=8�6��h�w�W���D!Nj��o��#����O��6����\�j�ϩ:�!�V`Q�rdH�6=�Qe�����C���-a_@�u�u	�9��;�U����7�P��-A�I5�Rʘ�
R`�l�#]���d�BC�E�`����kyg���	����K���&��6��C�d����z0���wڃA^�v,ҫ�E-_C"���N4	g�Y�e��G�H�(i{0%��K�h�8��2mD���;+��cY f/S��s�s�ˀ#���q��u�ʃW$�s�w5�,���7YF�3��<��L��,"�j�(�TY�Rp�'"$���eE�U��7G+9�*s�e���������26�W�m�,9�Q Ҕ��ջ5���AZ#1L���x��6ܨ�
(f��V�8^T��Ն�6�^��r�e��J��I����Z���8�R��S�I`�*E[�ڋ�E�k3❍y ؄� o��R:�.�Hc�ʹo=C����.T۾(i��%Yw0:B�<œ��aS 0:��d�c�ET�ɐ7�C��[��)��5@��f������u���}?���t�|��`�����t2� }#��F��l,�G_k�6�_~�a��/���g�矃�}����'��;�i��060� ���[����#W�6�o����`�����%]k%?��"��3�2o���cHYm��qYmdLA��^d�􀴿�͒CȺ4fH޽b]l�m	�I�O�t�mۂ��4/�9�f�1o^�"�`J����������>�2>��l %���M#Z��'�0��	K8(��a�����Q�Z�o��P�<��G��M�V�6OXm��qQ��H�#O�1��ˬ//����E]#�2�
)�I<���1|lPB�O'�~T$6+Ӕ 7�����d�%Ս��ɞ��98K�
���)�h���4��D�:~_۫GNp�~K���+��U5�HE�D��a5�O�^!r���$-�A�"-�^d�S&��hc�m���ݿ��o�No�čͅK|<����(���jHTs�~���L: �ՁNk���k���5��~�-�ᣏ÷9
?�5x�áu9����-�[���a�E4��c*4.q��/�OހR[ ��o����O���U3����G��%�x��F~��w.�ު��=�/$� ��2��H�P�h�hµ�=�5r=-�9�m�f9�ԟ��܋��%��m! 2}-s"j�����֜�ΜWMC	Sp��@��9.k��*.hܖy�H��q��6���8��Y���X!%N{0r/(�+b���,�7MX�u�c�*b��G���Ji�J�P��-cg$��$(3�����hM@���ɐ�%I���������/����C)�Mj���ՀC��`Q�gmY��%	��Bʷ�aK��` 4:��eUS~5�w��A��E���6�q6 �1�0�Ӽ�	!D�b��a�y��Y���(T��W�>-���hQ3,q'���iX���\ΧQȳ� c\��BViC BS�T�`Ҙ'�sN�'�D�s�ʪ�4����e�0;����ҹ�`�M��5}
ʂM���,��ʒyj�1��,��\��p��SDcbS7�3=��G�%"�6F~���Vc�'���/�;�������;n��d0iba[aG�i�H�2͏�\�I��-�l4䊴̻&6]w������>ӵp�G�_�� ;���#O��_x�~�Mx�5pf�6����qFM��.ODoҶ�51��5���ݤ9-�*c������S�\ч9S�(#�L�4˒֥������S���K�"��e,��N�~�#�SyE�^Q����Ae�J��ZX�-�'��Iד���5�E3�0��z��ϱ�p�k[�}̢���~3�19�T��[�HL��#� ���I�H2O��[ܰRD��/��y[�+\d�
{��]j�>�Q<ǀ��f<2�Q	Ι&��<���՚b�R}C�(��mpCNEsY������E�e$�`�1Z��1�3�h�q�N��.޿��C���o�������T�D�������]VM̯E��G�u<���,�&��{�p�6H�[g���|���G_�^<������������N���g:|7�6x���|b�ߛe�Q0���AM0䘸kX�O9Q�<��|�MG�Ƙ�3#�c�� ���64zz�S�ߚ�0ÜH�TO#)�2H]��*`��1��v���`у	�;G�p 4��1l���Eut1ۗ.�.J����ÓƩՙ>��#�-�����������^/��`L�� jK��+�=Ld>�e}�}l�<��|B��1����XN�?*��U����_�D����=�: NBN��OZ�rޘ�[� �G��?W��,�Z�ꈚ�ӿv�B%��:9=�?�/$:���G��5!�V�.)�Lz
��["�tZ�}�K���B>.�?�iF�d!ʈ3]@�O�>��tIq�$
Ɖ�)��O>������jdSmPY���¬${�5m��m�	�e��6�����6]�Bɴ�E�`�m��2�ї��\���m�Շ4�"�i��̸���7+e��7�M�Ϭ��ԅ>���M&�<�n��m'�^rt�������˯��������h=r$>�Zj�����d�뷅W͸!��5�޶�*�6l��v�ƅ��[o�/�x����Չ����=?}�{��������B�K|��h�Z���z#���	�h�Z�t���
�aFZ�D ��l �=	y��aJ���q�vNJZ\ϫz�j-z*]e"��E&����~��"nV�ӗ2�`��D8+a�d &c�l'�@	��*ad����a�B�8�0�Cb�t�ZX6�&��橑SQA�e�*�U�����a2�!m�}�+,�G��X��lk�'�k�J.�P���S+�c���a��)�OF#_�CI�W[�q��<���/ߧ_�:���4��h���5�a��b�0�T�"y2��.Bg*��ρ6"�H0(-Pj�r���>M̬�t�3[-l:��Ǟ��N������x\�~��F�.���.���K�"�<��e�g�T>}�ӣ��ޘ`���t��?;%�K���t)��� /����3��N�y����ק&�j��N�1#�}0�6�Qƿ�}.W||	�9B���R�B��&�zLF
��`��\�2z���耓
�� �e'�5e�2��}�¢�����mL�W3,�.	��VŽ貈�ԡ�
ڸ\�/�ʟr�o[�HA�4�i�7u�5H�eXI�lQrW�k�}�?Ґ!�dv��`	߫��P��f���6��$E��I{06�5���V!ufu葿"��ypĹ�g���{0�u�_	��rt.Z��^K����cA?_p�6=�L�lP�ɬ�=�G�������:��(x�FB��{K��Cǟ��/x�_������K�Z9���0��4�����'X1�A�ɲi_�7<Nb����#A����w�0-˒qL�97	ȱy�ES��CA'HĐ5��K�C1�I���u�*a�9�) 򊕽����COM���pqZ$�%
�h ��4�T�c4�cd&�^�_h��L�F⒐ �<�����X��� �-�r�?�`h�%$�-��w��Fc���g�{���|��O~�y���{w�7_{5���#�:g~!���]O2~ζ�͊�[HK��¼X�)2/�E/�+}��2[7#���A��S�������ͷ������<
��kx�����9��7�xc�3]Vc��9�w�[���`Пi�!�&߹�/E
-�����hD��MM$�Fvv�s�:� 5A@���f��O�lM�	c%6�E��/U��`���� Ҝ�{��{Cџ��������x]��A*6��m	�I$�1��S���ia��e�j:S�
���F�Ѓ����'��Z���~*��V3ŧ�P�{ju.NQ�Uf�p#K/���GO;d�Q>+���}FX1<� �V�-�@�l1�\^�EW��s0,�*"�d�(�r����!>C��E��|5�Gw�l�m�8�,�Gb�S�v��S�U\֎�zėz�p�F��ٶpf<�o?s~t��~����w�_��v�쒏����z�Gn��&��G�Xö-�'�Qch��6}���MvkӇ]0�-�n>r)�ɗ�g^}���c�'�Ó'߄���N�iM�w����pڲ��$zl��F�c�����m�ڬ������ �(�~��ʂ)�H�H�V
�o}a�(3,�2�j|u6�0������/���1{�܁��� TԶy�i+C��Y�օ�"��U�P
~���G�8��U��jYyTNi���b,�#�:M�	�=�G�d^��B���R٩YLÆW��d:HvE��� �>�C��./2+u����_q~y7AVKEk���w�K>W���:�$�[Q�}*�U~�	��@܁7x������a���Q ���A��n��#Ei�w�]���09,js�{�q����v@Q����x!�Uc�)>��zۄ	L1�Q��ޗu��a*߬G���S7�x-�D����ex�.� ਔ��V�T6A�ڨtG�k��R�ɼR�(ܢ�*mA���.8�r�#���21/u����$oiqG���:�M�=��m�bqԍ
���NKO�OYXq��;m�'O�������(�ol��:�a�u��0~��Ϫ�CN�m��N��֠�%jܕo��2��A�m�́ҏ�s�M�l©�'�	�lvQ^8����o|n�����?	���;���/��� n��uwMrl�d0����/m�I;���9H|x�s�`�xw ���gV�i����/<G���G��,�x�����o��A�����3��õuX����L;��#Mp;�N��1W'��>1hX[�1�y�I��O�`�&f����oA'=,-���3�1�qf��OݔA�,�R7�0\���S�3�;�^�
�݀�AcVbSHj\��n�Nb�r���D�|-R�'Ҝ��oUa��bQ�ii�d�Y@R�$���HBڤ���O�"��D��A-�G����F O�$k�'��tE�Q�D���W�����ZvZXf
�d<�'�h�؝�MK�+>Y2 T��L��|��Ms�&����F7���#��-���[��ag'����˔�"aӤ�\�(!M��ï�e�qM�3T��"�r�J!˰�G�
"Ǒ1At����\gRA�NHR~e���sҌ�[Q��g�l�Gq��6���/�O���6�&�앷��������>w����w�_��F8|�!�d�oW�3 x�H^, �G�acpm��3M�}��ۥ5A'q�M��ҵ�h����u���#p���ÿx�-8��������=����l���ڨ�k�D9Î&��C��c#| cW��(%&K|�� �loʧ��g�jb�Xe��������#��7 �Π�Ш	�2���ܾ�K�@O���	�h����0�v��Q,�m��4`�~6��>����^�X���/2C�cFF�{�Y�U�5����W�|�ʔ{0�<4瞮bA���ݸ�����U(%L8����� �i�7ϏB�ȥ�&�75T�c��6�6��E��f�Ur��P�)�����u����t<�bpʲ��s�W}�5��^��D�cU����M��v��ag�-f7�H��v�A�ʊ�	��`3=��V�f�@�vZ�����k#�� �Pu���t��}��ܠdJ�)��ӰZ{Ȱ�v�y񽖧�Y�+�`RI��|Gf.6,d���Πd`e�������\�*�2AY`����̋2V����
:�s�7+[2	)(��2L�InJBj	�Ϭ����"�*+�yA7��ұ)�~j>0{��9h�L��)��<�nC��	rr�	�i���dx׭�Ez���0�OY2Bv��.���1�!����qɮ�!�]���?�F'#����ᵃ#8��|���������^q�q��O�7^z)�`�J���_E��c�l�ƕ�6zZ�;+���6�q��*��m0����`����K/�/�~�S���o�/�~~��3������V�����k��i�y��p��h�~q��C�+q����=�Q������9�d�����
�緩ęS�u%ɍ$���@O,z��6�%�=.U^� _U���M;�t ſ�P`,��Ya����n�ZM`�ê��1�]�L^�;�J�0�'����D��iy�U9dX��D����4_-��0%L�flw�FS�o�#��=>*{t$�-�C�3x��Ǥ��U�PF�/F,�2�ʴ!r�uQ�6~�)�gVDs2����0�ʤ�g�,�C=k������2-�APR7�˱�(�1��f�?k:�Hf:�C7l��4��ǖ^B��G��u/�7AH�/�'�t�d�{�u�k�Z7���ٗྦྷ����>y��\��|�������x[�wsc('ZIx��!�� Y>��Q�r3+�!�{7�Мz��~=����&\p�|����]�\v���^��>�4���p����]w�ˁ1ؑ��i;i�s� �iB;6��+)�Q	@2��� �J�%��
�|��(�%=�&Rf�o
P��'Bo�E�n���޲*`-$�(\�8F��-l|"yss؊MQw�l3Y�U�e�(�qq��C�»S�KXB���ǽ)�D�R/k��r\�2�V~S�$���Ѿ��2��Wi�Њ7i���jh�B��XQ1�N�"㡛��� �T*��*����o)*����x�����/�&:�a��EO�%v����)�C(W'i	?��>��4�9�:���h�<���zR���Vx-�(&�&�uQ����\8v
��\`�~XX��\�JX3��IN+Ccʵ�K�N�qJ��SMX��j��&D���t�\Jqƪ��x��E���c>^d4tPC�%����r�G)GJ!�
���÷��r��H��
#�����uF���'���i�$^gP����n�-
�m+�<Q���@�ǽK��JmH�dE!5�ڤ�!�M_�!
�~N�yV�L�^JM�QHe��R�<�w6CV��RCͼ�	/xZ/���1��/nN x�p�gFc8�i��s�����7�= w\w��z������K/�Ck�7/�RE��ВS�&�(��Ekv��6�``�gW�������p�՗�G.�?������/�=
��*<}�$��SM���QX$���\�wWߑ	:�K�&n������uO]�~L^ɤ0@�f�}�G2)a ŠI�~NBQ(-��"���y�u�9O�0GpN�t�SSN�A�������̧�q1��챁��V|�5�j�H���(�%i�LGq��x�WiM�
���Wk�"l@:��j���Z;ЍL�tUM}��A%���*}Oq��F�-2��L�N���d���c3���n�5�� lm�E�(Ʈ�<(��_��_��xm#z0���&��6鏋���+�b4Ƚ�pZ��t��A��D�&�\���i�[��ə��������^H���c3�UY^�W2���m����S�������7��G�����cp�����8|�7��G��+/:���-��@��aQCGM/`������B���8�;�F%�/����moN��	\y���૷\�����G���1x��7��7ނw���fW�Q�_X���se8����X�F�1PH�]���O�Dw!լ` x24�1�{�r3 ����J-n)Q��G[6x�"a��`�𔥂���$�C�2�H3���E�����\K��F�ʴP�L��h�l1��H�B�I�rc{
�>S\%OԊ��8���Ҵ��:�Ԟ¯2��s�̳�'8��JP��ů�/Ao;S�4|�d�rl�5���^�s�P�9�V�C=fYg^yr�<Yџ����a���<?&�t�6�X,{,mqz�պ�(Q�k�>bG�M
�c�FA�j��`��5����A��
TXȕJ7g�4�fx���,>+"���ɇ��@��(�Z�J��)u�h�$��V_�u����a�!�CJ#[c�z��j�S�i-%߼���5��l���T*άj��b��0���^;�����3� �����̃I�{
��Zb�X'�W9�rQ�B���$���=k��5�kka�>{`g�,�1Z��{�������&�{���;��n��:���ð�E-��k���ck¬�[K�q�9eqA���J�Q2�p���_�ʘ� pAs�p�'�7�g��O��k�����=�8<��[���.����]�M83ق�3iF!����pz.x)	Aް�05oDB6���	�W�P*�Xj�>+i8i�o`�X-9���t�����fK遃�8������qN��I�S�w��!����%A��S�͛N[�,:h��Y2��)�3�9�����߬����v��q�}by>�z�ߖF����",$�$}>]Eej�J�[ �X6y<Ӽ�\�a�
���`zVKD9C��3%�4{�����$>�2���{$߭q"7��ƀ�� ��0ݗd Y�T���a�m;�aV��� ����x���x�@�;-���N��x�be|�&vN�����'>
���7�w ~�������\u%\x`�������y�h�W�I�A�A �Za��ƹ�8����	�{D��ݜt:QW��|��ƽ_���� ��|��Ϟ='>8�k����be29�5��zO����0�{=��	G "K���G��ZO3� �ƨ�#�J�>DG@Q�4�c�"�eJxh���j+���`^�eR\���� ���c��}w�P\�PՆ{��]	��m����������N��i����i;��m�6�:GNoE>4�f��F���r�O�i+�ΜƏ<1{���{2o�����?C9�
]��Ȕ�刵=��hG�����R�W��J鐛���Y�u�+Q�Sb��`N��+�=�=��!,&��`�_�u��"�/��Z���7�nH^�ԍ+H��H��(���oCQ����lYix��#��B�H:y�CH�b|4>`�Q�Q�@�:S4f�WT�O��C���C�:f�E�
2�ƻܨ)Ill�����{�˓��W����U���ݎ���Lr�\ �W�w���2a�4�lF
��'9Q0�8���d��$�m/#���Mb.���-j��A�������̛���Vל!G4�p��F#g3��h�f/wq����׏<G>r!|���k�����8|� �9#�͉���95I	�'��"J�M<݆Js9G80qyo�1��X������2��_��x�e��C�{��Ͼ�L�G�vx��v�m㸈�Oty��p2��#��o'��Td/L�x����ny�0��>g�c,�]J�<,�+�+��0��X&e��r�\<Z*�
,�a���z�8p�m�G�R�Y	Ri���c|G+ÇE>0뢿\�����ʷf�ot����?d����{fJ���lr��#@!��0zQ�E}�M��/&�#���^�6�	}!�Iu���o�/��h)�<hP��_�*���p��(��G�g&�F�Fsϱ���[�.�8�?:ĸ���3lA�T�N�-�`�s_��
C��YS�3���x8$�2��o�H�Y��c)�k^as}B��4�-�z���
o�"�l�j�_���<4�3���w��/���/w��o�z3\�ephc��ov��J�W�;�mr{Pt���q}�F}�A���臨ࢍ1�����Wn�^y������퇟��=���2���l�y#��G<L�b��+^lX��W\:��䞉c��kE���(� 7��t�4�>-���6e~����,慚�w�xc6��.��S���Z��kQʱ֣���2s�9�,��l�M�Y��mZ`����0�{0C���	����D�J�r�O��rĹ]�A�[��t�2��9�n֋)Y ����Xlh�"��^M��2",ې�{0AO��I�I�p�P���>l��R	Hs'���&7i�ͺ�$��LL�f6���^�98��F��v�ufHD�@�/pa�yQˮ�͞��d���Ma�{Y�s�	 �B�=A��# ��2(�W^5!��#��ړZ������t�W� �14�Ĳ��4�`�~f�2��*��W$Ƥ�I�}�I�9�Z����MH�$@�4$��koD�+ �0�y��ѷ賊c�A8VV�'V|�Y�(0�O��3>&e�3��(ܫ�9���8����nq4��PzR�3��Sj�Xބ{�]�#&����9�&z�������yp� ��N��G��O�8_���g_�2��ppD�e$�SU�t�TH�p]~2IqJs��U-�u�=�|������x+���/�}���Q������߃M3�fmOݵ���^y# ��ͼ��m ��s��Lo�^���i�*�N�I/Z�@&cL5���.���L��>
�f�{���ۿع��e���\�r�1�p�� i��&ϐm�/�_6����1��9�/
������czE�W���-�L��'�#Ja���0V�Hǌ()#�
���VNo�~S:d�0�~��U��;ٳ��2�Nc	�0Ѷ�v�k�ژ�@�((�UX�OH>9Ol`z2�^���%=mP�H3Īy��T=sp�m���RR�@e�%��33�.Cl�ih�!X	O-�  o4O6�K1���s�F09ʼ���u�S_�;!#C��A=;�Ώ�<����SF=Ѵ8��������;ޠ��>i�q�������&���Ix��?|�q��ߺ�r�'���Q��B�<�i��-�i�7������-x���I:�庋/�k/=��`w�S��~��1�n��7߆�6O�d�g���g��Ago26�IdM��fO!~J>A7��lm	E�J\[S��T=��0�x��dC x+��~�;�9``��i�i�%�� 7�3�:N�q涙�м6õ���,*U�rd|�e�Gr�\K�a�R�Kh��)3w��ٔ 9݃	A�?Pe��SYꏴE�D>Oe�C�"��+�Hr�@E��jGp�yXF1��H<�� �BS���HJ�_W5t�ڒn�����x罡"$��F��`���Ea�z��
�#����3ʚ����Y tqh���I���H�h�&�Y>�N"�$�iyO�[5��}���yKg���R�-��a��1D���ӪW�SD��-9�z�E�Xl�	lAE4����
`�H�0�L�$$�#�e�=u��vo�<�*go��3�/0b���m�k?��ڞ�cW`yڬT�R�$qu���3)�0��NDZ(K���&Մ��0$�Դd���i��Y�ֆE?M�y��A�+?|�8|�[�΃�kc���9a�xUJ\P����&�k��"�f�$�ƶ�܄qk���\�]z	����'_~����_>��:�=j�����x#;���ͦ��?�:��Mw8��$[(��6q�₨��m�-ُdy�:+!4J�a���3��Pc̈�FbL&�<]Ԓ�����\P�Ff�4ww�&�Ww�6h37��=cp��i1sR��O�Td�̑���4Ð�Iy�0���⠥C���C:�� 4��0�y�p7���}��#��Nk aP	���Yq<f@	(���ؐ�Y{�|���(KΆ�.�f�mD&dF!,{!q��Dc�H�W��qQ�$q�g���^�U�E9�(��:j����M>�K��6�)i0����G:D�'6.Q�M�9y�7��֯�`<�
�Β�2t���y�~��~�:}��.�'���t��?~X;䍿����j���v�74��I�46� ۑΚP6^t"��ॣ���3ph�w]w5�uõ�O�x���_<��'��?��GcX����L&p��Z��+��W|8<�!�$�D�Z�y��UC�7�� 9�D��s��{e@���_�2���j�7��c?u�6��"�b�o�M�y�WfuV�w��x,W���4����[�����}E^��2S�
�aEL��iq�v��rH9�F��X��U,T�F�0Y$�V:/�n\[�B�-�K��!TIܨG�	c�o�vB}��"	꽗]?�ʖ��G�����ox�+�zHT���ƽ�&���t����w
�60�p��m�I��� Zcr�[S�Es�65]��ҰJ^C�5�k�$z��k���7��s��B��n��-�όQb tq׬P�5�zsk��,:(--�l��SF��&�I�ސB�:CŒV��y���m���� �n��|;X�����b���@��|ϧ�H�@Or�S����J��!�-x*�MОӝ��hYA�I�H0�P�iEX3t.�C�6���%�@:�^���ƙ{4-lu�N�����L��M�~�,�lB�g��M���;����!y�i��� 4�H�;d7���_t!���{����<��k�~	�z�	x�ͷ���:�wc��؆��c�� �-Ύ�
O�D�	�ëh��\Ie3�%y\}>Ӿ�w�J5\��=e�=<�T��c�����9턬���]3R	O�P7��A��������l׈��; o��Tа"�!�,2 �<+�T�)��ۃ;�aPpa�N<�7,����B�~�)/"��
���H�$+�a*�}�b�?R9��2@�A�	\n*v��$�6A	�|�UdMfo��Wy��~�B&��6�'��2ۀK1�Gϑ^�v�I� 'z��#:�<I�u[�
�Gd��َ*~�2t�eb��%^P��=ȇS��ß!cCL�tm�A�u_[����ys67x�Tt[�I^�L,��6�Fΐ��j��#���!�H�C����G�ʳMhXc��-�\<j�k�]�~�:�Wp
~��Q��_�
~p�8�����ހ~�պ�g,��]~��y�2��!�i�7I1y}���%|��>�80��4)$ �]aNC)����C���4���b3�l\O��� �|��б�񚰮�u�������[���^+��E�5d��= O;%L���i��x5
�߬�.�a/j����2� ���g�)��1o7��^���B�`�w�:hÞ~S�����Y�
W���dO�b�6D%(�"~��7�φ�߳-�
�J��?����r����1�y �K�#�a/ ?-���� V��4��H`"����I8o��A��sdQ2�--\S��`"��~!$�B�I�y�b���Ri���G�ꕚ��y6�����	$�p��T�~��6����b���Z5*��T�mɨf��߁	���E���M�R���~Z6�Q����쭁���J�	�R��U~EZ4���'�/7n�2�o�D��J�X!BJ�$�
�e���&LP���.�C�&!��g����oN�.~�^he��,�L �6���I�e�O�a���	s�q������>4�f2`W���a3���:����߸<������CϽ /��6|�	�n�|����m��ʤ1Ϊ9ZU�mc|{�vj��"�Ԡ��K���^��k)�z�;מZ�
HY9-9����y�h�����N�Zk��Ý�i���؏�7s"�I��Q���Le��b�����w-X��kJқB_�ʵ����E^�-O�۪ �)A�`-�"L�O�	��MC����q��J:�~�E�J94�(�2ڮ�ᮕM���@��tb
U���<0��c�s��۵t��䢨QA2�M��Ech5����*�	b��2�RZ"u1r��ӶӼ�-{��We��e��ش&ri�r*�e�v0'�x�>�&Q�6Q8�s�CD{ ���yI��
��I	]��&k�t-��N-:��ѣƿ�B'��%f�ӓ�#�L�� ���vy5�<T6�+�s|���?��Z�X��������ߺ�S��˯���=?�t��~�*�����>��z���5���3��㾌b�[�}x��ޘO��>�I����F�w�!��.iHhD:R6���T�� #�'-����(?w��@pm�WB�cpv�׼cc���y�p|4�f<K0��V���4;
524A����Y���W�[�eNE�T�",�i�a����g�C�I���'�E�m�M��"�E��aY�'�-�kv�R�Yo����O� �N�~��]cڋ���e�Ʒ�<�QN�遣ifCbV,���qX=S7��p��z�ׂ��ͫ!�e�j#���)��%��B#p����**of�Ƶ¶4..�݂ٗl/�&��aيQ��i)٪��C�  ��䕹����r|���Xc�;;M!�D��2�MHA;+�t�9|�����eҍ?�	�	U��Z.l�EQ��j����S�q�Az���4�@먐85������N�.a�a�A.b�`�R��TvzØn$6����L�C���E�y��1QRO�,�ƣ�������<N������/N�V�M�WZ�t'ΈO̶i��lʹ�m�����ww��dg���d}c3�(o��{�e����Ʀ��ˊ(�Bǅ�6�T�m�ƶ��E����5=�\r���[��WO�?<�,�����Ͻ /�{
N�hkk��8����w͊hc���Vn���x$��t��'ˈ��I�M���B��mkJY?�9��_��$5XA���wB�ľ�)EW�=ē)�:S�l`i�1U���.�eT�fD9�;�_�d�a��r�a%O8�x�T��*�Ll �s�8��0�M넋&��t�q��3<L~#"8���hE�<5ܕ�(�d^��^�@���n��;h��p�)������+m;wY����$��F��qB�4�F3�\f�A�a&�-'He��R9Z+�+�{0Z�w�f� ��6^����b<6`�A�]�i�T.�o���yC���G�����8��ܡ����Q�%|�M=���2BA)�Ie�4(�#q��wIXfE�b��ӭyO,�1�9ǫ~	�be��A���6:}g�u�xKJ�'ѐݕ�ҝ�д[���io��÷����	+�t(g��uOj��Cf�O��u�v�����uݕ�����ջ�����O��;���:����dm���H��5���C���t�}�A{�s����M(�e�e��2%F�g��ge��)�9=��g���7 ��c�J1k�)F´=�Y��Ǌ)���3�������L�����f�"a�
�"����<� �"Q��)~��D.#~9&ɁF���й[
 V{(���c���e]��B�4o�t�&�C�f���E���d%��"��h�B���%�ơ��=�U��~ �]\�
�cG�ˬ�K�diw�9��tk��a6ԿY���Z��fՠbٰ ѶQ�1�E��T��m�gu#j���,�t�����W�|�c��0�B�[��	�=$��"Lc�F��S�J�F'�Zy,����B��Qе>�$����������&F����6���������͒ׁ��[�^��n,�}_��H@"D�")Q�V�B
�ሙ	+ba�����G�#�`�Dh��㙱f�QP�D��(�"	. 	�$@ A\�@����n��r2�9y��[��ޫ��Я�r=��%��I��uM��B�����CZ���\&o'˹/���fL =p4M�ҏ��,] Qq�p.�Y׈����C^(0�.����;`�e׍C⺄�Fc��6'.0:¨��	B<��K���9�,���O�K��{�KOGH� ܱ��H���8�}��s6�ͬ�*L`:���i�{�%����&��d6�'��c����w�z#<x��pە�a�M�Y�Nx��#���0� V��"����3��@�B�ܽ��������&��}��W��>�է�3Ͻ?��<�t��/�κ��&m����"gO����-�ma��r�P<�W���P�@�y%HNN��@�F�t8K��,K�Zn����ԖT��	7KC�u�Q<����?a&�1h���>�f`پ��GU'+ؾ5�.UXvnd	5��~�ܽ�G>�2���Ӵ2�S�D0Gq��+#�"d���J�e�z�����eWq�>S�E��LO��o�4�ܵ1)�E�vB�Gۥ䳵|#�L�WH��`}�m�Caz�C��� �rgi�IG�=�`�󌣱]2���j�$Re�6܆f��i���T��x$>t���a�A��n;5�i�<iy����E+s�!�_4�^JA�Í{ս��A��8(Qْ$�F��j�L�Ok��js[�Lm����y���N�>$����铭n9����pq��s;�{�p��)L�]:�H8��������@!�5�ɴ��LV�2�,�9c�y��Ix�-o�w�� �g���
���𑧿	���/`��;+����y�`��g���
�M�'��0�]Oǝ.cpб�)L:kk�r�И5��E���a�&�m,X��ٓtVYUZ^�V,0�xɹQ͏ӺE���������G��rj��Ww ���E<A��;�8M��qF|��k���=��j���2D��h7���R�fH!/�F�Y�.�mю6P3 �a��a���T���x���	>�fAd�~}D����i<� (w�h��B7��i,X���8�����Muʰ|��
�ڵ�.G�a�'T��M*���j���q��k�Yma��ܰJ��'�Kh��e�@I�0�o�
R=�X�ez���7�Rh(�h�V���J�(��d�<i	X�I��8"Ր�5C$�Mc*X�q.0P[
9*�P��SÔ` �ߐ�2R����lp���R>V7��m�E��\ڏb���Kܠ9�m����G��֛�9t$�2��BΟ��^[Z�����R�SHv D�*.I!e09�`>TӰ�}9a0~��]ny��6�}�6�u�v'H� =L`�[���;0�mx������x=�[��
����#���n��*8����	��3����F\��f���Όm���yBU�pHaڀ�MW��?z�#��x~��+��g��O~���K?��x��N@�61gi2qh4�%r� ��FR��A��r��[��@Ƒ'3��S/ �{�V��A^�sIY,�����H�oo�'�J:��t�l|��f8:p�TƂf`�xȈ�XT���n\����4F���X4��?������H���=C�i�/�GC�'��hCqK��߳bߟ���q�ی�c�@��f��,��zED]&^P�/��#�C�Hma��~ҤC^[�,Bi��ibs�("�<+��1Mx6!�a5�@�Qv;��iSh��'��l�c��!��rs���C���F�G�n��:HJC�H��1��kN,�m��3�5�<-�<��@>0r���[����������$3��3�TW0�h�E�������^��?��p�4�z�
��{��|�Ax��;���	8a&��v-;�vH��]�E/�-68���$�"��sX��68���:յ��n��o���w��~�G�ٯ?���s�͟�?���ĉ`�8�ϸg`�Kx>�&�E~剏���ʿ  j
B����.H���0�UС��� ���5�r	CZ�(EzOi�]p� 0����}�dؐ�9&����@~R&��˲j���,'��F��$�+�SO�T�C%O���˩1�uLi<�uШ2���Z�㲬�O�ig0(f�쪮�~�u���hʡ��A�8���H�� x�I�%,j,�����:{S���@����8�aI�y�B�FY]��:k��J+�K�k+q���2(쩸��!�G
H5d��o#Y�I��n���%��FZ�$�D��t�X� .�zn�@J��b>*٭T�F�'�0�&�n�����Pp��t�*��8FF��, �m+��a���5\.�|
-�����Z�ܑ��mn�^�?kD[��BCy4/��LpE:H�&��7
�,C6� ��u����Nm�ٶ��l�������|���?��>�9x�m7�o?|<x��p��gaǽ!�FFnsdk��m0<i��bT��>c�Ʀ3��hȠ����m�锴{�^oy�M����x�W���:��W��/��%8?݆�I�伏������#~�^_��k�ɕx��*)�q�Pgf8�F�se'�A�?��7pJ���>(��X�7Iq, Y(�5��Z>V�����Q���K��]~4�����s�GEy\YUp��%�bL�Vpge��8�D~��|��^f��E�K�	�Y���훘��D&��Xj�S�[�{�w�XYG��̰�鐣����$׬��t��;���F��P�E^X	�>�`f(%���O�����<��eu�gq�%bfsm�2%a��T�R �,1邰y�3�0��3��eDw��<�Ȼ��,tzҩ)������"|�K߀���7��믂��{���{���n�+O���+���=������p=��ݐ#�6z!����4^��v�]39��>�������v��~>��S𱧾��ho�lkf����y�G�[C�XрS>���yx�/A�45l�K��򉃅���
�����n٥i�1�ܵ��	mg�ƙ��Z��n- ��F_z�$˒�e�E�^-]=��[��(ߗ|���T6�����'�Y�gL��^�C\�c���bu�rc����3I�L��j}:t3ˮ�U{���� 3!�ǫn
�i�/��6ǬU<X��Kp\6�R�)�r]nvT�'����cA:	�Ay?='3�	"j�B^K{�7y��:��B�c�𸱠�5&n�@y�dN ��!5iL���̱�B�5N��巌�JG�0�>h�*�����
�41G#%R���`Hр~��k�\Z�e��ADa�v�~_�/���Q���C�Z�ϰD�{��D�a�{���7.K�=��5 ��
ד����q��(>i�D�$]@�@3�WgrS
����Q�M�!%���ť��x����T��~��3��H�'������
�۳0o���d
ϟ����.��OíW��G�r���_��8{�tWv���<:�hs�Q8�h�IG45>t�~ݭ8�I�e�����Z���t����k�������u����G?�z�9x����}���n�"��G����'l�K��B�Z^�� ���C��#(*���K�K�83|�9[��=�Me.w.a�~r����y9�1��mN���lg@'�8�gea�������c�d%��z�z������ ���04&�|��@/kl=THi%��oe?�ţ�(�2��Ƨ=���|���82V�i�M}�4�vTɇ�:�����B�aT�f��BFם&"�/�����>���
��4L�:�;��D��:4�,ɖ¾���QO��d�T��'�m��Y�Ɉ� A��S-�񔡵�V,˝e��X�}����#��Q���H����bv�v��SW���ӧ�m��L�!�^�}�o��^|���}����G����G�k���]ڽ]0���3	͋����6�}ט�e���}g�z�NuF]�ޞ7��zr~����{���?|��_���c���/�{f���뼍��w^z!��w*�#O�M9��1���-A��#�/�{h��;���N�Ǎ�=�檲���*�&�z�[Y��rV�mz>�VCg�`�Z��mTQ�!�E�C 
�5���
�6T����8{ᰤ�佗����O36�:"6/�� $���#��%`��2������dt��;�C����E8��MN��-��'��0�!萶�MZ'P;!|ybσ��?��c;���*��ʴ0��c�ׇ��J$�rs�JK����]pB5.���j��[���=<���q� Q�>�Z/��S�CMx��F��(�e�R1-�4	N�nFD��ؾȅ���>��H
��4��kGfs�����3(�
��J,�/�.v�pZjq}Vw��)V��R%�0�d����x�=�jem�;ƥ���S  ���I����}>�p��l��MxM��$c�� }��������n��Jo�BE��Ϯ o�s��L�7<5�4�wa�9݅��/cj:Z\�f����gsx�[/�Ǿ�"�v�
��;n�ߺ�~x��w�['҆���d�k��̡o,��}d)�`��Uq,��c�{�!��=�-�t�������n�?��g�����]ڙ��[sf��×�}��~���`ٰ�!�3�Qi2� ��� 9?R1D �a[���oz�=q�&w-�!����[�p��l�k�w0��`ȷຑ�A��U���!�Z�z�*uRy�ţ|�gX�����8��hq)#ʙ&���8j��Z�����JX���1��.���?K����!~Z}5�+��r/���׮�L����W�"?5E[��K	!]�����*��l,kW|&.6��o�%�b���A������[\��-M�4���Z[S�e
p�'�{[���^�����u�om� �[f�M&�#��eL�+u��	��)]LÄ�VH�}�Yы
="�9:��~EB�`X)�:��Lې�0����П�h����
:ư��$�5;���]ؚO`k�s�IW����N��W��}��]�ڧ����'�����w�s��C�}7� Sge� ��G�"x���EB��ϼ1;��o!�W=�$��a{�K.�=����'��ux䮷��������لR��ސ��O���-ș)�7���Ȥ��sS��K��`���z�v�}ss$������Ms|5r��
�e�1�)&��d����2@���~9�� �H��[Ȥ����sѸ��$Y�n�䫂�lD-b=����IY �H�1��Pj���9��5�#�W��{ʾW����!l�l%Q��"���m��ymU���� Vg��2�IO[1E��K�a��� ��zB�ą��.%���H�i`֜�o���CT�w3�
�x܎r_�6S4}�V>saX&�+9��oӡ&D,��HYc���B��|��
� "���X��x#����T�B��ĔU$��ll�����(8����b���?�A�ì!���I��k�e�"�E���E�c�1+[֏�)��k�\�O�����-h΢�����.����6�&�M�@�a�G�.%e�I'��f�з����6WNniM�{Г��v�	<w~�����'��=�{���C�w�WN&�եq���~e��9��6�y��
�vK� $.�s��hb���p��i�g��8yf���5���)gD���wܐ�2��?G��7!$=��L�?Y\��JY��H�������j-�O��!�ŕ�R�1��pT�
�m����J���IM/��3�ڐ|�L-DY�8�?��*��8(q��K���5ƴ��Y�Oi�� �x�|���L�ǽ��|W+��4H�i��M���
�H64�3ƥ��� ��� I�cD�^N>k6�˲P�T~U��D����f͸��pꖣ�ot��H���:/u�BmN�/xܿF�4���O�g�'��6��L�L'z���$"�A���\ľj#QvF���F�6C������3N#h;}d��RN����N��E8��[0�ԏW��������?��v������;��N��<3��l��3u��8=�=D�������S�>��l,�4�h@��>�7�K��	��?���?�����w����K��u&_�{�!>�:O#�8���:N}��y�`�$}����K���$Pj�a4H��}mevU�k#�x/� �G��,����0�̳��,0���>}N����Ӈ5�� ���HY���8��xz�J=2���-��Ob��>�Շ|M�2�:e~�2~O���F1��(����U�y�c<����[�2�Ь�� or��9F�Om]jȘ���lϲ^p@���ߒXQ�&u�"NDҩ*���2G��qs�KG!�k�d[5�J��T"4<�r��%-��1�Ee�#ó]\i�Q�r8M'�iƸtG��f�)c�k����C�ã��6�1�0�F~�"�A���t�(����ͻ�$������S��g(�		i�X�-t���&$�T��J~ō�e���4��H���/��Hh.Ő�Y��7.?�{ж�I�#t�L�M��	F�c��q��[�NOç_k��?�U������_���C�����7��f]ƶ�C�1	
B<	j�K�����i���a��fH�f��}?�5�?����K/��拏Û�[�\+��>i�=�G��<�B��Im�QƁ�%y9o�n�{����萁��g���1\0��p?�'Χ�Qӯ��Hz �nd�����JY,�*�)a��v��}�k��7�L ��)킞6kz�f�PŽG��1}��4���؜�����I}��t&�.�?i����V-�ӄ��{�9l��j�7թ�/�F�%uZ{\j�`�V��o���,~0 �E���UyQT6R!Hy%%4�߈#�(̈́��+�.Ɣ� �[1�f�,��C4����cq�ς��Oژ��
����Y�&����O}�fp�����N�q�9vN��:������󟄛�����{��t��ѻ��N��ʼ�=W�$<�}�>�E|r���@�?�0'�w��3��ti���,���џ�O���7ν�-7m���<L&�ةynSY��cNtO���J��K���K2�ò���4���x�����+:� ̓`��%&3���A�s����¥�A�Ref�L^d��z�!0
A��VI��{���n�em�g���Jt�fy�vӇ׀wc�3k@h�%( ����P�������5���4u���Ȋu���-Cs��]7p=���yZC}=���8j^(m:[X�iĥZ*\Hl%�>J���(�>@���Å)Ϥ�)��|�{!|E���h܁@7���A����S�4�J�J�F/$A�T!D�VXd�Z�A�7��Eό���hm������M5��!L�`y�Q �R�k�KnKe,*<]Z�����~� �`���k��.E��ɢ7�ji�jI���>r?S��oz��l�,HN�m��!O�~��WzV�Y�"LSXj](e��d� 33%��:��^�`�W/��6+��N4So��-���n�M�z�
N4�p۝A�ka{gf�v�G�{��_\�'��p�矄w�~#�ɻ�o��V8�u.�-����{�!mC:78S=��*�'���C�aC�㊂�w�+�5�~����>_=��we�Q�΅��s	�#d��L� � j��3�$I-l��+*�)r.̩2�.�i 6��*�޲^I�*��꼼���l�Ǖ�7㊵!�(���$�*��S�"�+<$�G��e�z�#�'���K�[Q�Fǽ�̅�*e�����R���U�?��vs-�e�X��ɤL7Έ���yY>����iLd��).�ִ� t<��PΌA#�#�qJ�lg��u���S����O_:�t�3�0�/�c*�"-Nzꚛ��-e�<�b3���A�,CyW�(>!Mh*i��t�Z�R\�:������4�{볤@g��Gq��К����Ll��y�bL��c��A|	��+G�v��w�<���� ^���#Ͻ��=��[�w��V���`k���v�kSg�-�Q��Rc�ap�^C4X�h��đ�
�{Z�ө���'��u�?���)x��0~���\����tY�o��g�xH:]R9��"+�L�Ե�e`����&/Yl�\�_�=�q�;V�����<g@��e�>�FCz@P^��}h`��PZ"�j�!�Xj5,"���'���N�򒞧�kƷ1��H�IP4�*���@�N6�2_ZK��!ۗ����݀h3���H!����v�:8����4�KCF��،��qE���Hz~7���Awj��
����Nh!���dϑ�.
nR��4�m���c	ј���'H����Մ�h�n���գ����|X3H�H���i�~J�ʱ"�1I��I���0fcid}u��4�F��!��Dȷ>�k�	��4�y�4l�5`s>C2�aT�\P�t��	�������(ɻ�g�@!��k)� �z�G�n����7��L��i�V�̥����k;�*jm)ۓ^%T����iJ����C��0���ُ}�Z����F���$����{�نu匤�L1A# =I�-c�>�Ft���nÞm����˯�	_���~�q�-��? ���{��kO��Mӭf
��<^Rvq���������p�x�����W��z�5�އ	���'��֭k�d�)�٤)~�8d�Ҳߖ��6�5.4�E��:k%�:���W��'i��_��Mg�ZG���68�V��/yepACrVG��8����<����v��Q#�/FĦĐ�O����m�����!�8�|,z�Ѓ{_��Wf�~�Y�Eq�j�T�N�q.'�d ir����S�iA���B�"��
m1q�iq�X�3�=���hh�R�G%�+�E�Z&��{�!�E�Y�ûøW��ͼҘ@�t=2�JC��7�p�~j�΁�Rz�$	xYd�B���pM��<�6|�$]��,[,\�*=o���a��QHlkK��祴֡{ѭ�$�!����sXG�ӂ��`�0�2\���Ak�P���CǶ��u�	3��N������E��K?�O��p��~��{�w��r�W�؞��5���l��߆Q�3����-~���X�W�`�Rq.����>�v��>_�睾�&$�:/���MC��@�y?gH�R�pU}�B5I��E>��F�0 &��{�зO�`���_��	�R�U�~"|��)e�JY}��������[�A0��>yj���7xEd���٠
,� &`��dQFQ8A����!d#����g����ܘY6�l<�~��^�os���o�a{`�_I��T�����������ɒG���QՔ���r�X��}r[���`�Kv������e���3)�0�v��|ߙVI�E>c��I,ղ*q�'���С6�=R�!Z?���Ez�J6T@2�3��{�﬑��#(�&���Z|�/4)�+o��eH!�n�%�Ca�զ���X�յ8��p�l_6���%��M$ȼ�D�&���C������ͦXi�sԠ��bm7-=�4Ip�8�+�E`z��dG�ǿ=��\�����T�Yp�MԗrCq��`�H&�;��E�w������&J�~K3�r�tK����hRl;o���w!�]��$�`w
/��
|�;��?�����
�����[n�3��^8�/0�6������P�q�6Ƚ{�x�>�z1>��u¯�w�y���Jz�ǴI��������Cs�e�������X@ᵒ�m���� ��9~Ee9�{�N�^X��,�����xC��$���.*k�M�Л��R����!1��3�4��B^��l�Ƣ��"�)�
RA�_��q���	ʩ�ʲJ=}8 ɇ�i�v��~cq�eUɩ�o�vU�z��+��Z��1m���@a�Gv��<��%K��cQ�����~';�\|�B��آ���1Z�\竆��!HCH;=�s��M/f0)�B-��RY&==H�]
�G�aC4���
q��d���yq�C�d���gH2'�kC
���ZC��|n��a����2>���͊�Bi���c�NM}�ȝ���4�p#{.�X�a��~���?�2���߬#���[���O�>��}��/�����7ß<� ���[��k��Ԇ�m�{�Y
!��6��y\�Ӑ�p�s�[��~������&'�1�k��)�ɼ@��tK"�W� `iJu��L�'AdaW+V��a���y ���yr�6�C��#��fP� �p��4=�ak�~�l��W�M�n{��������q�i��W�ҼV�JN��rG-I���� ^`�c�r���'�t�
zZ&�x�u��Y�����Z�wLCe�R�v`�'�e+�/�1X������5���#�#�HȒ�h��W�{�y��:�A:�H&���[:,j�q�X�{�[����9�$��G4d	�'k��w�!�7-%�Iy��q��"��4^\?���V�Vw�@	��T�,P�E��9�x��Z=8�Z,X�`D�P5	�Յ��B���6~A�(�6��*Bp�V�)6	`z�M�>��r��~�Ἃ��m��p���E�UO)P
���J��(8B�\�2-��.A2�_t��ޥzB�U�_�����Ju6Z�(HZg�0G�2p֢mΈ�����7ɕ2��6��{���0�f�������7��3�ka>߆���<�/��;������,Xg5ۂ��*l��ʆU|:��A�
I�P��5p��g����ɫo��T���P!,ԑ��e� ܀#�nr2M�5r,I<*I, |��߻�1�>,���um|��,�w����f�Ѐ�f���ˋ�,��$E��dyf��<�4�~�y�Ò��U�I���(��I<�TⴲH\�L�5(�z�%�>kRfQiW*�?�ڥ�m��Z��zzp�}��b^@�f����R�7Ŧ���!� �CY�x�ir�"��.��zmH���x��:�>H#>���A�3Z��b� (�)k�ʔl�Y�N�KS�Lۼ�R�U_̆ͻ�ԋ�\˦C�	��lmIϛ�S!��1�6�3�Q���x�d)ҫt���٥��?f�=��8g^Ϛ;����s3	8�x������S�����������_{��9���(U&�d�<qx���=��D�Ӻ��{y�[n��-��lo7�S�t��K����F0��9Y�A�<�=O����0�1YRm�pX��Eԡ�G�4��!�^/����y(��$2:&`�������}�7���=:߁���1L��
���]�/��o�3+�`HX���0�"6F�I����'`JCe7��PY����Ċd�MZ٘�r��f�*��e�({�e$*�E�Kt]���'Y��!'���3��|�%ê&v�7MLt�XdY]/�n�o�A���~��@�� ]�F�T覤�!������6Jt�zQ��&�X�wfiu��_43:#{ސ0�i�'�����7F���J�-�H�D��t@;�y@�:7�߸D<��k���`S�6w�F�%��a���.7���(�Ȫ�u�kRp���5Rn$�	Y�4(��OԐ!/\���!'q�Gz���<a4��c7n��J�e���z6O��4�mN�Eu��?���w�wn���;tp�Ҧ�3��;1�;ۅ�^טmx����w�������p��)����P^eHF*y�<�9Jh�Ѐ����cgr�����	
h���L#.l�I�B�H2�9�=,]V댑�3�J�/WHg���@=�(S��_7h<5��4
��sf��}��Hl.P�0��	����g�2x �o��+����J�0�d��ie*��vi��`~
��[	"n��:�ȧC�=&v w��S���U@
ԧzH���wi�f�Y���!�0�d�QCq��<�7����}��JBK�c���`%2�X�|͙",���f<�@�ɝ�,��i��`)��L[g��5V�di���y2v�ޫя
��ґ�%}��q�"�b��c-�Ȑim0����-�ˠ(̻4�/3h�H�l�
؄���tkN����^�;�n;y�����¯=p;��X����m�㨤��Y���)ю���AZ83݆��m���E4j��3�t;WW�1���p..�!��b{���f��?$�8���T�� B�o3�W�.�K�(G�=��Q"���&�]2�@@�Y
ଓI��)coB������yKq"l�?M/���	LM������lF#�,�fHb��~%/ZvYxkrM���KI|�ls��M<$R�t�YȀ#o���+�I�w r���jPo��z�pJ�QK��� �Bk��f!a�O�����}�:AX!��Xz*W����>|��
d:lOc�Hb�85S_�P� V&V�:s^/T�V�"�:\��k��gj����LR�>h�&(�@^�x�ߖr�jk���ƍ��V��2%��@�Iݟ[�9�,�m>�e���ZQx�����O�r&i���-��bm0�3���q��dܐAe��K�oHǰ<�ӫ�i����?�0�*��Bwb��	�g-L��)�s���ˏ� �v�m�+��7_{@3���3�<{6�s�C�ےt��C�d�wc�ܼ���y����&d�I���2�j�MmJ�t�$H�~��#��J��8֘<�%f��F���2.GZ��ͣH��A�&+�u�I��[pp`��z�h}	� SB� (u�cD@��j���k�-pOZ�Q�=��IT\,�Sڅ=V�.�o����3#�S�P�b=)N6V�S�X�&����wm�*�*U.��P�7��HK(`�Ф���nD\\'��m*��%9%U/u�����<d��b�<ω�4�����m�IvC�涢ìt��Z�������~��.�7�� Ȑ��n��=$�ů�g+R�UR�������PM�� |F��2sīu�lQ�4n����Hc�8Yg��?���A#g�[`�.�7��fwm���o����[����	�z3��b�ӓ�:�hC�h�<Ӈ�*�:��w\�`����$�xB�a4����.�l���n�L=�@cy�)ur~&3�>l<��C�S��"�Rk"�39�>�%-��4t�1�#ǐ@|ok��B^�f?�;�L?�,Q�(�ٷ��G5rF�Cu�gDg�$���Uj*q8�Ը���)1�����Y�F�Tr�����f�z�]������>\�=>��Q�j-l{����IDXZ�wڂO��Y�7��mبZ�P�{�aD���O��}zhAi���hC�py��������{!��a�~��F^؇��k�q��Z`ĝ)�B�`�*�I�q��#q�2*��}$	����s�&����W���H������z:o~ Zr�����v����9;��Q��b�>�����/�R��2dX��0�]�ᆘ������H?�`�G	Ƹ|��ۍ�Ci��HKגJ�d�!�Lt�s@�ԡ��u*q0XFe �A����wy(�WI�5o
B�=��H�#�������@g�[���[-���v�9������ʲ�&����6or�j����=��p���}����>�z����0q���g��q�2�ű��4�O���@����f"3󻜍F�98���?	?z�U��O�>t�6�|n�A,���YL�7��Dʵ� MY��HW/�f�4�@<Aʻ��v1��#�t�hU0����}��� �$��>8�a���E�#|+>,�P��I�(pc�!
5��O�5Z>��`�Ez��)2Β�0ô8�O����w���+e�����1�q����t�����:&�����ź���xb!#��ƙ���Q�t&�mRʣ��o¯��[L�P��\Ҳu�$�;�z�}��eZ�|e�3N ���1��A��5�;n@|
��3���j�L��"�F֏���}x(r����A�YT��f{��R��}���C�y�N` �T*��B���ܴ�2��yl;�O3��������^�s����Y{�u#�v).^�3��t���w�>����o�S[�ׯ`���<�C�3�G_���\�f���l�Nڂz�3֘��ş��ǽ�cM�6�OQϲ�(�:���E��J����x��V�{�-��/ɫ�/���e��[;f��"�z��O��zF��1�Z!�"�B!�R<����A}���`F��W��@�������X�ވ|��ZgQH�O�6
cY)%�P"�"�Ӗ�q��gI\�r�8CH���X~L�
r��32f9S���	g2U2aא��?��4('�,�	������w�y��֢|��x/����F����@�&�&(J�u�p}����	���M|��0��O-,)h&3��I� �G_}Z���iy�F��ג��;�G̈	Rx qUR�kJ�KↅQ� ��������^2�,0؈�%��
O�e�z�Y�ei ���7j�%d�,�<���UR�㐪pi�jиF��dP�N�!y,�bZ��4B&�?N�2�?T<�ҳy������&�c[�4��osK���(Ȑ�67*ܦ�iM;�FYgk����u�?:����(c�k�L��݁?��_��>|�q���sꄓh�Awp��i�.�����gXL~�$V��&�'�Dk�w��'L�cB�حm���~������Ih&So<��[��	��L��=��4��r�pҍM̲_!K*��>#E�-�x5C�c�`�3������r�C���@Yn�F/����z��FOP�s�8Z$?��U�0@z�u�qF�������u��O���<��K�� 3�]�Ecj��WVeL��(�vT}P���;9�}ެK^:T�ð�]�d�ax��	/�垤k�Ć��8h�%�غ�**孋�-�<���!�.�s�
|�7��_�5�M��e=��Q��X�Oa�G�XgB�!=_|!���<�E��$��F��m$�������7md2L�eyONO��M��oP����8��i��*� ��/f�?;e��ؾ0��'��{n�?|�x��[��k��iG���g]f���,��#o%5��:C0�zOM
'_�ȭ	Jӫ,���W��Op��4M0����kWC戉����<<-Y+I�Ĺ�t�Q�-_m�|�$LD�
�u�a�h�@��q���U?�2��j��. ��{R��7�Y�j���qk��;&�}��cD\�R�+R��̈́����t���8�/yޘ��o����{��3��%�'��C��d��G���~�d���9�aq@�%�u?۰(�z �N		� 2�xXȀ�+�N̦��&��-���
Y�V�$�MI�HXkqwfJE����O1�����̍�bB01
/�����J��&�`�s�)��NP�6��|� �s#��'�7q�ܑ����Ʃ�/c�Ks�ɐ��?��(�ԝp�m{�z`�V�y#��
�dH��=(2�0�/����I"'K�>[���	�����b��vPPj�a&�c��9o��A�)���������w�yT"����}w�f�o
��ܜ��f����;���o����9�H��z�p�M�mq����&��	�1��z�ț���xt&������܅��3����ß��[r[S�v�mh��7{�aρ�qd
�9�oT���ǪR-��?<L�R�?L���L��'��t��v,˿�K��J|0�3��{F��M����%�3�!	��Z	��Ž LRy0JY? �E(��S���kT��wC�+ڪ�����*�X�I���)?��%2=Kx�L@׍`��o)��������3��gͲLhE�9����1:¼����܀��Q�y����Z6��"ce(�ByP��n@�9��(����Ѥ��������zJN\�p�%� �t_jP|^Ę`���+,՛���9/6V(͕�����1]�p}��ݿJ2�⛹7jw��� f�����)�=ל�<�(��o�;�^��]����P�6�G9υ��H�-����E0AO�<�?��7�X}�L�|�?�����?�,�N�t��mh�I�qo�s�tM> �}eE�L�m���'6�0h��,��S�a�>�k4���|g4�ڈC�ʧ��4V�#�8B;��;3����R�7ח~c@�4��!]�{P���w��E;��n�Ә긌E�����<K �3�WlH=�D:��Lsؤ}�,����/ɩ���s�|�YK�?7�M�FoL�#`P�1��*K�2X]���^Xf�Qs�
ڂE�b^����g����&�C+�[�x"q�{?*@����J�D[��*�#�m�
΂��1��aL��a�'80��6;�%��ujn/�����c6��s `ߊ<���
�r-�I�|BoX��o=+�NO��҂�Mb�"؂��#t3KI����i�6�RY�=mȖrZ�_���S�&�] ~YX.��d��U��&7ڹn��!H��I��s%�{shfn�r��=�%�ɣm��[��(����a{vn�Ҽ����x�cp��ga�����̼�hnᙔ����mmio�M"c��F�7p��I��hh�K4u7�<�����W}櫰{�4LNN��z�@:B�}�'�����
4�#d>9����&L����J��M��y8�n�7�(�9s�$������H�t�¢&���F�"C-�<�t	�Nq��`}D^4$���Jz�'Y%� I�8��|��8F�Uܡ'n��v �F�"�D�E���|
�y���`�."�r>���HR���7��N�	���%��R�G$�����q�m p<����w3��d�|�}D�{��}c�5A���ȼ -Y�6����KI�9��đ3��E�Q���
PМ;�
@�r?�,�0�OV *9��)ȩq_� �bI�$����pg��)3�U�:��=��w��BN�����k�N�x쮻�������S'v���v�;]�����F!�'X�|���k���$��&51&H�liO��w��W�܅�|�k�g� <w�u����n|>|j�D��t�7�D�|��$]��~_Rq9�Ą�Vբ�=��j�DGF�c��R �d���x(e�E�[�!1+T��O%��OI����Sϡ�d����hIgc:�F���d�vn	F����U���rCy<�����w(Ge݂6��1�[�9��Ft��(��57����)��a_kp�Nу�a�.���FYKN�XЀ�z�r�M]��E�� ��7,!@7��P��s��{d�cIǩLd��*��H7@��p b1e'ӎ0mr�6TOo`�Q���-k��ei��U�S¤`�t}�������1��(��
��,A~_V bN��=P�5�o�ސɁ�;E}`��¥�IE����kB�r����9���A�h� �8o+�~z�%�,�g$)>������tAtk���X�(�$�!LPȾN����E�"���L y�pW�&����s�.�t5m���yc>�7a޴S؛�m���3��x�<ܼs~��w�o>� ���w�m�^''��vY�;�O�4���䩨�0[|��62�|�'*ZM�pDO+����4���}�Q��ߺ{��?�}���o?�9��n�뙳��+}��D�/Kܷ�|Z'v�����Tz��`��8�A)b ����F*LV���Ko��\���he��/����=���h$�F\�<��q������<����a6�}���<B%K���I��Ckϧ��,gi�V&�3�ĥ2���#Aá�O�+���.���vi��t%�������-����(B.���Oг��4E��/��e)�PFץ�q��3A��ӻu��A;��E-#�6\n�/&�71�]�C����'T(��yJ����X�u�0�yEi��,C�	D���aLfsI�	�y��=#�~���0,��?�j!��3��| �l���tl������������:��]���ޘ5^��L����uq�x%���o�w�{<t��p����/g~q�c2�{	q�dʼ�u%C�8��"ʚM�81&����h�H+�(`�g>됛:E�]؅�>�<���}>��w`��Lv�HO�4��')M�j�ȇ�s��qUZ��
0rdc�+�_3*Uo6?m{��{�P�8�-d��c�C�%:���=���<xA�%��DC^%ӧ�9���˗�H����}�:�
f L�d=8l8P��|�b`ӧP^��~��i�A��"�΁{�,]5}y�"��p��U,��-�,r�/4��|7|��y�]i����s~/Y���mA���j����g��v�B��Y�=����xi%�w�/g�١>Gf�ݏ�&��C���E��!Z��D�$z#ڿ�7���F�2b�W�VI����T�7��f���x�BC�uaݧO�?@H�Q\�Ddة��L��c�>I��\@D��L�|�[�5��`�:a��om�:����	�aK������6}�fm��Sp�^���`��X�êƜ�)6��t2�@�Ȍ	�z�J ·�."�!/��8��
d�����w't�J
�����,�lp(
�u�G���wl��m��:bo~�'VX��b�E�I3ق�d^��pnr�]�+�p��mx����|;<z�p������Sݲ�d��<�6v�e8#�lI$l6"��<6��q2�}h�e�֦��P	y��+�g;���ν���7�cO>	�z�9����arf�ɩ���r4x�M2!���(�!B�f��d�rv`�c��9E#4!4��#�rC^�eB�w���S�E7dk.֍��˒� H��>��������ߎwR9$I`���gY'y4riZ[�AH�H����a�����w��H�P&��G�(}�5ʓ(�5"�qDW�8e�2���.�
~}�*�A������Q>~*}���]�[���Z�gSxP�E*���q�w�p�ם%',#��$t^��a�7dӔ�L�!&�W}v9CC�(��Q���:�ږȽ���j��
�~W_����=�bY�sB�!�0��[�*�`���[H(�Y�(aR���@�Mi�J�d��EZ�s��0���g����L�,IV!��V��-���6�d�=Ob��b=�o��:m1v�i�К	����O^���83�g�R�z�x����=� <x��p�W����*��%��d�ʹ�E����o�)4d2r�;��O�����[�5�n��������|�ix��?����mN���ɀ�	�MХb��d�ԆѰ8� ��|��K�t�Y�K4�4�  ��`��J����xš ���j������(Y,����7�B���-EF��*T����C�к�W�q���q]j8ni��"n�����dh��o�7"�����&���b��+dyd/Ao�8X�^݃��Ͳ4A�'��ȢYlR��[S:�u��p"E�2����x�t5��Т��*G�&�0#~%�,��-O82��g���2N+�
4��'�e�Ou�Q�Q�a}��
i��aH��)��Y�n�ǴOR)���w^8IK?H:R��RD��G�m(BW����a6�9��
��@�/�֔��ϖQ1�tg���Rq6�A�A�o,��`mQZa�H4,���6n�S����	�e�+]�o���|Y�wo�4p�B7�:�]q%<x�U��M7�����V���Y8yf��������j��}� �����J|#��aせp&���5�m&�^3\YS�uA���s��|������x��٫���'N����30��+~[���?�҄�L�E�2E�?ߔ�Qy�<5�"5�;p]*��Z[z y��r��o���M]��_���٢��u���C�G244��\}�q��m�?}��)i��aP�)��Wʒ��E�Q�S*�ͧ�g�|R%T7��8��U�I�Y���h�K����7���'������ky�4cv+�	�e�X���!����&WE� �e�N��2��|	GR����Xa���iYO;V�:XX�ޙ>3�ޤq�rb2���&Y_�A��Ll	�P�G`���}�+�8�*aL�0݀�	�&��>�uN�§�O5z���E��h���� �N�؝�������y�-���y���7����L�wh�qp�������Go\DkD�S���hpD7M�,��qN���>��s���/�G��%��3߆����t��ɫOôC`�s5�p�x�<��Ƣ�������!�:(|���m��kYY�}��+Z���#@�PG�����,�1܂�S�e_�'�V�o)�"a�t��U�W�.�eK�@�5���r����o�B�cL��p�f��3�Z.���bI�b} �5�o�@�AU�m��h$n��!(��
��>/(#3��t_h���7�XT��ѹ��m�(�Iq���R�닣�G�T�(��Z�
��8�OK�R��Z\~��&
܅�I����G��Z��,���+���K�7����F[h!������r�`���Zz�M�Fc-�ԙ�>@�Wa�8�� S.'�t"�2̦a�%A>j��љLh�a;���FO�b� s%A�w������1`�lN�}m�,���3YH��`�w0�n�V�dPC3�Ŧ�p�c���Cw��_�)�v�up��ih�~��n�Ovq����s@h���6�7	�7M��n"#�z]�����yј���w�����_�~�qx��О�85�ɕ'`˿?m�<��/�{ݘ����"��[�@��SY�I��D�K����Ȥ�"}n��PX���n���n�~�B�C����-l���O苬M�o4}�dr	�Y[��tK+S�O�X��'�B$�U���zT\F����ߵ�a}�� �B�3&C�d���^��neG@��АÐt��%���`��1�T���㍩��S.�K�o!p���FK����K�q��f� ��3����m��a�EtVdj8_�Δds�#a!p���+����b[�ɲ��+{��dZ��L(�o�7�ض�7fh�ӊ�$�%c�8�.s�K�������ǿ�^-L��`.�u�@FO��ז7��A�j�̗k��z������-*&GW��Ѷ�³']�W�|>������O×�����;[0�t�qcj��P�=�2�7��6B��ǦE���  ��IDAT6�6}e�&F1� y3Ȭw�ss_@��"ǆV��q��v��0櫬��X>�Ȕ0,ӫ�,� FK����>�M��0F���!4]��ÿ���c�K��^�����ˁ�,�~�e�>���3�\�~�(����$�t�p�Y\ۨ�?H�|(?.�W3K���ؚ����@�8@5��o���Y�e!@�~d?ˢ��$���⡖	;�IV(ۢX���jy%�9r`���9��TFEF��6���Hw��"!k<��a�����8������ꃁ�1�&h����(q���A �G
g�-��$��2r:Kw�"(o��8"��[o�����蛣���̠7I/EȮ	̸���M:�ǰ���C��|׈����Z��1�W ���ד�{�ȨA�7}4ʟqJ�(��1�Iq���:�f�7�F�o���9o�-�O{��`�8:0���@��,	�	7ܜ�������x��jv�"L����s;�aS������Sd�y/��n;��i�{���Ĺ���6�y�"<��ß�"��S߄�ν�譓'a��Y�vϴ8�����1�晫�!�"��"��(��J�#uS1N����~���I�
XV�D/WB�M����H����q�A&kR����!�@�%{��fD��l�M�DV=p���8����H��ce!��S�Ui�V+�,��,� OO؁��2.��t��yQ��x>q1����i����&�	�&&}��jM�e��kxyC7�^�4`�W3nL: 6��Ǽ�0�0]��l�����1�;���0z��	�g_g=��2Xw�ͩ�y�۔iD�B��F��~G������&yt+.Bxj�v��3�i�eD1�*��I��k�����{�<-4�ym0��G�z����9�l0��q��Ά�Mh��ve����_�g��|��O����`�"̦[p��+a:�`����p��OLХ���~�+�ް	�<�R�)ǈ�B�-_�ێ�yB����s�M�a6�
�T3�:��mn'JMdނ��)a�N����*�V[�R�]���|0"�0��|&Y�~������(eХ�ʾ\:[ɹ��2)�T*�G���OC��:�nVo�����&!?�,�+�l�������oJ�n� ���8��3Z:��Z�r��������%�D�ZY�\-�u���5u��6g�t�f&�k����+�o�Nɦݤ���l�$̐�ih���m��fk=v�k�����naWZ��S�2JT~�&h�4}�h8���W�*a,�2�~j��)��%��(����Q�j:.IpU�I����i�Ҵ�H-T���4�t���)���m �7+�&����}�c���<B�ͳ>W�!����!�SS�)��9z����q��#�U���&_��T"�N�Ҵ*k��Or b�0�6�����o�%w�&lj�x���mf��������n�nֆ:],��}X�1����bă��`0Ҧr�LCʁ,8hp�`˜�gд�Y��������1|ꩯ���|���g|��[gNÙƄ�<ўz�"I�LP�hn4\a���9K�%	a�G�36��NE��%��`,�}w*ik��.�����Q���Pt��ɐ�ܬ'8���vz�`��mt�2��@��z��d��~�9CĿ˨��i}=dzeH=' "h�"C0R�X9~R�Qh��gi�P���v�z�p��L��8ٷ$N�=d���N���M�39�/�P�q�p����;�o3´���yL�m�'����~������&��ż�q-��_f�Y��*�q�0x���|S!�/���eL��\7��㊾�j <	|iQ$��L�=�9Ix����D�(���C#���*I�5�����y�8�u�9�������(/��f�����^�i}�{U��� _�tF"sc�չ�G�N�&>\��{�S��y�q���Χ��W����|��O����<�x�\<�%�t��+�D�t2	y�|���>ɒ9 ��޹�T�������\S��e�7gzr�
_#�y�t�c��6Y�$�)7�7d��u�;�D��8F����֧��ɭ}m�2k�!��Z=��o�W}8�k��e�I瀪Z:~ы�'��ñ�T�Oc.�_�y����
�j��$���i}���� (��g����ō@!-zU�^�m�ӅJ9i6��[�O�#�I��cDhm�l��n��.���6�߻�$ �(��k��G��3Z0���v#
�� �وC����6IA�)���O���)⤰�~��C���(>2Ne�4N(w���8��U�Y��A	�S7�wtv,��|����Z>^f4y�1:D (!א���B��M�vt,ݢ��<X[�r�ڼ�%�(!8~��A����u͑iPQ��X᫥��7
�&�e�oUC"،�Cڵ�p�(��K*�G���%��0�^��Ql�6>���M�?]�,~���v�����������h����|>�6�+_c}�@�Q��l]`ǲ<�1a'�楣�m��n<���O��
��O���S؝n��ӧ`��6L�`H�niB���_GM���6���W7�ln&�*�M�t��3TfI.H��������Q��6�h���[�˵��ky-$��c8d ���n���>�e#M��*�IYOI�ÔqT� �m"qL�֔�-_�G�(M�8��Qj5*�b8CO��C�mw%_�(�*�ZY�1DH*��~P�,������ĺ��"xaJ�},Tu�3�C�"�EDq�e}�/i`��
��4�ˀ�0�IrK��%�#�r`��a4��Ԩ�o]�����Y�D�}�:O�̐\r�Ӽ�5j����A^�11�e�|������1o�Gx��W�y�l7q��:}���&'��#�G�ͬ��H&� �"�?�����ok�W�65&a�g�~�&���M��K��xC�f��� _}�%�w��4|�߂Ν�t�3p��4W��������F�������"ߠi�l��U���>l ý���c�5p�,~?����&CZ������;��g0����2h�V|��[��@+dRE.�zOU'��T��*�寀U~�J�[7`�����H�D�BC�e�pzr��2��?�|�O���k5��h����{�_��u���8���+�S���Y�:s{�h�o�y+ڼ.�(<�||?m�u� ��������c�$WnQ��q�����q�$9��R%�n:�I��`�qx��F�,- c���L�$�֙~��pg��j�4 
�N-ê��F@��P˻��2�eˢPpj*����G�Z�����h�ևy��bb:�d���1��޼9�e�䓞6��/��o�]>$�/�e�샀@�[��<� �m-"F�:�b&���R �J�)�i���	�JKR�pm�����M�E��7��Z�4��oT4�?|k­4�"y��`����~���߃v�<�;�&��Z�r�I3	��l\?Q1�o�#FQ�i���43N#3D2�h�F��K{~s�{��S؃-��k��񧟁�	��/���_ 8y
v�=Wx����M�4�D��@#q@%�Ȉ�&]S�Q�0c��1��Z�;�����bks�͍�Z�@�.�e�6̀���3��|�3=�UzI�<�70�����~�h��J�V���ViV�Q2��05���Y� ��T���.��F̵8V�����>"__�}qcp(Ƅ�{�o��0�)�C<�cF>"å2M��@.+'����W�O����zb�QJ˂Q�͍�s��QVm������!���km�p���J�%�9*=$h�Bx�M�<Y^�$]��� ��U�Q!�`~�b�~�B6����5"ú��ML�h���#�DΨ�m�ڽ�����7о�{�ހW߸ 7o]���#2�G��O����mx�'�<B�F�N|� �?����x��D�7:�����f�~��W��O~���/��.���I���8����$��e�d���P�y�3)��6*��傁Χ>Cj0D�*�� S�ޓ\�Z4h?�/K�c���7a8����G�K��!�\^�!��kTʤr��r-/{�y�U`?=�P�SIX�Y�ξ|˖I��SHl
��j*��Z�Z���<_Wei"o2���+�9Sy#�A�RE9G���c�]J'g�߇'<���B� �y���7�h�Հ#ᲦΪm<P�	pRB���2)&Wڬ`1�e�����CEΪ��DghjT�և!��nȌS`U�N2�j��"0���/QA �EA��u���}l����"������;2lٲ4�����5�@���PI_�ITm�8	�Z=&��4�N��A��\P��ue�o�򍼰0���է�zJ��X�����cX8�
�)x9]BY�#Gi���Ħ���;[�hA��UYǶ�q��d�
�Q�#!�H�������n��3����u�p��6�:���v9g3����g������㮷 loC���#��ͷ������o
���%����M���cHb��������+��+�>��7��z^��/`��wrz��<�$��ƴ�Pÿ��+��I$M�B��`�Q�
[��x�NC:���!֘Z}�Ȍ#��	cdh-P$-�y� m<,^������}`T�t2ذ,���L��"  rC��� ;�,�ě�ҭ��
s���T�qB_a�*�����%�$t"Z1:�~C�^�,G�1u��WUq�U�!��x�8�g�.���oI?����r>iE
)�gHq$�eq19N(ȴ,L�!rD��H=	7�ǽA)�4��c��m����ၫ������(-��/G�|���P�X�S�l(��C��rVK�b[�҄�nA�&Y��Gk���ZJ�Ҁu��&x��q��&x6��i��9�uӽ�p��I�����y?\s�*�O�׉l�O���L��洌yԁ�����[䷃�H�1Y�o�qh��1	my��מ���g���~���K?�W�<�V[g�a�{Ԙ�731��6�Y�����=~�˸]:�Y&��㬐j7MV	��u�g`��Y�BY��3��g�y��h>q�`��}�?}����0AʃEd!~��m�'�gD=(�z��{I�v�B�g�?Qբ��!���,���dXߊ��}q4^�7�鳾�_�X�=a�o�4��r��+�f��o,�zӻ��,do_���Ot��r��S{�w��`_� jˊ�i�z���3(���,��驔^K=�Ʀ7��fBڀ-D����لc�h&{>�Cp3���u	����~AD̗8�V'�Q��������R}R� �Gn4&a��\K�?��4�������P~���V�W�rS�J�$l�4\�E�a*qeƂ�kZqt�b됲�l�f��;ݟB�@�a?++׀Br��X��{�@v����:f��n��(�'' F�]�KW��U-�f;�f��ӂ`cc�6�׌�5������|�[���~�7����^���<���f��#�c��gw����$B�=f�n���)�AJ��4)[�`��:��L�y�pN>&]����9|�g?�~��W�{�}�簻����
������]ڐ��_�DE!�録b�7;��,4�&D��ۅt7�)�s�4?΅)��%{BΊ�<r@+"2�8�༨�3�$���'��-"㚸�����v���o��t����cXp>'����s;D�����L)m"�CqC��X�B,�.B�cz�бgH��a�Q�O��pxJ=��0"���6w%H۴��0��~_w�j}�P���}ej�"Y�^��0�9��"r�M�9O�{�)��|t?��h��%�0����q��zX��m��\�t9��#�d��նj��E�ݼg�R+�H�*r~: k���y�J=�.��J}��Z��ܩ=�R�3�B%M��B6�k��F�����L��;w:��c&���?ΐ}�g����=�]��.x��ý�^��&0ٚ�:�|6����D�;M#��x=���l�X�@ܔoH�&�����+�w�K�~���?�x�k��=غ�j�9s
N^���,1&M|~�b��#�<F3?��ͷ�XH8Rz�ی��Y�;����4������$�Wqė�T$���탖׼�i<�"H���xC֦+��課���j�{�z�<���0�V�%DN\�ep��(������cz>)�	�����>EE"g$��@�D��ɒ���0(�_M%�C=�~��)@�;㊾�3���SO��2Fb)����v��]��/e�������MP?<؏�Uc���v�H$��M�& ��w���eckT���mLq�؁{���66Y`I>Mp�7�*���N���ލ��D+��n#��q��mZ��PWU��"�͟��E�B�|4	�d����Ҽ(}�i݁T��d,腄���Y#�z܂�L��	e�a,�h���ie�@\c\���_������������k*��W�6$�cr"���]�f_1.��.�q������$���oӇ"�NħF;�"�YJl�K��h�W$��w$i6Jl%�p��G��F��جj�,����CA��e�H�"�"���N6����iӉ�~�C/��r�\F�/H�d�d^�V";eȓ�����.{Kֿ1ܛ���x��7�&��s��=��]0w�ƓSx�7���~���঳�������q�����<��e�ΈVl`����#�'��(�R7��L���pz����sO>��G?O��}xs��|��ӷ���`�d���YS�.�&ob��x�p�̞88�b5��ȃBƃn�9g�1ܦ���Q?,!�)kD���G���Z-�*����i�-6����X[',��Qv���
��>�,�"l��c�hZz����V(�^��/�D�QPo 衃P"6���G�1��ӬR]�whqC�h\I�H\���[2�rF�Gp�(~�o��t��e�~��q(�J�V������O��m�(ʊ�Ox?aP_a�DwH:��kX���e�=	��{���C���\��r�XC�]l�^S�'���؛y��ADyu�즱�#AP��Tؙԋs��� Z=��eK���"/jJoh*|nQ�"Tc��x�6��r�v��ws��HD'�G�}i�6��z��<~:O�y�����=ԅ�^����kN�;�~���ᱻ�3;�;��l������Pm�Mz�!c��o���7i?<�7~o%�C������Ζ�����c��瞀�����+��������t
�!���1������G����4�=u4Z78�D��-�3@h:�+���C�i���@���R�1�d�}ڰz~�cX>���c�B���VȢ�
�E��O��̫_V\�,�?(�B�M�"�WWY~��@���RO_\~��Z=�k��5���pS	��p�.���ٳt�q'�u���V������J�%M�RP�8����px����y�����?���'G���8�σFό��D���\P\ �$H$@����>�>�*�~��U���w�nw��%+�*��<U�6���B�쏌����I80[z1a-�i[h��̗l}|N�`�= O���q�����ɲ��ȇՖ���m�����d\�����}�w�#�����kQ��B���OΣe�Z�<o�����*�ҋM�H�d *"S�zę3�i	9�<��G>9+aQ�ˋ��n�|H�0>���%�0a�3Êj�};eT�A�� O�4T��sƢ��ʡR��ό=��b!S	b�|�z,x��p\���Rjv}�4?�~^Y��V�̡׌�Z}�{q�y�� �vd��ωcPuh�6ڨ�b��F�#��ਦg�{��6�ūj ,r^,'V
I����0�,֙5�_��|}��E�="�Ji�Fyz�r/��#�a48�S'�%
�E���O���	o�1�Q/�.����g�F�D��|W��L���[ڝ��+R�q�ӯ�����(}��|��t��1����Ǽi��d.dH�@�syj ��qy2<��;�]0�]4�}�Bm�#7������S_�6��/}����_���x����m��z<.�w��
לl?�4v�.�M67���� Nٶ���M5k���d�>&�V�k���1;�Jo������ �Dpυ�s���鲖5`�/����5\H���W�w�]D���d@F���!Ս�	�o�|9���3�"�I�T����i(h'B5D��!����
R�Kj�e����+�	����R�n���G-�1�#Q����{��NDf[���������{�I���#u��v�OE��r��Rt���Yvni9��n�o��n�4�q��ڀz!O%�Ҙg�A�����o>]Ή�z3!��=կ��G�~������=�?��p�`�Ġ!7�Oº���Vn�����4ﻳ���W�w?�a��������'iխɟl�{TF�g5:�DK�C]�3���T|!�}���!$���K!���QV�!�ъ�o<=�×�3_�*}ꩯ�W~��d�	�;G����ʍ��kzy���_�.�yF�݉s�	Ỵ��kp�0��|�vrٟ�6{�va����C�z륧�"�ك-�a.�S@).f`�7���R��õ�,͘E�-n�8�2���U&��\��C�������C+/e��sl�j>�{b=�$��A�D@,Hux�F�e]��e�'֜���lE�<�E�_���qn4��ƅ�v��&��s��+�O���O+���iB��`� �I�כ�<>P�Z�sF*,˙ ���p9y����)���ڎ���A(t�#���A����on����O�KJM77o������e�����B��������5��jmb����&蛃kA+��4����-zи(O �^V��Q�%e��.��+ۚXLLz��֊y��(z�ܽ8 iފ�IC�Xs�*G�._$8�y���f���<'���vyaF��JS�қ�\�w;K�$��z��{I��KsE���1�F\z�J	}]��c���������G~�-������_�U��;�No�y��>x'|x�|��d�����̓y�َq�i�6s�==�n���,qܯ�B�&O�{�������П~�����H??��F�o���-����@�����	ˋvS����"P.h�$��7e�/��K�� q0H�͗�U�����Q1�Ǝ����	�W���\�8�p6��<�3�MCW0�7T�������ZcE/��4��A!#����Uza��Q�#|�w��G�72��6�ԇ�r�^�O},M���'�ӎԗ֡���8�v��lm��U�@����
N����Ѩq@7&c���\U?47�Ā����r 3.5>��s%ۄ��X�p���,�OHtK%��sf���뢫�8�+��*A�F�ܿ�>�I��:DȢz ��;AF` �]'�4�۟ B����HC�	���-�!�b����x��p%��w�Ozz[wD��w��Ư�?���ӻ�x�n�o]��y�&�%�G)3o�\���>g8��$�%��?N�(�<~�y��+��m]/��}�;ߧ���_��|��ҽ7���ZߺI�۴4n�y�sX���Q��o�+<]��.�m�Y�Ӡ'*�6�������z)�����z�I���Y��̗�}���S��x4^��l� CU�e9���bLݒ�Bf���9]��툳�=ۧ�98�[B�5f�����e�y��R�����S.��
�x�����iĩ��
�	�F�<�h�"u�����>�7��ek؄��[է�;Zv�ŀ�ר�~ ��z+#���$��T�arTߜ�SR��`I֨��"�����h���9:75�����k(�w�j�ϻ'����\?O��z;�D+�6,M��o�R>��G+ '�#��_(&P�M��P���Q�'�Q���~�YMy/���0���!�2T0���+���}}�|*+vPsF:��)B�[p�,obB��xcb!�qZ�4��tH���߅�N�f�~��ˮ��IfS)s��7à��I�W�-b���F���h4��M@�p��}68�Hݸ`9��?��&8�tkz�����=zߍ��[�y��?���}����;4F��'����p�F�B6�Q�n�V����|����D*��c'����#����m݄�V4��܏^�?���?�y��^���1ݸ}���K7�9���]���l>�sy��~�㌣�O����_��x΋�YO���{�m�2p0VP�;�[�a�Qc��<���HD�P��;m8��U}�:3��yi�D��>`���耊�[����q�@���L�~�*e��+N�P�F�ö!.�#��{�bʫ��q����Y�Z�
�Ώ��ؠ/�Qn�>o��V�K�����z=�s�v��g���>��s��q2�[�o��J���G5��_����X�x��UW��A�F�M�Cs _���\mO�_b_(�Q��i�Ϻ�-�ʩ,�hQ89�F�EP��&��$eq��3L�t�.�Ti۪����OJݜl�	G���gِ���塣�>�$����*���[�w�"����a(s~��6��ד��x�?�7��͚�&�\^���>�;ҹ���W^S��m}���Z;z󡧿�ڳ�o>�W�����~�pظy똎n>FG�5�~,k8	d�y��V��2]�s��-���h�.;*�~9��g*�\��E�<T���S:_�O�����m��JК��~m��;�e�rg�^[Qm�j۲����k����|�����L�@�>eOk�g��>-�(��%R���VN�-�O"s���k㐢����ũ�L{������O�|U#�@ۛ�ڞ:�c�+_Prb��&�����T�8�*�.����}��
O�^��g����lx�V�f����qO_��!]���
�CY=.c�R�Xo���i�c���:tb��i��~��ݸ9�r8�\�Y�>��7:��e�����"����@h4/V�����xR�_z�MuT���-��qZ�+�3����׮�C_�3�vX�y����e&XO�t[`�A�>[���}pS������*8di�9�X��U�}�,�� �����`�$*<AԘ8���<P^X2�2B^���*0�ȫp�՞��£����h4���j�X�-�)�,�M�ld�QG��1%8���ɉ�(��[i�˛%��>.d���o��I������!�������/��~��������wҍ�4Q�O��oF�"ȧl�����>�(��A�D�-g��]|3ͭǓ2�nX����ݤ{{���^�?�ܗ�3_�����''ۚ�t=����t0߇+Q:-�Q�uy�ǹ�����]K֘�c�Z1L�/m#J�@>(��}���v-�)�R�JJ��a��G0/�x������lġSR	��,�*j'&,(��g�f�7��W��+l�o^����KH�6͔_�W=Xv�\�qzl�o�g|>��� _����,ߧXH,�`��Dg�[�t������+�L%�,�*mּMP�A�a3y�j��5�&}B��O�\c\�ƌ�. ˖��Fb���1������ݰi�Je�zK*S��({q�2�W��pI�l��vf_�~١8)~�2pv�eι*ߤ_��H.���Z�#�m6�D\*+����kpv��z�7�bMH"����ͦ���o��?!ZmN��ɛ���|��o���>D�����/<��WC���6>��A�
�nⵐ8����O��"�Xχ ��c �[�����Mz��}��3ߤ?��S�w��}����-nu�=y���໬�h�B H'N�q��%_4oT�>�cC*n^7��/~ȧ�*I4���}Xԛj���q��,JD�4�Tl���s���G	h��q����5�.DY���qN�lf�q�|�J�4=c:�vU��܋���n�i����A�i����sMJ-_-ϡp��H�RP^C����%�iȓ�qf&�r�Ӄo�A�5�2�����S��X:�,���ϩ)a_$�ryH.f��'D޳�U��x����lUet._�����S-<� )��ԛ(���e����b����Y֓�+h��S˻���$���9JGT��#MJ���}�߄�7�3�M�$;PA�3.�����%В��͚r�0%�>�I;</D>��hk��?���c� �Qe��N��R�5�j��O�Y��0 =H�*a�i���P�1�M��
��KJ��%��ʽU��[y�g��H7��d��<�v#��_��.?��_�!�)��S������5*��t��B(Y�7K�>-@ɤ%M��'�2�N�p�ӓ���k�������=�[�7�m�+Q�x�F�^e<68�>���5,|8q�W[�E�wQ���)<�r�+r��o���^����7�?<�M������$�[��m��!�3`t�*�;8]��uh�3�����r/EZ&�30r�T6>�e:����rR���'��4�`aS�х��!�$��<�5�v���Ȝr����M�o�eY�4��<ZYh�I�{(.��k�056�Ա��������{W|Z�)�3a�k_}_�W�|jTZ�5�,c�̂��A��l�C�M�6�����|�>Z�+��ƿ�<ۗsp���c^;�*v���'�N��J��hs����kV��Cю����<%~�HFlC�!�Ͷ&���Lvј�
l���:�b'ǴE�(�KÇa8z��L�nR@s���7h���^ׯ���sx�'��ѕ��W��_Å">�����pJ��{�������O������?NG���X���|��Bp���Gyפ�d	��H�����n��F0���pGa��������}���ҟ|�Yz��?��Pƍu���I�������w�ϲ_�O��O:%�+���=>Nc#��P²�s�����Q1��ʘ����T�ܢt`_i����Q�8S��.-�\�� �M�彀ڤ0?�|.�K�^�Z�@SٲdЀ�����4&}hڅ���ih�i<�8Qf#�\�}9�>�a9�>ĵ�j�!�:E�X�8˺Ӫ�$;�܃a[�m��p�^��V���c��k;�]��d=�N������	�4�i��h��`��:��&S6�R����8���f)M��%��m����K���8������i���;��b�f����o��n���]px<�7�&�\�ג�SYa`f'!�YIzk�j�^�WI��K&�6H����F�p�8`8M�p(ho�BKqI�PrP1�����>_�ܥ�V�9��o�%K�kI)� �H���,V[�*�@uVh�ej�t�gG))g��Yo���ǜQ�b�W�Mp@'<l���C�q���i�_��<�F�=m�ǿ�p�l��Lj3Af��tU��H.
e�C��:=�e��nB���l�/�����	����I���Mg�����âf�2�s��e���<m�.b���=�DE�׎n���k��+��.��O�%}��o�O��߹I7�E�!6#E��t|m/bv�m���<'�<eZSC"_�->����S��P��rY^d�g��8J��?������>Mv4�j�5�ڧ���CӼ��C�ެ����|�\�1=L��p<�}\-��[�ߢ6p�����q����q��5p;�CZ���<��z��K�d25�q����|GӸC҇�3y��K]��$���+����wy��r��	�P�V�r~A/������\��6��ϑW.��d!H�7j	m�=A��>n0�a��y���J�����ot�HG�o]��iZ�t�������G.�~���Ҝg(�gS�Ӌ��d&�x�A�I�e3���|��cw����%}�W>L��!�^����'�c��D��y��� ��f�q`F�υ��aBu!�|����l}�{6������K_�?���_�׏Vt��m:z�]Z�lP�!�)^�B#mC G�e!�6`
]s�Ů]l�94�G^� /��>)�U7�R�{+>�8�{�ϗ%gK��R�έ��q4w�����̾ˮ./hi�4/��dʩ�q����d��\�#�V�@�Td��y���e���5z���$?�z����7���4�z��.��̺u>|����Vq��2jR�#)��܃����O�&"��iqt,�8�}��?�L�x�/�A�Ѧ�>]WX[�R3��s�yN�)�1+΀3
�Xi��� }@a�HZǾR2�ӻ��A,9V+r7no��5�����
���QI��co�j-f����o�%|��4�S�X�P焔�v3pԠ}�=44}��'�R)��[�ۅ8�oN���'�R"���~�#.���x`-�;�pU^�DGH�������:'�u�7r#?�3e�G~�pZFmN-��(^��S�%�ÿ��Y�B|Z�1���l4f}H�Ō`��!Θ6Bf8��O�x�E�$��&P������eQg���}���K����t�?�>_��̱~Vr�=_�B��e^Q~��EG�c��)�::e�j�i����?��|�9��g���~���{t��6�c7���x�0�1�cq�(��f˿�X�|SD,B������e����Y�E�h�(��Z�b'�촴Q��
���
(���hWH:��g�"wP�t4��w�����,�D�o��7C�ؾ�����m�j=��#����sp��ٛ��1��E_�v4�ҷ�v��K��AKwJ��4&�(��-�"Д�Ѕ����"�0'�@��i��V'��t������
lC񘳚t�L��8iQ��o�z|��S�ک^�6���!���o p0]ho�L�M̳�=���WF��u��u�u*��D�bVZ)�N�O8ȼ1��pK�۶����_�o����Ane_���G{j�ؓq$ud�`���<��r|E��ί����֞�=$z�?�O���O}��{�'�j����#����޲�~�M��B@:�;Ïn<��yO��'���I	�ؘ.�J�7� -.l�����F�S��W!�y��o��E�9�3u)���1�k�Q0��w��
Kl���ŐS��z� �V�q	��5`ٟ�S8�ik�(��O?�ʔ�$���&i'�����!-3�c�/�G���N�i���|���.]�����̈�Ɂd�?�w�c1�W�{tۋ�D�v�>�h����4�m��9�+������(�]8��#�����v��)�t~��x<�/��$Iv��s�,�<s��S/��DK����B�#t\t8��=͝���^�ʛ5Y�$'��s?��--~	���ECg�>���Kib}:x��.T��zv��q�����"�5����=���dRV���*X�!�rYre��y� �Gv�?��"�m{�[W�	�L��P�ᴌC��t`��f��@<>M���O�9�$$�=NUJ�7�St_i��L��S𑽸)WB�!�8�v�w8`�o��q=��o}�������@s.��̰1�%釁o|�|Cl��z���<���=���O���L����o��=\���7���ZuÑ��azi�%��;�Wi&��(���]�^�����r�f����r�f���{�a:'�ޢ����N��7lg$�HC�k��)i����c#N�d�~K�G�w]|��@?ꭱ�(˰�E;(�N0>�w�w�['�P����l�&�N����c�@xZ4�ʜ�)�,+_�7�֢ł*oi&�A���D}����m��0��ϣi �F��b���g�u��sO̟\��:יNꀲq�]o�?rp5�p���XiGޗ��B�4��	��~|���H��<�d��~L�Y�ɹGk��K��|�9˓�b
�'�Y��T
�v�{��V��x<h������`X�al�;�b3��v~`ݥ�p�ɶ�x�e��/~���Oї��}����tt�6�x��n=�����c0�[E}��G=?���i��
�D�S��R�i�������������t!�{ ��M�b?��I�`��A��~�O�=7�v�5���L��1�
{~&}B,=�T�uxm���|�ǳ\��3�i�C���#�]������+iw�}�]��V�R��v>L�<��ҕ��%�:^��
���!!Ӛ��G��m���zჿk�i�f��g�3f�i(��m;����\�I{��/�q�t�;�&�.
��V�V�L�8o�v�tH��W��P'~�6mA Q
��ʱ�Jx����0�>1�O�w|4��E9�z���{V۾y�z:van��-�o1����0�٘.�5|��>�6��CN�Y���-�yq)r�<L�."���Od��P,�����$PY8��ab�VIK�>���e��
V�p���e겵���"��9���S�9f*�����$皧2#����|��[�k��[���c�}�eu��J@���.�����FG��*�b��V����ָ��N��Y�gØ�	�:��"qڸ��N���B(����Mme��R�[�΀���8F���o�ݿ�8}��ek(<���Ć�(E��eۥ�ԁR����Ѥ��h|��|�w��U����A��s_�/}���m����t����
N���G�;g���TW7Fs�[�"��0��b�e�������i*l�8�:M	K�3J�ӵ�/wq��e+;���$߃=樐�(SC��K.��l��#q~&���pE�d��cP�o����ԿX�#
��e����Oql�ܧ<c�D.��yI�KC֠�Su�m�<���p$|���?Z��e!-�g⸬E4(�k�k��3�`/W�|,K�Z}o���E��U�O&S~�{�^g�<�D��-�,=�0?����o9��C�y#�Ҟ�a�L�=��+�VN��(5�zV��Oy�@��`�����A���<*�"Σ0�K�G鸟}1O���qi��!�e�n+�Ԗ3�0�"�H)�8ȝ(��p
����o�����=��|���p��x���׍�^��1c�z�"%D������}���_���/ӟ~�)����ã��ܡ'�n��*����4��.�G�w<�0^��E��֋�B��N�ჸG@�q�g�_^�ʽ�e7�m�D�S+�>>���1�إ�in�;��������n�������=��h�k>�T'�,(%K*5ُ�a�:o.���E�l"��C4 �;W�O�ZP[�_RV�������J]-A�9}�$ь|��W��<r���"�'�|1uF�W(�hQ��lU�7��|��o�:mJ".������}l���u]
��fX����a��e=_�=��O:p�a�?h�]bD��_p����
a���o��g��.��b`=��-B>�0'=7J��@�N��DGǣ����=�1��X�$XA�fxr�tPz�]8VBT6�~�f!��{�,�8����XoJ�R��J�a=��kў|d�i���A�~p~mU�SMmA�W*�Si�g�8�+��H��i��ۚ��H�����O� ��>G��A���*D}ժ���Z��N|Nt�4śx����A�
)�!�7�=͍,�p�h����0��l�S8JXd��ђ)ӒsV�b�I������8c���A��'��[��$��A���
$*�H���
���5���a�tH3`�m�5���o�g��u�����ͷ�K�mB���xEG�m�����:?���?J]v@/��1LNt�C��5P���"� �+s�R��w�a*�������6�ҭ�iT��~�W�X��N�-��+�=�+��hGsW�K��XJ���n� 	�h��ލw�c�Ǯ������]�Y��n���iFYS6t,V~Z8��F��"�f�7����7�fK�j���`�9o�O
�uZ���f-�>�=Q�+�C<f����5��Ӣ��y.�!'�]���mC`.U��.W�+�8c0��2W�뒶���v�¡������]\_�4�x^{-��k�w�i�0Z�>�N:`�R��p~���@��Q-�A���p1�uF.�R����/��};m��pMI�[���O~s���:�HAß���e����f���kz��ߣ?�ܗ��}�Wh3аͻ�s��É����!эB {
�w9���������:sO��n1�z�t:�?˪ӳ8�З��^�=�s��KtX��n�uM6˕�%v�u�ݥ� ������~���j���8�c:�->�N���oq�[�@u��8��,hQ�i�\���L^-_�7��hо�S����|峖� '4��,|�GR|�ن�-��O>'���AT�J�M�^����Q�d�ȧ7�3�#q�I"��A.!�*���S�4��CZ}2�E�]��8ƾ��ǅ6ܮ���Ы	� L�h���r������;��ߺ5��À6EF�d�Q�g4˕:H���8�p��Yֲ�QV�V�	��=�Obx̧+YU��Ƃ���f"�S7ȏ)ä�Ke�-�.�R�n�V3f��
��8���?��{1&�6%��Kd�7&� ����U^]'p�0\N�漻���t�o�T��r3f������u*�Y��V�R��M�p�ǀ	G�����dED��!��"�ǵFW���E=�Q�������W��}��_��~�z�g�уm]������1��A-c�Ȋ���2��821ߦ��驄��b��d>�"�,��n�>7�7,R"Me�څalN	���MR�n�t ��}��Y�:|��,�V_�ap"����~���5\�"�&��}��Y�>¾Т�"s��*���U_���}GS�=�W����w���ѓ�ry���#r���zr�V�L���>����!�|��Ot�Z�	�mă��>�Eyr�5R���.Nz��2c�3�<̑��8����2�Bi>����'i	�%
^jSo�)7Vk�;8� ��I�c���Pؐ���ؗa��=�y��ì�wr����S��g�O���/��''�nݢ�o��[}<Yٍo���j�{R`�!��c?ǹ�"���n^ʛ�n��H�Uf���ة�qe`���[����+��B^{��EM�s�l͋����KL�	<7އ�x��쯻P����b���@���X�[К�5�؋�g�^��1ʴh�kaj݉��*i���g���l�3��p������tQ��Z{0B�Ē�� C�"� L�
"�G���l�xJA����P��.��;o*0U-�N0����������p�7��e'p82niiW�ɦ��z��ul�ͱ��b���*zi��BaPC�.֟#����6`��<	����m:9>�~s2ăc�x�.��+������h��vM�!0�YƇ(N�P��]���Me-ɹц 
�^�K+)M�}�ȇ_
>x��U�.Ӥ����e��ў8����j�U&>�ТEl/�����PlCM� �2���A��ocY�Ѽ:�ڑ=$;��r�uA �+J�9�J2��f8eƁ�@��=p���QO%B�%�~y�(]�hgl�ɖ��ܮ���>�����~Q�	o�� %��1���V���7��������oҿ��W���!��������Һ�����yB�x<0e��y��bQ�
2
E{�n��}��~��q��U��Dy�(Em�7͔3� X�Jr)e�ʺG=Sq�ĉt�����y�iޝ&�t� f���p�@[��Gk��T��y�[d��Kq��S4��M�`�u��[�o��Ή>�[@ׅ2
]�t=�b��>K� �����$�Q���CN����\m	x�X��Z봀�}<(8���c�K�O��'���O)0p�%VN���"H�C���	�qR\��:�ș�9�q��>�<}B���~�Z�ˆ���a ���b�ρ+GW���׿���W��?������J��cr�kZߺA���?	o�!H=`�1����q��(ǌ�|}�J�y<�]��3�d$���� �j�k�*%�W� ~�ɳPEZ�E((,u�;���חe��aܔ��X�����11ה)��d#ڸ%s��0vY�~��������|�S�D�/iA{�Ȯ�z^��nG��}]�e�ު|H�ୂZ}s論�� $��f
��G0QaH�I�VA�(��8��d���NH�z���ߐ��E���HHc��[��6�)юu��I��m����EC�F#�&n"{�^��uc�C���&���6h�����bL�Ǉ;<�t�����x�e��>��ѐ�:�}:Y��=�$=��~<2�e�$��G�Ю�
���B�Z��d'�N3^+3�,��)�6,�$�����JJ?��T}�14�A^Q�U�}�V���?�ph�3���8j<��&p��g1�Y�۞��i���K�k{� ��%#�r�x�[���]��M!�Y����%��p��e��W�p�cם�=&E�������%�DOݻ�y���#�z<f>��\L�<K}�ǃ<�ARٸdE!��//d��?<�j�Mn_N�4� �A����������=����׈���1��6+�.|��c;7A����ܾ�ßП}�)������Bo���:z�&��&Ի��p�sx�̅Hhp|:\��ldg�Ot'ȥ�y��	o�梯�1�|X�-�g��DI�+�pl����g_�m�$cpq@��,ref�Mj�:�+�s��i G�9-�U?�և�d�=��Ȭ����.OZޙ�5͗{���.ֳ�6���V���s�I�+�$)�6�[�#X4X����eM��O�E��|U\���E��G�y�k�l������.}�(����Zȴx	*T�u�IүI��Z��9��E;���e0�)Zֆ�^,]ȳ�k�����b~���K�*V�� �ڠ���!��j^`�ڤA¶�5%�G�K�Zf3�;%�_�21����_b�1�Y�é����_�����w��pMc��1<����x��p���9�oK�p�:z��}��3ߡO~���S_�}���wn�z���;�i]�X�����2�n�l���ځ�ܒrF|�*Xz�O�6�m�J���B`�kL�M	z�6���@�9E�l��Ȥ�X$eN-U[�8�Ƽ�AF۷�Y��ظ�s���P	��R+�/�3�*8�!O�����&��A�-P_e�m^��20٭��w�Y���{tY�ڿ�y
?b&}�?"�F���"m.�'=�g�%۱�_�kg�#l.����G�\��sVzF��I_K����.���˼��O]Q���d��Yw�X�需׆8��'pL�� OKN�I�����& �#|{�Y/�7ZG�$�,Iݒ,���G��	�a�ph�њ�w�҃��HN
�4��eD��QY�c��&*��<Nc�$t3}]�~�"�H���â���tsh�C��C�'���o��si���ʤ�8+���R�l�:�?�PAAB��D��~͉�F�R��	�>,�k�g-seHm�E�UpB�[Dٰ;�69J���i1|W�|P1���N�st�w/�l�ˤ6��IZ<���^ԕ�Qٟ��4�\@3��?�8$�֗t���ֈx�dC��ӟ���������16$q�qs���Z9zp���/��>��g�S_�:=�Ы�����w�F�
�õo��Xݰ��APlc�y�v�?,�|����������vO�dj�Ycא{F}Nwjn
M��j�^U��M�B@{�ʩ�H�E��6+ k.��d�ϩͺ��>�h{������k@��˓��pk�*s	����Z>)�o�h\Z�O�������X��Kӏ�D;��!���U)���;.��\�'�7�=B�eZr�n��.K�z�!���n�������D��p9�6	l�Z��/��s9��.�L�C�1��Cc!�%_q��(~���4����o;�C�FD9"[�
�}��s��~�7~�2���|�����1k�G[_�H!�c���K.�G�xz��oޣ���<��_�:�����?�)��&�o��ɛۤ�q]v(n=�u��(f��(�˭Gy�߃�E�Gq!�Y��f�9w�(�4�kQʲ�J�E�!��\5��"_�9V*��0֋�"�bph��k}p�t�y �[!s\�僡��hSg��"�{1`�i���s=�L��*�2YN	�h'��Q^���P�Xe������ғz��o��Vו	���e̘���Q8�k����D@Md?��:J+�N��̧�Vن��?�<����x=�֎N-�����>ژ���P�!x֋S�� }l�zLn�E�e_Ow֠}�t����� �HD���tIl��E��Mt�`�y��ᴍ>���c4vO����9�Et��p�J�5�u�i�W�A����:�ɾ !�ͤhD+��GmYn��e�����z>�|N��h�iڅ�S�	�S���I�6���4���2[횃�`n1��ГV���N�����X����I�O�J[iR����C>���s�9q���y��!	����9��3��4�P�R\D_Nl^�B&�t:a��p�|�M~"�.����EH���8�������?���_��������;��d�7q�x�h�����'���/��}���+��_�z��{[��V�q�7o�z�e�3n;?�q1�#��%���v$�����:'لb��<�0�Z|_Rϼ����z���߲���\�ϵwFZшV�s�p%���u��(�i���ѓ,��	[��;����k��`I��}N�o"G�(��[@��0JT/k6���KeZ�m�N���Y��S���j�[����!�tqZ��C�@W�m�Á!N�D�� C�d�^�q������v�����6����-pEr�������s_���'�b,��1���8N'�d�=�}8y<��K�'	�҉pΦ��_���lG��9�I���k�4^'='����aS��K���}�t������t4��C�U�|��������ӷ^���W�N�����O^�WNzZ���k�M:��i�O�>o4{�ј�(�طI�6��z6���/�E�/?�[a���#�]O�E�<�����:��\	5�|��Jn�{s��lp��<���k�|P�.�'���$��zY��TY�1�6�4tUh�Ƨ_J?��S��k6`�S���bZ���f<���G��2�Gs��>'�4W�19��?�Q8=�|��D��F�|���
�z��o��[y���s(PGz�������<���Ӳ��"���8x�	�X
�TOÝj�h�х֓K`Q ��r�?�U��Н�q2�'/�_ �xy�}~��91� ���\w�ύ[��[�J�ܢ΅�
�S��G���4��$�Do��S���`��`5p8*}%_'�G�w����z�p����N���?�<r�,?�v����[�����E%-�yj��� Je��ʅ�|�|�3�xm���`�/��`�#d-Y 
8��ӂsG f<��*�u	쭃�I���T��c]��}�O��9D�/~g=omN@M�0�s�f�.�dY4.���ܯ==\ߥ?~�������?��'�7>�Q�}�6��pC/��}�����>�4}��/���!���;>�ۏ?N�9�}���~�H���W��	�S	@��|��~�S��A$�MU����JoISp9��7�]u��r��`	TA�AL^��.�T�����j�9�ӧO�e�m8���#v����e��_����8dz���xTb�G�p�poV�]O�^��p��
��z�AJ�"���i{p�>��F��.�4pM��B;�C��Y���.ԭsykҮh(�E�u�#Uf ��%��yd*�ݫl{A��������~(^���Ig���?�k���o*3�bJ��x2o|8 Ǹ/�J�+GPP8�sA7��so�<\����>������Ixfo�s~����<(�)�m���;C��#zy}����$=��s���1z�/���zM?��}��/�_|�K��o}��{�ez}�-wR�u���r�G��i |%$���O��:��g����W6��L.ia�VC�_ڣBʶ�ʨ�}�2.T��͒�t�,^���L:���>�� O�z��~P���{�.�&/�)�q� WL`+}� 0}DM	8��\�ߢ�dA#W���D�ꓤ�P~V�U������%����3B�d����z�'N'G��zW�My�_�\쿹l3q�l/��x+ZI@;N>N���*<����p>�.�:@�n�b+�� ?�H8�U�~r���_�>d�oL`�ͥ��0 ����O)�ca��M���'�u&�|�C��jM����1
�����`w;�C�u�Bp~�w�h]b���B�R��w'���
��iEG�|����g�����,\��4$�pS�F�Z0��*N���S��,�W8�ʨ����P������`���Zx��Q��,� ��||D���c���.�s����$Α��_�'\���� 7��
�4�)`�;��^}w�t�#(̲��Ϭ���ٻ��r�(�MG''=��Xѿ������׿�_|�.=����o��N�6�6��h�o}��N��Z"����l0�]��j�H���S�����`�2���h���y�Т�-���D[���t��E�e��ͫ�l53�Vs��\���BN�Gv�Ŕ��{x9��i�s�n�7�MC�a��l�ݜѻ+�`�͟G�r1}N�H�X��!�\�5K��o�Tp�L����9W�W�S�Q��T�|���A_�]�Π}}-��J{�>�pԠ�v�-�)I���|��5��q��z=��/�����tN� l�
�c���9R����/�fe4 �56m�.>���~׳)`�������e�F��(�y���y���kp�	��O�:0z� `;�A�X�p�j�m�Wv8Zm}��oh��~�p�}zza����S�������=9&~��酟�I�v�j��n/�s�p����l��U������[�(ϗ����A)����S6�쐜-�����\Ks�+��(_�柕�8=���joÂ9���s�.�F&�e��$���G/�#��p�e��e�h[L/*$5Y�-���|陞�T��3!�*�i�Z���~J�X�k�(O�O�pe����\���x���~2�ſ�x������WhGP�I�((��Ǔ��~Qv|���\�Ø*����Yz���C��0c��>?X����p�n�Vu�=�Ei�Ԩ��S���h?�jπ�W��\8S���}�vz���}6V�׊��X4��<3Q\�>���Ԩ1w��G�tw�{�-״�'c���F0|G�=n��d3w�9���}85�Y��x�P�F��Tn������ɅR#��G��O�>]�кK��B�/l�6�]B	�ҟ�h4yECa����!U�l�B"S����v3<-��BȨp���nWa�$���J/H9��#E�4/��p8�8R:�噋�W��؁Ԛ�A=��CKXQ�Uv�r�S͞8F��@�;�r�mT9��Z_��О����hOt��t��=��5��;zv�N~�҈s7���*���>g7~� ��G�%.�F{#��8���Lj��M+jL5�Gy�#Z �i>׸�C��9�e]�*��A5�����LüQ?n`7�tt�l��E/�7�����N��{�aJ�mr���`���S`���*Sv��Ǽ�	��������2®cp�77����[�G'�eY d���lW��������Up��C�Z�A�"�L��oAC��Ns��C��O��)I��9�(1]�`7���3��K]�Ki�����8��s��kg�m�����O::\����w�iR>��%f�%��	�Po���x�;@`���x���'���6�y����e���\? ��I-Qg�o�]��stH�6��jkg�������ً?{e\[������p$�)�C���n���r����$_uIq���I�A� �'h~��	��׶�k��2����T58��@�&?������
A��S�,K�q�N�E�d�� F$��p��x�9��v�.�Pp��Ƃ��ȟ��Qcw�Xv�}��k�0������U>��C0����k;-1-�ծ�lg����^8lW!��[�E�Bӥ�h�v���h��90S�g=�w����8k���J�f�	�d`S,��´�;]�����ϐ?I)Z������`������њ�p��+;th��c�6�Z}�F��B�]Wi������5��["�C�3��q��zi�견�8J���Íd���c��bZj?��\Z���[�×8H����e��1����<�zx|D�!m�/;-$GڒTsd8N�<�˗���3<��!�$
���BA)Fx�e�ά��
.��t4�3k\&�6fT�x���|���.Ꙡ�^�'x4��f=3qKy��w�f_���+��Ɖl$/i�q�geDc��S$��OL�L4'T���
ʌ�x5�/>��E��@���W��i�
��~r�Ft���	�6x֦7�"�=��bo$.��YR���j%�[;X�n��h���6���͐�v�9��͑�IǛ1�)��1�#7e(?	<n}�r.��p�e�ckCMZ��w*E��R0[ i��W�Xd�d��<����3�uZ��.�Z"�MEQ���I��R���8�9(���;M��1�x�¼;]�p�����?g��"�R�I��!%�ه��>vg،r�on���|.�4M;�}ڵ�O�>��,�-�)�>jmM�B��B;�W���Q^�o��e+�	��q�#�	��|+'����Yno�>���l�L��?�p���a��p��'^����m,���G8�P���(��"�B�]|n� {qO�~
�w��¶W���!�+�Z����S�Y������nݍ���-.nu!O�V�z?^����y>���Ax�x�b4���G���E�z��]͟Vz�g�S�S�5G�'v��J�,Қ������d&���@j$�����NP�����*W��	|ɬ؟'���̀K�ڮC���Eg��F�T��Ս���J�P��$�$N���H�@�U�A�hG�M]��a>^��C��ܯjѧ���ʦ'�w.�����LW�ݗ��JzF����+�?�3�H�X�V���ڊ�V�A�TZs������F���d����/An�W�u[[l���]=�]���/N�i-��w/8mU��qv�����ׂp\|`ǅo��z\1Q(�'�,"����1����x�z~�b������x'���?�7G����=�CU
�]�`� n"�SG1A@�#���^�қ8��e��V-�gFV���6��ٸ"/*C�}V�Z���mxh�YV���_����4��=,>8P;����R�㛀�|���o����@i/�~���T{�K&׮&�qL��&��9����^�����q�E:m{�9��tdɓ�%�.��)Q=J��h#�E�8)�c`���t�����1�����m{6n��aE~�h�H\0���6p�����W>-����1ތ�Y��:[�R�(KR��6�}�*�7�b�'�y�
�s�V y�>���񒙜)%����X!��(q�8P�e?8m�r@-X���]DA럶Cy���^��u>���=��"D�K�M㜪��,Q8��-\�]��ͤ��#��E{�[��Q�>j�6�W�4���R-&o�?J8��#�9[�x͔dg�`����:�P>�����M��7��Rc��.'L�����޹�\��ज�EW�y��똣}\عJ���,c�xf�����P��e������8ǧ�A��1�ʅ���x)�*����0�я�²��%�q�Lqu���D9ۉ��$:_���|�<Ѭ�eA�(���B��^�]�Σq6��x�|�:��G�:���.I�����t!��V��RL�=:��X�ル���4���(/��3�)S��ƳE{*���L���6h�ŧ�y��X�`=Z�X4X8--���3�e���A��Z8�8%�qO[�i���^�g�s�z���0���r=�^��/m*@Y�$t��\�[�ԑO͎�0��Y���#rG7Ơ_��m�U�!\h�'׶�NZf��J��c�I��ͅ��J������i��%c�C4�Q��s�=݇��-�\oZ�e�MO�������^��¦w���������s��L�d�;�C��Y��&/��Vvڿ��PR,��82p���&uJ�y���s
�i���j+����jW�>md�)޺��`R��#�(S�A���T�@i��?�U1o��CE������L�ƥ;�Iӗ���R	����j��_M]\����(
vY_\D���E�5qT��<I�i;���X�ɤ
<��3-y��M��`#yvg�_n�T�'�1����3�\�7N�)Ûg���k��p�&>��	\�!���M x��S�f���z��gi^���9�(�l�A.O����1�VYH:�[FR6�fg%n�P'���E�V���c:�Y��
[���ϳ�9�9�p� ���WW_5���r�>�m�Do�j�BE�åz2�7h��;��hL�>��hߟbEkoi�A_�c3B�;�v��s�-�	�0�Bv=�)�U�N��$m��#֗�<�`�M�33��j����O���Q��z C�>��8)q��\uދ���X�\���Yþ��%^	 �e�#�cJ�����RD�T'_�褔�s�״��(@�w��\� .�[v���t^���A�M$L0��X㈉w�'�8�7��)
�!9�s���=TIB�S_Չ�N7ét�󥐥ҭ�j%Nɼ)�\���I�sʺ� �����.��A_C�����K�n=^
�|�Bef|�'�m�Z���3���
��Q�2�*�͠���r2���Z�����^e�&�!�����?_)KWS-�qH;�h��1�����O�U�c^�{0��8��b��������x�ZRt��_@?�8|%>ڽN�8:��ܴ1�6_�M�+�t5�,��6bJ���Qf��N�覃�4,
��2���S6�`]�R�_ha8M!��w�7;�o���^�o�n-�q OcD�f�l��z�.��l��w�����mV܄��9|��k<���T�9�Iy�i3cfMP/[���^T~�9�!�e��������o���8��iP)�v	���E�
v'�� �l��e�ﭾ�V�E��pF�YO;�;i�4hv2*e�Y��<�n�oX���Թ����1.��phȲ.gAI���I(�u�
ε�4�,�~H;��Q�F�˴�Ie;��a�2긐����
B:+��6_�Jf�(.8|��2"�v����8�6J8"���{Z�u~�s˝��#�1}����'�ԉu�[�oR=��T6��B!Ca���h~�[;�sKқ�W<F`|X���ݡ;��6A��%��X�%5�t^Gi����v��уCm�֠��,ƅɇ6��8?��g-\�?��>�K�����ǣ]�%h��eYn�,ڑ���i��
������n$(�L?GW�4B�:�T��q����r�w.XZ��w+ߩɍPx��v���s���}�/�a�2�/h��L6d��"�}���+_ �f��TD��O����M����)Uv�K�c-.˖��L�/ĥ��e��� 4T1�ĥ6m���k&E���/.\�+����'~c��2r��I/�x|�%d��q!mP<�)V���j���$}=��V	�YzHc��.d��5,@~���W����U�\�t�_��A,-~I���+�q�E���sp�y.�F�,���.pjN�|^%�E���I����S�<��*��A���O�"��
Z���
o'qs�pL�TAZkp&��Q���zCs8��gIX�ɸ��!��z<�ɧ�ut��e܃��|٥��փ}:�o������z��(h��f�њ�.��u����sr"���b���٠�>mg�V~>Ac��	3;[�	V~ٹ����:����������_"�6��ݦ��1�r�0��1�v��iGT�iT�A�:Ns1:R���&�fL6�e�~GJh�U����7�㖥�7�d\���)����xq��Wp�|ZA3ogѧx��h%�">�q}5Z /�`Z�0J��P�,Pn@2*]�b�&��I������g��[Rw�t):ث��7�ذq���A��=!��S`���T&Зa.��N�������.��,#Nw�<��bNR^P4x�e�$����]��z��o��>H��8�T����~7ܲ]��/[BA�[����ysBPk��sV8�M��<�d�M)�3�������O��j="�5VH��١{�0YvS��Rj�aQFeQ����r|�b1U/�q���{�A�����I:����g$� l�N�Sa3�8~�� m�[��]ͤ��iT=s�┨5io�Giw*��~}*��é�ƌ�J\ǥ��<ֲ_�SƼn��������b(�<~	z?]�zw�z�v���F^Y��{q�,�����~��N��s씃��O�<a�q��Ҳ�k�:�`�q�#�?�"��,��)ln50������|�I��fcZ�p+�hԔ�"}ٮ�u���2Wia[���,K�9�O@�Y��"u�,A������5Y���R�4�D�1R��-�+I���q|���x��1��},,O����˹� YG�'�_i��H��?����(�g��K`����*�q�
�]���[8��2U�-\�L	�c�~8.��*��n�X^�'[�Q��7�>�]��$�;Ez/�%��팄�}�}���-�)�j&��<<_�b��E�C��ׅ���a�L��~�s�U�~+�����A/vi::�էn����n�x"`���k��KdQwSL�V�s�鏸���ƴ=�	U�n��~���i��`�@�S� tjKͥ��h$46Ĳ�5�W�C���'MPn8�9��j�y�����J�o�7��h=�u���096=�!���o����3 ��]v��٥$���Ђ��	f�SP���	\��N�c��#���]5\Rr�i�G�,�L�E��i�>�_�G�^�	p�}b�K��19�'W�6
��齎;Tȷ�T3D=JK�⦞�L&��6.�.8K��Gh���(�����Bn�?.y�/�~�#}��׾U@F,;��:�<��>l�<��%E����� Mn��1��P���S.�m�V �XMɹ��7�m�U��ZbI���? 	�V�v��i��X���>�r�|��v���j��6ZlTMw������P�eg�I��[�邌���Nฆ����66��{�,q���;/�.3�s�3q�X��
��I�}H���6��%l�P�O��.�K���{h{E{N��l3e�l�.�Ǧ\҉�ث �=�X���x��3xa�kP�Ƨ�������1�G{Z���A�F�oSm��j��pPz�B��l��O/��@>�q�rT[���������rBh`(ͪ�f���e�������>���TD\�O��*prIZӚ�J5���3��2c[#��Q�vՅh������g��NM����<��} �d�WD���Z {Ϛ�!�΁�lISbF�)�B���J*�Y83��=6�B�)��(S�ԜU�I�$o�v7x䠬B}k�iX��xeiʩ1c���\Ɇ�H�/x� �$�Uk��x�z8~` 2٣�r����X�N��֨ٿ ZݾM'�#�M�g��C0��M'�0A��{�]�U���KN�8�ZE=�����1��p�X����g+����H�����n�6
ic'�0v�~C'7���������{�h�>��A�nhu��ë΃�1=K0��=�<jӬ��F
+?��A�(��P�^����rD������U����f[8�]3i[m6hp*��.M��.��M���mA�n����_�io?�sƳl!�C�b�a慐h� o�L���Z��$K(H��p9�� S.���t�L��9�q'H^T�<�����x�Ǚ�dG'��֞.F���Y��&�ϥ����ی�iJ�c���F�p�r���q�$��$%�Nc��(�
��?�o|+��<G��'�ת(�M����J�r��J�IR-�62����yK�a=5yp� {�f���-f��ʃ��wF,z_q~Nd�<�q��|dדq���������E3۵;���ay;��4c̐A�k��6�,�I��8��ϑ�FQz�ǩ��Z>~%Z
H<ɳ/��5`��E����E�.:`�~˞��O?�ɗ&���<&*b#⺜�Ps\U"��S���]����i�0�ۍ^��c��XKLߢ[&ۂ6�.E?��I�5�˷x3O�����,>���a�-�\���m�½��=t�N}.�Ӗa���G��i��#iܐvb���e�u��r��@�β�L�A1�]~>ʌصɦČ��\��L��	�gѬ뛳�4�Z�²,�7�y[�G�߉>�$��Q�v��7pE��@���Wi�xF���0/�G_B:4�X�v��S�b$6HR���	���t��P�+��ZS�E����-��<�Qq����}��c��o��Ii�9�u��(�h�-�h.f����5�r���~^��� ��!�j]��;=%W;��ߊ��gV�h\��r>�m�ù0}8���n�B�|���=�����J+7�����6.&�5n��s�~=� PHwʿ]����Q�P4��*?W���g�K�9I�o��g
�S8P8�� �z4�,���[ksj�S�����{�T�|�����%��+��8��#��
nv�?��b���s�DZ�$6�fY�����jP���1O~9T�B	������h$�.p���ל�7N�pe�]k�hA"�����<p��f�@�:$��cxq�6�aЄ�� )K	��_�)���S�}B T�-7��'�DaD��k���i>� rBU�fJf�ְX`4�a�%� 9��3C^0Y%~�;���vƸ�e����~"�-�Ns�]f[��_]�X�*�o�+�E��{Yun��v �0���3��p
��� ��{�UAd�&�IL��q�䧜F�)�Z1k�8�|����_�QF��$G��P~�����.Q�����|���;X9�Dp��.J<�C���[��F������>~ ��F����v�E����r��$�F���,Jm����TO�K�
��WeB�s%��|�+�@G�VpR�&�ڽ>8�7�|�m�e���F5�eE��<���R'��~��fߗ�-R��f)� xUU�:#�g#O�<SX��|zM��J��iR�2�����j\�ۣ���^�T���pA�M�Ԍ�d�)�Q$+�c�5k�r&�|&��+0BV��jϫdhjuSX�9M1�m�h@��P��D�ʣR�N�kv3�X{V��uR�e�_Np��:'������?����+4�e"n�-�!&�Mt�$c徕D��k���g�i�YO�/g+ho�Ck��l�\�vձk���f�v/�ö� �K�Ϥ}����<���z��x��2��.o���� ���9���y���>V�e%��O�D�Һt��i�f8���}���1��v��".�˧�nШ����A��w��2ڎ��<�wb/�W~�X��>�D�tǢ ���3��6w���5*��b�7�R׃"B(�!�a=L��Qy��`�����n}����c�'�Pڰб� ���d!3��,���RL���|�V�8WƩ[�UҶZ歮%G���HtG��:�n�����R�B���B�+%������@g�g�C��L�9��l�.�T�M���AQ���lt����ě0��49Y��`�K,̳l\�#�iK��H�c`��<�n��a���/	��ޞ��*�E�y3����=1��9P�!Pֱ:�4��u>,�k��o�#��8�{r�I��/i�&���P����T.��	S�Ʈ��G���E�Qn�7x�,�YX��8�]zZ�b	\HWd�d%��:�� ���.]�,��°c$�_b~��&�H��$��T���[S���q�؇��.�K�o�֯����v��R��c������\����o�Y�5\h��wl����-ƋG�wL+aUO��$���I��W'�A�����Z��4�6f;ا�E��ծ�L0�l3ױ�_������ ���േDK�]�:ы4�����uF���q�b�E�M�>-�y�'�Xًgj<�q�-��ę�o���9�P�b��2?�|Y��Zϲ6c��ut-]=����q�t�cX��p����A��i�n<-�� lڽ��f��Q�.�/�>!rdc�l��(��X�Ojt��=��6����툋y=&��@���?ּ�d����'��ƛ0�^[�2]�ߠ�r�lk�D�x�e��� I�H��!����E������2��\垵��"c��e��k־®u]I�ӛDg�/dB|NѮ)'�x�������L�m����$��%�s���z��B�eq>��j��8��kL|�_�,�Ў��(K���T�����)4��SF�C�&iWm��b�A���x[�91f�S��ߋ0-�NK��A vSd�O&�F��pH�H�pY�	T�Z!O�C˧8���(c�Z����������~|���Ƿ�^
��w2�鐏��ܖ��G_b�3��/w�l�t�q8 ��TX�Vs�2|���9��;�ؠY l
�_���$;\���5�W�c�Sxւ�^|���A�1/��p�ግ�;_������?9^���o�h�/�V�7��&�3d�D��{���P(<P<�2,�?�2��3�(*Q���u
��{���
��v5�Aԧ�|��E��\A�������K�[��G����������9Ht1]��X�(�y��&'�
�#x����-
�&�"�\�yT�V��pi��13�|�sY|XV�qy��Vx��4���R�k�΅8�3)V(ګ�B����B�k�-�V"����W���r��y�-2��t��vE�j{,e[aA�<)LY��h68�iAF�J�j�+qD�fqydly1�<i�;#��eeި�[��"Z�.�MEw�c��V`̣l����w�Pl��)�\(_w�c� |8Jx]-|Of�9O��4���Q0��_�{��8O>��^/��"TĮ�0 0�d|eQ�ӕ���o~;V�av&: F�I ��x^Xک�ǧ}�z�c6Kw�5��� M
�Q�ҩ]�<o׹7��R\��ۨ9�M��]�>�����e<1㇌�/}��E��j���0��g�J�8�ŕ���oY�'P�}2�E�Q&��e	ړ��������"�A;�v��ڴ���S$��n�e� =���A�&'pN}�R��!8%��"����9��K�%Agk�H���Ŀ��@�4P��N2~��^Sw�6�+L���b1��fC�E:���{1��x�͕����V���V�C-F��'d���g�!�c$C؋n!�Nk�Y�鎙n;��w8&p����oz��=���뛎�6
o�D7��&�K�d8������� ��%�
L@��3P�	���u���)��I��2�&�|p4P�#�v����L��
Lc�e��ek!�"-�`F� Ϳ�'N��O'��̀�����>i���\.Zv�p����_'剏�PUt�Os?øƽ{�sr(�Z�5*��|�=�*�F�@�xn�/�.���n�4�ђ����K���(��7s�<l�U�fl��uR�ђ^١�c�B�(o
j�6���
	��������C�5?u��<��$�y*�N΂�f8wj�_϶S��.��m{8��(oFk+�8����]r�̗�e�������5?��!��Ƴ�q��6 �\m� @Yˇ�-�m���<�{:g��S.�fo�L?�[�o�b�K�jM;�w��y8h��l��&,�8��ى�k8;�Q�sQ3��k�t@($'���s7g]] /�T&uk���R��LS#(�u�*yj�͢O�C�"��4��(�(k���|9�d�����i���%�`p-������D�E�fq'��tq ���[����,(���՟��j��J;�M<$�f�����J����{߽7�],{#)�WUQi��q=ے.Ɏ97j,G��Y�0�:�I��8v�p�e�{���ȥ��H��Xn�p��p|��8|�7t��wӭ'�F'������(��>�������!'�E1�Es@�d'�+�S�,�"�g��h'���y'q�ۓ�j+�Q��\9�Z��V>�̠]�Y��}sh�3p~
W�{1�-���:��"
=��D&�4��L!(�����Ʉ����x,
�5]�7�
y{�p�6.}���K���y--�7��.g�@�9#����!2�ӏ��S�����9�#��#�s+)���-�*!� OI%Ћ��J7�
��e�8�~Q�XM�亥�]������,���x<jv����YI*��h�>z�P���h�?��a�x"�A�p�����Q��N��9�a	\�y�l�x-0�)�Ǘ�|OJ|�u�|K>�X+��#+�ȅ7D}Ɗ���|��41.�;�Xud#�0i�>���*�֛�JظFJ�\>���a?²�q�+n�1#P3��㐟'�S�;�F�G�;����P'�6����1��#�9�q��Z�q����q�$3|]�Y��[ƺD+�e8��0�5}\��������XbQkݓ�-VAR}�`�5^ή�L-���A{k�%�H�
�g�7�/�(3��O�kr�h�Kp^�g��U��@�!֩�`0�%�� �/d!
~����ր]Β�h�̓�h9x\C��*��U����Z�*��王���x�A�������m�'���>"�0M�t}����s��*��� t��q(��{���u��v࠶�k�����ɶ/,=rf�����q`�N��.�қ��t���׏�h�Ɇ�ׇ��������GOʅL�Ȇ�M�r!$���p���{�_��>h�\{߹w��r�;���v��vw���1�D�%�$�@<A$P$$x�����E�W^x�%DBd)QL��q�;������}�o�f��U�1jT�˚k����9�^kͺ�U5n5�&2��2`��4W����ԩ�Jr'~2��H#�6wM+ڭ�;~�t�������p�~-�}E��.�P<�G�?�����eBr�\������ ��I\8�4U���yޅB��8�3O��x;���Rk�̀�E�D�4���{?���}s$���T����'\��aZ����r�~��\%3��g�j��
�k9�C0�.�^u(&��C��]���w$����K{�WFG�r�hg�.�����+q��pw��Ѩ�5��CK��@#���mSH�h�=��y�}�,<1@�aD�=�R����Z�.�-W�z�0_Ӵ}X���p�vBGoɇ{�96�}ا�������*�C��u4ʜn�k�������s��T`o\/|Hihfܼۦ����(^R����tv����xR�1�M[^8T��6��D�i�l���ҡ��O��2*�l���� v���t����w�n�D.ys��%@�3聶Ь)d�<�nT�h�:9�D9�$�iwW��D�loҰ�a�X������i�h�K{,>��BdS���!����q�8��tI��پ�`6�k~�Z�jM�A,F�N�EX�-)>`�-:py�aF�D� �=�jw]ג���d����on��� ҅��$�"
$=C1��l1H�#��p)�ki䓝qH���o��� ���Y�p�������������o�I���+��rM; j�D|�r�W�[h����n���ċ��̃�F����\s�kQ G^
>u$Olg�bH����� �,��8U�;~�����g#��9;N�������z<Mw8�{�Ǿ�^������fˋ=uG��=�^;��.���P���p�W���o��Fq�	�r��tR�2�]u�"8��y4o�g.@ģHcaiT+��p�7��(���Fc�ie�b>���>Ϣ;Z�X�C�K�H���Ԝ���o�y�ח��^���XG*O�����됋r�؇n�f*�����(\��(����(�����}T �X����м9>�`V�Ӓd~c(��ұ����XI����WS8�z�!��*�G��i�ZӶ�qZ���Dxۆ=룎�·�ϵI�p�ֲXu��O�Ʃ�x ����nA=k�z!QNէ�*^��k}���޻�+���hzb������V�1��	.1�a+����ֆE����F��k����<���|0�!����9�w3��1�s�s��A@����v��%��	���?);=���5��������)N�z��I��Y��)�5��yY����\!g����j�9��m8��Y��ӸN�԰�漮���o���R�kf��S��������<,�,��e.GX�;��I���#XS���dߐZ�w������w<�
R���V�/�`�)���Y�:�Y?���j'坃����g�~i&��k�Z�%�V���H�n��p7p�D]����a(�c�Sq���NLQ����M"�]��u�??�-���!%̘O����?w�_'��G��w��ܮ;fQ ]��x�{�I��~��J��e��}S)�ii��Q��t��q��Ӱ�w\�ZX+g����`����6ȓa(;:�)\�-Ɠ>t����-�t�n�����_�o���1a?�S�+3>D*��,��Z�S�ъx��9��N���q���gJ���X��3�F�ӌ�-��4d(D �$~~&�\D��g���JK��tOr]�ki���ϲ}��΢~���|癏�z@��
L�s�����2���F6#9lxC�eLGk�*<4����ۨ�w��kcA�F�R�(�ޥ�R���>�����ؖ��rՔs+,�R��c���B%�z�d]�˗�E��6m빀�4���w���g���Y;�?�{�#���	�Ty'O�ǿ�Xv�'�x����SʍH􍴉��5bg�'Vl�X�%ܗ�l���<w0X��=9_Q������6�������nO0��ڔ����=Q�3���UZ5wj�%�$���¾�Z�*���;�)�oE����+�muF���6޾!�`�'pr���E�tҳ���З�K;�WD��	���V�LO��^��)�hs�Κۈ�춴�3�J�Q�]rf-Іɇ��r�6�E�*��(o�)�lK�"}�\6�c��U=�W�5�x^x~8}FK�K�iЎ#�4�f��[�4��Ri	��J���4��~^�C��Kx�~YiZ��=)-/��Sw�v��xp�u ��4��
��@�'�����}��0�l��~�b�Z=3�i,���M��F��ʏ/8x�:=��'�;�����a��j|���&�t�J��9��Uȡi�o��gu��H/��	���z�}Z+_����qun6yꘫ�r�&}�����k������>L��ܾ���$}�O|���~���{���t&��C=�|�h�N%���-aդ��5XG��95��Q20?�wg��@�R�"-

�=�:��fဂ�r>!؝*�*���l��f��ݎNs6��%e�`�f��}�F���N���]���YH�xu&#	��@��+Ҽ�¥�bDm�C��,iZ�n%~.$_y�����f��	�iƳBN���d���N�-.zՔ2�K��P��p)���5�Q)��;eM��š��	���vr����y��sڨ${K)��P�zϳ�^&2i�U�$��3o�_�qYR�:�>Wz������h�gQPq��bU��5œ	
�M>�+����z��Ò5��:CI���t�+@��c�۹�i�i�V�a�2��YqA���>+W�� �Q�yW��r�<�W��9�<�9�&�]��ŉJb�R���y��ˤg�*協Q/R��8_S;��;��	~;* �'�n��lm䊒6���`�<�;ӱR��<���7a7
�$^�α��B�PN�:��e����ͿҾ&�=O��/LK���WA���se]��,\���b��[��G���e��Nĝ&p0�c���4%�E�i�&T��5pp4�R4$�4V�T@ҋ��� G�>�ax�܃�z���p]�9��}�0��m���G<��wQ���t���nw}����0D�����G�'ݵuI o���r�
��8�#�V���3�8\TD�*`�p3{=s8"�E����g����p�퟽No�t��'��~?N�!�h��q����.
��� }|-�JXs#�Y%]h=���l���Y_+�Ъ���G�O��`���4|��S0U��Ϭ�9������̇8d���D��{s�4p��N�_�C�l��*�;1��H�4W�џR��|�j���8��1�������1��^ �J�ç�9A�ЏO�g\=b1@>C~�g%ґ���υao�f�2Wa����>狁����O���h-8�W �*�gLW�Oe����m����X妪q��y���_)��{�4��6���,tD>yݤ��Հ�3NT^歽va+���E¿pV	(P(+.n~����9�&~?������n��;�V��� ]ڏ9��/�AO~�p��,����\�_}�lR�
@����#]�B�1��&i��l/uJ߽zz�pk�s���8�v���c1o�qn�^E0E`��#��t�.d�pzh߲w��6O�^ ��[����,�y,�A�{ي�	�J�3��p��j��?2�ˉՈA&i ��-Z�+4�	v�������'�ӆ��j�����я#�o{h�;+-=3}J����S��N�q9o�Y�v�%���O�?��Ҍ~�ůQ���
����h��u���n��_e�C��TZ��@���t9��-�L�/�s4yG�'�Ūp�|�=!��Bi��4��,?޲At{�ѽ�az�S�R��o�����WA�ln���{���:}��T�s	<��8�U08W��$�� �t O����q뺔��2��np��Ư���h0��w������{��>�}��o�o�9v���PG�X=a�F0v";�\h�Bܷ:�҄RM1���d�����\`�>�6�<�H��d�V�#i�}�D����KE�F7F0��,�<�Y���of��Vg��-����a����,��f���Y��AZ�jq� ��d�����m3О|cgn�C^�K|-ȷ'�����X=�v�2�!7����6�6�w�ꛯ�� ��S^���(i^עa��U%��O
?��8����>*���#>�@P�I���s��[e��L7�C�	��CYY���mp9�j�sa1Y�R+�/�W�_� *�<qMO��-{نJV��%С���+E)0jZ?���WV�3��vnA�7U����^�h�-������������$>b��j��t����)��C�D��>'m.�,�ݚ�����=���<�U�\��<{�l3��e�{O9�":BZǦ>�,���t�<�z�����􊅬�f��3B)?�`����B�(���2a�z�P�l���#"�g����<l�>����$�YS�uZ�_�QT0�#�r�ʋ�o�
��#'���X�")wx*$N�R�@ꕁ��դ�E���u\^�ɟ�K̓vΌb8s�ޟuu�T�n���Ƞ��E�J���g�w�O���r���GZ�^�x�y�M�Ge��؉�o�z��r���{��L���EN5���/�r��}N�V�L�Y��Z���َJ��l��]��N�V�ꫳ>�^���7�����z����V'���[^�'�
�CK^�I��LB�r� t&�������}�ޡ;f����k���8������ۏ�s��@��OՍ�E�q��/���� ��)w�G<������P	��cܨw�l�,����QT��Ȣ1��Q%�n�98����ç>M���^{N7����>�k~J�:���{���A���b2.����4��f��g�pD����\��i��B�F���d�ui�_��1�l�b�I����ur�JZ�ɴ���iz^8h���GL���?�-@*�����׼hZ��#..}
�C��v	�>t]^�Ut ]6��+m��!OWI�kަ��.PwxǷ--�q�� ��RAV�}P���NJu� �[�䒷�.:�yAR�����i�*�"��6�<��W�j�r:2/�m�`����B�z�*�ŨF�>�t�,�4U�sURL]�W~[�~!߬�`�V�T��K�%��n[m�������:�����-2J�tX3r�ГL�dX�_�9ڪ��u�=��x��=6x�4�sa�-35�c ����<�#��sd>E/�6]�dnGs�$���*
߁��>\�sئ���'Q������/�N��1X�%��#���z��ܰ��.ү5�=&���t��VN����nO���Z@��/�;����k�H�k,�Jc� Lc�n�r�]
����`�[�ْv�T��q�#+g�z�j�?CmiF��y��i�g!�����{Ξ��� :��ġHSt��[j�*ꚉ�d�~���UmG�Y���iJl�y��w��N���<�T���ua5��N���-��>�)x�A#<��5,��j�]��J[FƉu<�ޣ��nG���8^{�v��!��]S76v��ks��:Q�\`��T�g����a��y� ��u��8���-LE/-��O�Nѱ�Ɓ���!�~�jx~�����n>�a�ȏ|�^~�c�-8N�]� ����R�6I�69/I�Q��B��5�G�^Sf��T;HB�f�i
�F��'��
�k�3�;�3��o�M���ʵ�;wL3�Ee���G	/�*�T���F}2�C�9	��Rp|�>Lhu�B*xT�� u+O�6�Z���V��'���XN��D@���c��댕M\Y`(p����y,'Z���x	f�~<X�_r�/��#41�1��J��V6J��_�~�=�Pw��,�B�X�)�g�Z��_��֟�״$�!?I�v��T��fprB9KvlKXՒ+���x���ż��!��@��h��-`�{�'x��p	�kO��׳��M�Ϸ`e{���	�Sl_��:�
22��9 7�7��[W�P9=��v�������Y���������w0ա�g��7���g�.퇩ɪ��CL�UÔ�L�62m33�͜Dr�jiVy������c���r��־�Á����_qmo1f>�x��{5O.�50G�Y#�̓�źm���h!E�N+��O�uZ��r
?�{�_V;w2>禑z6��T�L�-�m5��i�/��&pH{YF?>���w)��b\G_���L攞{��bq�p&܅��<���������/�
�z׏/Ly���O~��w���v�l�����p�Ҏ�q�tI>�z;G5.St�� }9��2�����TXL�`a��C5���8Oz�﬊�x󆏑��X߮������;o�[?�U�z�n��x���9:rC�����]�
���)m b��hJ�y��~���B�q��o�H
up���M�g-"䷠.�H+�+4*�t�	�V�\��p�:�Ewc-�LÆ��ȓ��M��
�ҧ*|ʛ��W�Q��<�hH��ꐔ]z�%
�h�����h����)� �#�sGbpể�K�i��źcj�(�<YK�4�:\�|��pL�rŘ'��v��Y�\Y�v�gn�
&�	��ě1��)[�"_�*�.������J>�4�/iȳ���A�Up�L�^�sW�.��ʸ2u�fЯqH������V�[r��aO����*��W�̹����}o�lM��6>��j��9���3�op�~��P��:n�����Qc[��g�焷z�ҖA�Ȳe"��{�hc���=���(k��t��G�U����(G��Pl�.J�g
�Fk�^���%e��Z=K����N�"N,�N�J��0Tz���8�ll�U ���٪�N�*�Yc1����%Ȅi�&|ں�Ns���aF0Z�6���,?������Uy�O�)�8wQ�jςJ��^���8;�����U���]�	]��]�S��V�r��4��sJi?�q�$�vr���|��E�Li����qi� �b�>��؅�㫫��v�kz��/ҋ_�'�|��>���)� ��g����%�wM�;sj,��$�ǁ�����q�s�oHc��3�Y��'��X	��~zr�~�����/|����/з�}?���a����w��IA�G�y���<ډ��y?W!94;-�jn��[f��2��z�'��Si�r�9c:u�Q
7K�)ڡ2m��5���4O�U�Im
tA?g�#�g�i�N�\F���3/!�U�ρ�I��O�ǵP�s�W���clz�=n()b��!���K��ۗ��5_>�On��C*K����>=�M�ˤ�6p�9R*�#��ֻk0��ґGX�a��=��V�$��Z+h���M�N���|�
ޡ�O��gL���{|��2�鐆�l�G��>���K�h���$���!�x�f8W����)�C�+ԟ
��j�\�Q8����%��kճ�2s� ��8ƙ\�]�Ƶ�6�E��`�ҁpΚS`ɫ*.�k`k]gm�vT=�*�� �(s� ��4�nN������|�� 4O;+�3�7�`��!��7�]D��+�B���j�5�2�i`��GMo�to<CM��W�D֤Է�yJ����5@;�Tv�4�51�k������g����[ ?���]�
ϵ�Ӳ�^U�:.w^�,���ث8ҟ'�Bd��1Я5�+i����,���7�%f�Ő/�n��ڸ�Q?�/�VYV/ǽ�Q+�A��/�1w&�~q%s�h}�������m��������(Y�j������oPo��G����dT+(�\��>�9HVkX�t�棞�']s$����OP��/���~�n������1�sG��p�]|�Jܯi�	���T��.=�cfK8��s�f���"��
p���i�b@��q�}�=��`"�?��DN2|p�u��ϑ�ʗ��#	o���~�<Ջ���^�w�8�O���z�oYE��lCB~2x&͓Zi�a4}2�n��Jh+W�礱���m5�R�TZ�8B��t_-��.��S�_Tª4�VhGWӦp�L�2&b��4��y�͜�1m�	!�2�i�A�H�#���,~�s��1�Kz�N:p �5o�Ϲ�Øt3�k����n{|�'��6C�dOJb�S���u~�!���BF�(�T�= ���s�PG���G
�ha�^��<X	p$��l�'qm?��o�G�c\�9��{,�!�K�%A�+|�E�>I}��p������-�>��s2�bwKy�\9�5�8Ű����Y�S�S�=L�%},��=|��'C����8�U����
�?G��`�J1��M�5<�	s֤ub��������'ݧ��d�lM�����8?�eC�1�o�L��(k�5�w}��A��I��4s��/"BZ��� ��K�?�r E�6[�:pl�|�}I���	prPY9wR��s������K8�9�.�6�Wi\���_z��[����H`%���6�'C��� ���J�j�Y�6
(��z\K�{~�-a|����·ٶY��X��eO����~zK5q��:��vL�e�ro��10u�B��ei���I6d�bZ�Ii��/]>}��^m�¡�NJBz0~s�Z��o�{�_n�_�Ղ�}G�:Y�� &�X_���=Q�Pv;�N�g�\^�u9!k���Zf�݇��`j�=t��It
��ո��t���}�w���_&��wD����COW~G�n���e�*�@����U��-s�Ηt(��Ga�+T i5�$�pQ��A	��ٮ��rN���s�ak�5����;N2�ߏ���5��3W_�~����4���3��y�cp����;i]h�{�J�9m	��c��R��<ݠ4Hȴ)ki�wVl�j�V�_���ZP��t�E�)�D��r�����;��(�xf���_�ˆ��rR��΂$Շ�)H�Q2/rN�3���&����u���ޜ�_\2�n�871p�z��_�!� �",��]�,��]~��\�٧��rq��#��O_G�(`$����6*�B�+�똅�䒬_�H��@/�F��@1QJ6�)��f�ԛ�y�Y��@����dm:MN�[ +��&XX�E-k%`�>�Sn<��r�����C���g��:�t��ܡr�dN	Kn�XV`Z+������!o�Od /��tY;^[���ڲ�s���C��<|/�Y��]�_�epg7p���(��PSg>��(�f�Tp�ZV�uI���,��m7ti�9����k��Ol�f�ԭ2�'m�.s�.˙�g�g̢|7�?��A��t$q�w��P���ޱ�di,�f.'�j2?�h�Y^� �q�wy���pN�����_]�O��`3��o�[k�#��+�����].��`v�i��Tq�4���i����d���+Ҍ�j�Õu�Ҧ�a�O�1��F�3��S��D��l�
W�ʓl=�L֯�������v���^y];�χ���'�3 �^4�cw$����ػkr��u�ޠ��I�g�v]G��Qo�뢭���i�6�%�=p_� ��׋_��9쀞����l���]w�
?����!.nD�k�:����!�����=����@������7ޠ������8A�+:�����>��h}�<gqk��F����v2�!�
6],�>�-+�+©'�5_�Gcx*1�gŲԳ�$�4~�pw�VU�e��iܯd�YZ	���"��J[��Y��f*�>�;�2�5���K>_E*#b�k)<R�UZSr� ��(����.� �����97p��6����s�7�s���n��aњΑ�{iՌ�Y��j��(�F͹�5��b����ܺ~"%�v9t+J��kl w����G��t�����ׅ�g�Y�S�U�&{g�v �l5�w�>~�u����o��Ṭ�d��K>?A�����z՚����]���u�ʜAZ>�����빤�Gw�b���`of�c�cƛa��^u��ũ��|c����#��O�)s�����KFyJ6�k�q�/�6��>�m؈�=�G)�%�-<9�{+�m��W9xn�I5���o+��]Z[6���5�jӪx���e5m)7�c�-�s�̓Y��s�^5���	<��V}w��`k(���#{׾�$G�q��~��G�*��nݎ��a��+MT�r!��F�0���~�t��E]j�����DU��TΙ]�Cb �փ����5��v���/�F�D����V����{����g�;��/ҳ�5\O�7�v�6�1��}��B�w���^�}������F���d^�)���R� ;M#q�U[�4�Ӈw�o8P�w�?�}�����}����8�x�-:���ͮ_�¯J�!�#4T��5��t�p*;Yѹ8��f�FZ��s��K�_k.(����4����f��a��4mOr�H��b��?��H�4&D��ߠ�P&T�[t/V��~aw|�=�@-�V����� �/ݴl���#>Uc�
d�r�{`���߉VDAY6#�L/>}Rd2��2�$�b*��s�91ӹh��>��O��ʍ��A��<'clD��C@4���E�&�LK3%o<'UN�� \E�\p�lE�,�+���h�j{=���ܥ�c���FUC�Lխ�CE)�!���lXP�:�-�����������7P�]�C_�M72���X���_K7.�� ���~��֞'x����z-n��S�(E}w��ЏN�Qvm{���e#�I�v�e�w����8&��~	��F]P��`˨��C�(�E_r��(g�
�޶֫����5�ҮT�������:5Z&ڎZn��n7�h���n��k�2M#�3l�ŷ�C�?�͢%��O����/�~�:p*���)_���{�6g/�ڳ`��\�(:ZN+M�d��>w?��{J��	��>����W5M�S�*DU��*�{ t���J���S������?,�Y�k�s*'1���(�d9��/p��5�� q�C��S^;���zH��n�s��щv_�^�����jK���t=��s8]���v�������;Y�g��hx�L��i���� ��
q�N�t�����᳸y�����=�0�=gs7ot��ۏt�l��O����ا?<���K_����p�Ƈ���Ǭ:��O�%��=�Z�O�t�ꔃ��m<s����&�ZF��*�����u�b��i�#L���i��I�������LC�������nڎf;*m�˪S���s�V_����+��q��*~ �]?�����S4/� tT�<��Q��TP��?�H�*h&"
��KF(xA�h8���K5<�NS���	���p�i���riUW#Ϗ��|婧��Bv��C��8�\�'���<��sqG�C*<rjire.������HX��Љ�mǅ
���Ld�Y���[�s6��"LS�n=�.q�<���%;٧ٓg�S���(�ҵ�q��g~֏���w���5XV_��^>%3e�u����5�#���[s�?���Ճ�t��e��k����:STS7L,��{�U���|��)0�6��Ƶ�G׋�4�9���Z����L3}[�)|�C����#�p�nк$X:���M!�q�]��5��)���I�c;�ϗ;s��9!�2�sFja�Ѿ�M#��{/�2��9P�<��	2������(�������ňZ����dcf����iV����&��4�JS�	Cl���^?l�,�����8Lk��d���j� �sCY��@��9��4 ���GE�)�Þ`�p[��y�M�
4I�JOV��$WOꊑFD?	��9�Y$T~�j,�܂�X�Y�qi�n@�_�_|�_�����e��S�*�Ԣ��ً��3'21{�re3A}�%�2�.�>��FFQ��SE�5�){�\v��O����Y��<{��q���p1�w}����/�������q���n�i��+0�W��Z�l��ڬ�"��{����Y���cX�-P����o���J����������@~����{Ǥ�������~���M:'���~� y��?�O/�^ܚ�m�Q)���*���r�\v��榕;K(Y��P�^;R�}�Y��i���m���ծ���C���Uc�1PE9�(�6����i��i֘�QA�V�����8k ���b��������i��'m3���'-)О�.Qė�x�lH�|�9��l|w�c%�@8�4��pt����� ol�bʍ6A�.�R�j�qPhI�����Ud�`��>�Π6d�Z�rQ�^�/_S�l�hA��4�%uY��B�m9��	�%w7�lN���ɭ�T-؏y�Һ�7����v�P[V����/%�5��Һ��s�-�젼\����5��政�ul�ހܼ�K�}T�}����o��{B~xoNn��Q*m�`�i܌Щ_J�����F
"�O�8�X�jL�{���U����c��U��=��|;�����o�^-����4����J�b[���}�0��~�k�[�1�b���H��|x�Ӆ��K�4���Z��O<+�`�Go�Y�Z�~�*.�(WaM�}�
߮����J��pm:X�*�t97�;��:��~�����zL����%��TԠ'"�1n��r;1�!�Q��l5_R[�À�Z �]ȕ5vfڻJJ�@���H�A%}������o��?�����#���� ǎ�(,���w�>Y�^�l����nk-k�]���P�݊���� �Ơ�p��?(n���p�+z�G�F�����^��������0\��ëSC)����b��p�쭝�k���O�8�{��9׮�ۊ��W������i�Ҁ�4��S׉��bF]Y	2�Ee~^&~T���j3nV�F���	����� ��س�V�Uq�?�o�� (�"V��I(�0-_��t�N�����ƚ,����p���@���C��� �� ��v*�\`+����1Ջ5(��]Hh����܁��NK���m:]"Y	y��5<ob�����y&���3��70V�IZt!����w�����g>�u�2�9�R���F3��N��aau[�.Nkm�o��,�g5y�>S��G��kB��ۧ'x����K�����;nE�K������m�W\��U��͑$�1��{�[���y@Z��6�L���j/�U������d��rcSA�W��vL��kdk�8�QW���$�AK��Q��@��фHH�'���N	��� e_K3~*�G���{u�[��:��d���֫�ܷ��r0�7�6B�ɷ�!��6�_^q�`Z>%o����I6)�X��, ˗�ߟT�7p���p]Y�Zr��糰��E�b��2&�,h%�]�=����9�#n(��!;]G��p��3�=�\_��C5��#��ġ�^�r��!���FC]�4�TS�;\�k��p�����?JϿ������'wؓ�}vL;d_j���.E���kS��9���=���7���8z�B�<]�i<}墼����:�q�oI_��8���0QD��ыwޡ�~�t���ou�i�m���8an����1o��4��&�\��b���N���X���`2|���I�k�=(��%�VI��؊����Z}.�3�[̷���+��\�-Z�S9ӛ�b���$�3�^w�=���w�����3�Aͅ��|�u)����6��!x��yC(KUH�Qy�U��,��	�H��YߗbK�I;��?=R��	�0r��&�#AR��� �����*Vg��q�ta��Y ���X� m��ΒH�W�`m�@XO�<!M3^�Ӥ��Q�r�g��a���l��Z�]U���jg����RBpl���z�c9]?��j}�1�x-��<>)�f4L=�྇����\�sd�c�kA�+z�����&�c���C�q��-���U���S��\�Wq�te�:��}�1\�]wd=���2v��E���C~��$��Tj�O=gB�B��MЖ��j��CH�Sl���@�G񦉹����l;S��(��R}�m�����~隿�[���|e��<�$�xh��6X�k	�
�����F~���gڥd�区��:͕iV��X�ʯ�լ� ��^L�_�`y VqK9���RV���J9KnZ{1StעAo@'�-�:�ۓ�'!�e�	�m�#�6��ˋ�ue_/�ϭ�ܷm�H��F,�Z�Wɏt����>�׿�%��C7�����oniw����7���X��X���%�Q����K�c,���č|$���T�w����5��C��·���fxO�~�^dG�w;z�_��~��9U����������C���u��q�Uͳ�ʅ���$�yd�� �n��ZpJf�d����}e���i$GG�{"�7�M��y|%Ow?Nk�eo�i��.�T��/]�Iwg����|܍���c�I!͹B��ff���$\=�*�`�L�C�
Ò�3,��>$G}���CZ�-i��cHc=l�����}^c\�nm�%�'K�5��-^Β�o|���|��%Fr����e��c*ן��8��e�ܵՍ��Z���"��$s����e|}�QK7(v��]2�����z-�N��F�-�'���De�C�t��K"���}:;O�FlԂQ(3�2�	�(�_�#m	��\���g�sm X��	�V�E_\
�w�3-���A�S��*_����������e��;���t9�x�Ӡ��0�ǹO���!��
�6���ɑ�ٸ��F���OFy�]���WE�����mA�	W�q6��H���[���l�>5se6�l�5v̔ݴ�?ݗ�3}vy��9ɷi���`��)�P��Y�R��3B��×�8h�
�,sʅ��os��|��K�9p��^�S0��-�N�'�'��C9�^�#�t9�,���l^U��j�i��Ӹ�z��p
�Ze-��*�x��ԳZ;��*�j�q�4E�Tt*7k���jK2�S��K����ܷ�us��ǜ��4�݄}���%2L�.��ź������?����/�0]�����zcL�.�����.�35~�S�kݮ�����w�o�S�W�IlD�q�E�L4�If9&��!
�g{ȇknvC?�]'��%��ݼ�iz��?D��������<�C �!ܸ1�o��W�?�@�0m�H^�sa�,����~<ٗB�h�>҂�F���
��'v5�&��Lc]����+�b�+�6p0%%�%�t�,�����A{�oM�J9�+�}~Q�-�ʉ1���(G������S���9��DK�N�!���]�N��'�w��42U����ch�d�~ஃ�0�>�\
�t�>\����Gی�]�VpP�A�G���)/�KZ�P�CPFZF���\����s8�#�W�Jʏ3��*�si���F���RVђ��J����P҅�V���S�E����R4��TB��m��m$M�ԋf�dLJ:�6�X:�8L���fn��I�s����] �k6az�/�ʟ� ;&���Om�n�o��@�94j7t�~�x#��z�t<���>�����E��O7~,�����њ�xJy�p��y9��N�A�n]���u@O_BD�{xJA��K�B���?i��e?�ǫ�I��ù���[v�\�y8e�@���ryq:6�ύ�X���,��[MP�am�-^�>+�5��	��<?\j;�<g��a$"�!Z�QV�<��e�C��d䒺&m�G.�F}�ϳb���|x��G���
]'Y�*�x����u���pHj�i�k��/��@��_�B�3�v�3��Q�c{�4���W�FN�3�j�#c�o��4N�+������hwk^`SB�!�2�zFf6��D�<���x*�6���qM7u��(^.��P��j2P�몶EQ�?}����0����t��+:��~No}�+����&���o���h7�]QO� /�.��m�
�jh��N���p���I�|+3���l��kY`%���Q�w�bwM��O�[?�D��}��jx]�`����C E���C�>],�{�cq�}�=�����k���UdCx;����A8cҸ����u�p2��Jw��+iB0�~5�Ҭ~M����~Y8��%b��7qP���k�=|XtW]�@��p�3�8r~�p�7y+�d���W�%xS��\FB{�+�v��R7E$��� �;O��¡G��C�c
.|�����&tjAQZr��0p�s\�c%��zs�I(:�Y,%�W	��v�wz�">�sS�pM�Ga�����'�����:��!S*�/d�W��@��D��j�p���R#�ğ
�|���Q�,ŴЯ&ڙ��[�Z���C�__�B>����a��=�O0�c$x����ī��9�e�tz�Pb<m��_�����*��CF�Y�~�'0�Ȕ�����\�ˣ� ���;ڱ3�'�<h喇�Q�@�S;�:=I>���`<����hc�U箶M�gSv�U�+;�)_��c�&p�%�p��� ��8�D7�W�y�d}��y$�a+}��W�-_%�+}���<r������<<�*�Os/�(Wc�I&H��x&�b:�gh�5�ؖQ�گJ��O����7�}C�,�k�� �A]E�4�1Ѣ�q.D��㱜�9%GnY���'";n2)u}	g�I�G�����K-+�p*�q^\�`�s���v{z�zz������c��7�7�-���{��?]�a�@�vyJ-D���~��l��H���my �j��aK�YB���e
Wx�?Dwv�?~��Q����G����ߦo��4v������*^�B1�(p��"��+y"bʚ������v�G06"�pN�ⷶpHBqSrY��zQ�40v�g��H�ł*�q��[�9i�Nrr܅� �4���_�:͗i&�	�q7�7�t�t_��!j,E�JG�ʠ���b�1��`��.��ep�p�Dĸ��O��M(ǈ�2�μ���[*[��q���%�qm�q�\��)�}Hp��D�ŉ��	��|UI*����~��S�a�<|���}�}s��i1)E�rSv1��u2{�������V|��yj��H�ƳE�̯�ǻ�̃��oA��2�U>�6<@��&����$
���sO��<N���$t/�K�S���3:k1o��1�U6��ȯ����'x�'x��K��K��w	g9�Ū����ə���f��{�YG�'��6�3�G\�2� ����`����j.N/+������Aw�ͅ6�V!GeKo���>������&�G��YJ�ոe�X6Mk�݌<��F�+��A0T�]�h��|)|p'�ܺ�o�i��%��D���8Tz%��:��E���'ȐeC�}ZM�>�#W�����>���~��H[�M��i���W��=7��x��~U�~�N?��& �x1^rJ��T����T'����U�8�)dR>=�W���lv�ߓd@���{`��6o/T~D�l�ϮO�Q�|v|t���[��z�ޣ�_�Er�D�WG[�Ї�Z�>�ñ�.Tх��!+�D�J߼���we�.if} G4 ���H�U�;�5[�9Ĥ�x��p�FK/�h�O|�^���?����'������c?��ƛ8�h���i2�Ys:]������3F��t���M���d��:�W�3���z�����.Xv^��D+����N��v*i���i�ҡ��V��lzL�M�>ER�M�ܩ��}��0M�.h堆_~�3/*56�C��� �v�uE��w����{g<�+ �t�ZS@.-xc���y��t��#O�2z\��\���s�C������w��:B%-r���8rZ2�T����G\��򰤴8Q�F�B��P�F��K����
�k�ǢL֝�-�}��̚�����tC	��	�Y���
���Z�K�S����S��'s��%�����[��&U �[��D{��:��A��������]8����q�{�|D0�#���c][���'��l���gK`�t����o�L6�x���ӂ?e*��>�"�+�E�
[�2�*�*�'7��Np#��U޹��3ʥ�n�5�ݙ��V"4�~�v�bY���j�(�LK4���9���͈�U�J�5k�9􆽱%O�s-�+c�zO���Ȉ��.�B�� �K<�6��'v��B�گ�Y�F��r.�����I�:M���?M�g�������]4X��V���;��X�iּ�iY��{1�<R]x�.�F�#��S?��a�"n�/���B��Iz����^�{q�p�^��w��d�v�+����Ϯv��{��nG��W����?�e�/)��f*oL^�ҍ>�x���^�m� �j�}���6 ո��+�V��S�8���;�B��^���H�wc�S��z����ֹP\e6F�׷D��U�����˫���$�~�t让�}9k���Áv���\R��1(שvF0-XR��'
��E��2��͔
~eJ�6
A��^JT����!2*҄�	�THO��f��Xr����T�sB��B��l0)s�?1�iP?��ż���(�RS˓�ln#��tH���o�N��^������I�c��kZIB��&���K��/��� N��L�]���_��I���8���t��ON �kž��O�O��.WF��u�<����	)]�
��$g�eщ <@S;:����ا��+�\����=�Q�dU;�芐y)��o	���H��y�I�'�l�O$0kHFŸ�|
s�M��Br�#5i���Ug+�՞�\Nt���.O	��4b{TJ��ڞǚy9�3�	�p>�����u��eqkZbZx�u0w�/A�+u�_`{a�:��.A;qOۘe����3�V �΁�1�5`dfTc��U��<���̲����t����m��վ��yU�e�a��o�y��Nom�Yr���]A�_��|�f]�l!�x���4��������ht��<\8�\�*hc�a�*��ࠬ�賈�N��
���x�)(#��.i3�wY�P���%.l�Zv���ӈa`=̈́�d�g^�s"5���q�J�7D�'ϴ����l%����6�l�J��ԧ�C.Ze:�`�(w���l��a��K�:�w��ȵ�`�^]����4h�T����#s�7���`k����ϝ?��SuO�3��o�m��l�~��H�]��0+-�'|<e~��Ҵ����`���Ȼ�_3pOn��dW�v��U�XtǴI�%e����}����T�������!֕����N��$�p�&>�|}�.ՙ��Xw!?���h����XjW؏�2u�ݮ�����u��sG���������[A�9���.�3�B���"�*�1��O��cZM��Ga[��%ÿ��<9��&޵(��sw�@T2ӆf����y����KzquM���0�^�h��|,����~h p��m��p%�zܑ-,���J�yGҹ�ΰ`� ����u�R����N�%����<:e�ͯ�_�SiZp��H�s�4-p9�8�rV�Z9K��P�z#�qg!��ą��*i��i�y=��](8ݩ����'v�/N(YY�l�0�8�L�����n@ည������4��?� ��v���:N:��XD�Pii�x޸iNІ_�9A:��hX�	 ����o��>'��+���k7�Ұ~�V�!����"KjM;��۹����o惾1CO�l}L��jG�S6�)S�������z�������	>ٸH�n��j�չ9�&��u<o,
s�o\���"���S}�_�E�-d/��_�y`d-^��*{���	�l07�c�S�e(`ʑ�P�9��2'0am�W6�/��w��[��>@�Z�ԍOJ^%��JԤ�rh�]nȢ�Ȫ���Ȥ�脥�g�27�n"�%i�椳�CD�J�*Ͻ�G��f��w�f��6t�lF�o,
��읨7B��<|!К�Ð3J������LlKXQ���� �ʁ��I�ku���n}����܌�lz Ǩ�(���!�;g�>5T/l��M��k�V���� ,�i��t{��7���iD
�~+�����4~��P��o
wk?H�Q��b��T��Bw�V���F5����N��s�̽&�	�Px�<i߄m5�[1�!^F� �{0YO��`��	���	^�3�p$���`�YKN�Z��k�8��`�t|�9�xه�ొ>����r������ћ��/}����ߠg�����'���=sW�w�j��΅6Ъ���R���]���*��g�pr�E�[��_��\���HI�pu���:8�g�	�������7t�=#����gC��O؎��}\�4d�6�9���\�D��ʑ`�h���Ũr�sV��I'�tI/5��g�̶Ĭr�̟hg��Ђ4h��r���P%��7��E̕m#�	��s
�J?���BR�^�	�i���4�=��Y)ɩṜ�m�l۳ p�\�и,��	ߋK
N�d��I�p�R<)q:��l�?�`8��݂^#ͼs@��>g��yHc�B.�8�b-�ZJs����K��P�7�rD�CT0�lN�������T|�s��H�x�f��R ��J���!�IUI�)ZCH~h'�)�>8-S8%U�,b��3_=�����F��HZ�G����XA�~|��n�+�Jv:��[<`S��	��};��gs�a=�&��nT�$�~̵[[e4��4��R��u*��=b^݂���t������\!NF�gԏ(�#�>ʯ�\���l�tIw�'D5oS
Cޯ@[(䱖A�7�N�K8����7�h��z-�L�Ě�b�Ch�h���l�ʻ�/*p���_He�k<�n"�m0\	Ɛo�~�L3�����S���:$��~9��]��!��?:}.���^Q*�E���,f��ă�)���J��n��hk�w�eե�\fZ�2~�Ek����,V�qfW�y�_�8�v�`?�p�!>.�W�3%}�Y��(��yQ�3X�@)�{#��xMt.�~��la��{l�&|�������)zHa�s�Ė��S��ꐼ�%t�_���q���.�9�4&�X�?����=���Z�s��7ޠ����������������p,�u�z���C���8� �W���A�����>]�,ڝ�li G��	iWG�[i^9�D/�X�&���q���A;���7nnni����5��6��W�����ÍYIHJ6 ^]���e�f���¿N�늂m���*7�J����U'Q��WC�0�t�s���.�弓�A�k��J��;Up ����Y8X�Z+�L�@�Z9��H��Z�S�Z��-��4�H#���v��S�3��$�Y��d����]@�� 1��z#)#/6+��+ךϡ&q�+.���e��pQ]*�`�%� �m"M���`|�]y]�zIk�����Qb���}RF�q�h���!��bi�ϠP�7fJ�Jg��xv�нj1�ǜ�afş����ë=�S�}T���!@����6��+-:�%�L�7 ��J	����Q�6�2�"�i�KqLm�eۣ���{~?����'=�`;�Z�.��cn{���K���W�]���*�:��:���`ꦕ��dsvQ���1�����/_۹�M���ǉ�*�fqU�}�}X��$�W3���aN�.�<�/��`rPR=̄h�L��f�s�pi���>�����
���N?�ߧؤ�#0}����	A�4���]�>���cK�m��~����~�:���Ej��9@�5w�	��i���+#_艃��;	� �`M_���!�f�Wr�9�W7��J9�#��-
)��f3�	���A�a�o�c	��~K�~�~��M?��-akԙ�;#�ǺF�x�yQ�S��uf�&Ţ���T�k��1�������N�_�y�!+*dׯ�{�l}��(�+uGK�p�^s>>�_�%�C=��+����?��O�[��}���}�����ut���ݮ�s�oʠ�-Iq���[�g��&�����C�wi�,��c�o�0NJ~��8��Ǩ`v�{Db�`�V)�Ч'
!��SK�����z��whssT�t8�;fSa�
:DŷO5ƫ���}
��G��7�ؙq���CΩ*�,V���9ȁQZI�g���|kp����2���\s9�N#�V@�&nҰ�@h��,!':���3f)�n�i-��:�����p��o�`i��2M[|��0����i�_n朱��1�Y)��W^��>�QxW�Ɋ,K����(~!�H��,�s����������:�!0F���:B���b�HO/ߢ�|���9�O|�`%rX/���l �J��4�}��|���u�eVbe{41gt���(����e�V��[mI�9�T�؊�d����Vm� ܤ�~r(�ǅ��L�{��v5�~p����X�η!t��<��|���=�����+�*��t�y�kݓN�Dѥm�lç�<Ҩ�ɺ�\ɛntF��N�
��rh��@X�gH�о*u�n��:�9���u��������l[툳��m�C '�ni���q���~������ķ��5�,z`�˳iHC�P�S�Q�t����ӴN[��S�F�q�k�kq;?d�<���AMI�����_���a�P�ׂ-��HvONs�T���^�5.�&�M��׶q�˾�j�ʶr`7���({1��X�:�����=���2�wcPz��}�gn�c����ї-h�hk[�N��V˷횩Y�S`�����Fvo}r�P����?m��y��
{z�V��+��KwG�f4~8xƋ�����~��Ei��K;4���#�3�Ҽu%��x���&�Q'�n�#�}w�ge��pu��S��_&��i��?��xL,}���� V�m�r>�Eٌ���zcI�B���N1�����cs�)}W�]� �J�������o)`)35����_�_�����ۏ�K����\O�����1��C}�D�?�.�㍋�q*���9�4Hj�-bB�_�;W�{L��S%S����P��8����XIc$A���at.^�'����I�HT&�ᰧ�/oh� ���b�n��x�3̮B���.�­�>�L�̿�%ij�jZ��%n]/�!R8;�T�)Ҍv0�s��\0�@ש�w$l�_�7�f��T{���`7pX��ng
?=�f�n�Bw=��{-~�� x�A2�J�fCQ�D�T,���"�"+Ǹ�j�vyư�#����u�����P�C���S�����2^/�\h���`x�0�'9�����Y���2��H�u؄H�v2��,��ߎ�|�te�c0c:M1B���4������gB��|�t��7�&u���m�1�v8�v�W����۞vݠgc�|Y���r(}�ůs���=>��/���^�y�%o��lV�jM���t�k�p��p��=gS��p0�Xu�~oٯ���)����b7�mc�1G��;O^��5��A�t�7��C{8�gM!��K�及q�읍�v�pc%'���g��-'H~UF���m�I��|�`�p,/,.���2�,m� �ӕ�K]��Ġ.�҆���e�`/d~/�U6��~�B�R�i�>y��/�؏7��xG?���c��xql��\����..S>H7'{��i)�]5�qE���	�kbb!�ħ����r&�p�{Ys5����ۥ�T��&$oH�3-���<�2����� ���'��	.���:[�Si��-*mj�H��*�Q��\�g��s��b4j����~z�	���3�$�Dj�D�<� }�b)I�Ȥ�� �da-��q3��<壭?� |������m���?ߕJ?��KG�r�K�~���5}gwL����ǿN��{;����N�G�~{�w��>������bc�.���}'���wD^��5k�5.MV�ܲLlt9�����[�]7+� ����9�{�L��y�Ab���p���/^��vt���ޥ&�pcHG��ց�9�^k���*u��m2b�w�TX,��s�g�W�?��f
_�V�����B��*u��A�[�C�\��
O���fН�4����]�V��-iy� *?����1(Y�uz6���8���B�\t�<hW��PQZ0��8���+HR���OMA��9�s|��"(h=�u�17��dy�%�l&�è5����ٗ��O�FV>E�o$k&4�	n��!|����D?=��s��F�Ym� ��Nw��V���{QF�G�GA��*��o��65~v��P��nG���o���o�I��;��n���|�F�y7�G��Z���2��c�C&O�3>!j��ȓi��_ꉡ�3����-æd����Gv�w�@��>���:��"���%�a�<�Mf�r��u瀩`���Q���v��F[��Ї�~�^C���`SV� 3�ϩ�����\�Co��5���
� C6X���$�?���K�;Б�aUҊ�mS�Jē�+�[9�Zi�죹y���*uw�m���:�28��ǥ�?��>�zFW����7ߡ������M���+�[�?��v��+#���Nh�O����3>u�X��Xzlx6a'����F���<�\��,rz��[���L\���o����;��(���.��/��,֯U'I��܋!���
~s�b���p,��WwZ����c��_-M�k�9��9�O-[�!/٠8+��}j�ҭ��HPO �G���>J@���<V���CН������ hkR���1`���G�^���}c�����}�+_�O����Ʒ�t}���nyS���;�f�4_�WK�`�P�7�=����� ۏ�� 綺d����y>�TK���`�pM����u�!�ʁ�N']���QHÒ�\V�5h����~�8Ys�x�	w>�W���i|�`�g(�A��_�Ki�^���B@��Q������~ܯ�8���\���4�{�_S������C>S��:T�4mY��f�2� ���2���GNT���Q�A����D�XC�Q���E�a-<�!�<6ɀ��_�࢒B��e 絓����H�Ű����̇Bj��hײ����qb.9�?������4��s�̓�-gY�$�+�s�a�_?���>�FfcMa�S`�~�6�#���.�>ʎ�O6$���n^�W��g����?K?�����9�������ߦ����}zowC�מe�w<'�DՠE�/qOc�h�����+ʎYMIS$;~�ϔd�����/��ǿ9�1�~��}�8��>�+
���}�ko�y����U_�fKn	Z:��u��8�Z�\���n��!���������p&H:��3�ûXB#7&�4�{��@�Fh��� �'o��42�0�ҧ���׵��Iݍ��Zo�'��时Ei��Ӱ&K��3m3�!m-{=*�N9~b)�'> �<*����������������'�z��_��_�����M�{��txsG6�>oQ�M�o��a��3"8�Z���&a��C��^N��E��*���J�n�Z�_ѫ�7����mm�w^g�ɘ��wj'��e���F�k����,c�'��lj/� ���(�5�-޳��.���C��){�p����V�9�����\	��\�֌Rvt�S��W�ڌ�r��e�m�ǁ��į*K;1�߹p����}[H~�"�N뻗�84>�����n���;fx�ut{���'ޥ�?�uz��zz�����|�^<�������t���w.h����K¯�7~,�7��O�l��۹`i �L�u߰���ͤ��j�+g�צ�x�")����	�U7FŹ�'���<�Wy%
�{�¿�	��c�~NC�F�nn^��IG����))�7>�h��rfy����K��3�_sq ��*�Z�-��_Ik�[��e-�H�9��z�/�,�DV���m��ѹ}�b���|X!!�[)e�܅�<��ꖬE�#8�|7؃��[���_�~�����D����,�Mg_�:YBy/�7��H&K�pj zb���G��a�~�����0���gN�8���>:��I�Ȓ�:���m6C+���k��g>���¿N���w�uvC�����G�Ɵ����������kG׻�M�A�E:b�!S9"d���|%�B���4TX��?�!�l������Y�.��פ��a�	���\mH��	T��5��A �ܐ��Ђ7�>��������v��X}�	���J��T�m\����Բi�雧��-�
gh����
T
f��գ͂�m~.�I~yKo�$�b.R�yr}���/Q�����6�����s���M�P�*�;�ő*�H
�8�9��W�K��?������������h�����>�O����{�?~�����qm�1`x�S7�	��S�أ�'�K���vv��h��6�Ѭh��]��	��1�C�t#!�ۈvN�I���z��1�č��7��Ȯ��2�ѥ�ti�H���V������>�-��?����G򙖰|�5�:����u��]E���Ήk$q�+�Ix{���.�/���,g�H�8���W��e:�ó!�"�Fjxv��v�W���h�t;��UG/>�!z�G~�n��_i��z��p�ϻp���
��q�BҘY��J_�*cE}cn-�S��� �?��/k�<H�E��1�I�;��&�x˩�~�LT�[5ƀ����>����H�~�u�y�w��}�,�����П}fc��e�{��m/ߕ�.E�c%�Y�]i��.�����+_�Y	�Π����͇͘�=Ӊh6�4�n���l���V9,\D�lgQ�	�����ז����攛E�9tw�qO0�\���p�DE'�M`o^*
�������h�b#��˖uKIi�9����՛��ϴ�7$�������0\M<�F�LK�0�,}3��@���4�y*�LK��R�h`��x����%�ĉYpy�OTJR�9�U��g�T�:�hmFɥ_�^X��x�G�����AfJ��*K� d-�Ӓ�U'�E�1=�����ǯ"½����چSb�Ɔ����}�zG����i�ޏ}��۠���^��C����_:�ߢ��7���M�q�	�M  ��IDAT�z}��ݠvc�]BN�aD-96Mo��Pn��
P� ٬e�i��s.�o1��f��0�)�_qt7���M�B>�h��Y��&N����E����}<��ړ|���dW��f,�'�,�i��p��/�޶��_O����	�Ƒob�����:,:�ɣ�;�q<��ɵ�j�O-��u�߻�8'~ajN[�i��w��k�O�Bs���K�j[`%*��u,T(8�N��5d�)0
���r�z�<�g�:M���0�WґYh��@�<�e����ڍ���w<��6�4��~�K�NƜm-Kv���sf�;����"M1������%�i�@O)C��.jt�w�$��Ƿ/x��d\��6�~�C��zv�g���џ���п�3r|�
��{g8y��������W�=����N��˗tx�,k��>o�~vx�2on�ؾ�]I��O�|6E��v"|Z6����	�B���x`��QgY�\99-}������8�F��iZ�[8��bQ,+��w�~,�,�(���]�J��Öi��;K�V����1��}�:��Ҥ�A��T��8��)��,я�z�u.�t61C�[�]�sa�O����"<Z�>zڻ�/���@�������_�?����w�/���J����vW����٥�&�a:�i��tI�V�/F�ծF����E�-�.c��.�ůPI7O�lpN�%V;(n���~��:�4�)dA��,y,0�q�8_db��Tũ�,�����E�Ӭrr�k��2���*G���:��T�U%sx�Z�B92p'#���fж���N��%ㆾ(����<�u�'�+|��2W�%�AYqC'#e�(�r?��!����ؼ#�,�-�f�S��y�0A���g[�܍� 'ҟ���8{/�KZ��9.*��H�(�W�M���o�β���b���+:6�R�|�����E,�KN�h��H�ݚ���f�i9T��G☑�����tj�S��9�[�����?����|����vq}7k�����������/��o����~��]�{��?nX�ƨ�n�������'S�$���!u�w2���I��<��X;q3q��X3����7Cs�j�~�n۸8؇���,�e�Yj>�<� �'��ĸ:�Ԡ�d'�7>]@��:��.����RW��%Go.$+��Id�(g���������S�g�v�b�ޫ�;�yRw�4��u�Vm����~b�7��ɓkN~���W��������v�i���>��x���������I����][/_��po�<�������'�ߢ������wn_R��`�!�}�u�)��=�Wh�I�,����Ϫ�(h�������x�;���d��}k	p�m���զZ'�O�ܲ�=0pkU�z�Ҕ誹�����H��p�g��Nk�Si�.��
�*s,:-NTi[)��Ư�{Q����O�Zco���ec�]��ރ�P![Y#�)�*\3:�+�S�����?)e�����];H��.�&�)����G�Q��$�3�Af�������y���}�޸v���_%��=w����?�n#�x|�����m��4�K��I��~�����D�-��7p, g~����jp�����)|�a��iEQ��p�*����@���G ��6R+��Q�����k��AK��ʴ��3�_���ʳ���r���Ķ]�OV���˻:���+��OtP0���� 7m���г����E`��!��ό�|6@V��u�ũ�31��n�;l�)���Î���^Ţa���|_a,z]���
�]N\E������DD/,�|����+p1{��;�+3�nie�(p,+��_*�<�s�DE?߈���K���Xƥ����_T��Zr�l�����П���P׿��ڴQ���E��y�_�_����߿���o��������a��
�D;��`l0-���ș�@H?-�in��ց�xr��1�!/���.�g����͑��d��� 9�������M�z�W�����'������颞���o�a8�8�ڣr�$�n�qR���L`ad�������?�>1�����Ff��uƄؐ(
U8}�+�$t����)�Th�ڟ�yB�ɞL����KDa���Glg�����a���������?E���G����x��?P8g:D����{����W�+����������)��u���h#u]"fj;!T(�jv�q��He�ϭzg�L3
�g2˞��A���4����6lš3��Ķ.���?��ْV��R&�&�5��I}ִ����W��ER_���TD�4�����bj������Z���Ee�7Ր4���8����e�N�3�!�U���Q�v+�^�x~��r��K$8h益^����s��羗>��O����!���N�����i�k<�7�K���H��V��՞0�Z��{�4�c��;B:�Y"5a	��a�y��Q��	5L}���Z���n]����X|m�Ŵ��P�P�f�E�1̳Ҩ�FZu���J�`.~��֭�}���r�ҋ�O8���d���g����K�I� ���1M4�T�"`�ɾ	��n[x��7����k�Hƹ�N��U��E�}�\��L�a����&p<���P2�y]��>^����pL�L�ʕ��y���mJ�Ri�R�ۡ�u�
�H��=��U:�Vl$��<?}4��g�X�k���~���gG��?-���蜌��~,�S�������_������1FwF~��n����k�m[U 6���;��pi�) T� 7(i��64j'ݱ�V'��$U�JU�J����G�I%�J:�.L���&�vl��H�"� � * xy��}{��5�9�\{����w���o��k��xͱƤpx>_�"�*�vr�\?AHy��A�-���3��9;�� ����F�^�#�t:*��ʸ@�L��ׇ��ý�c���	s�`�e�B��3�<&ӽ�ӆx���c�,DpE��൬Z�W\�Y:���i��U_�$��� ĢV�5`>z=W�U�\V�+�&,Gi�3:Q���z��ԕ6�W�r�R��>��t��j�}��k_�"�.�Y�5����C�[C���7��>�a��W���!���j��E��Y��r8�U�u�]W����E����L@}�3ar�z�i�ߙM�m�ß��Y�� ���Is��m��ʹ�r���6mۦM�_+w���e���*�m��fA~�����r�h�����q��T�����i�F�@":qp�7�I}�^Z�'��i�^�EQ�d��`�]^���W� ,�����#p�-��-���o���
�k���(/���/s@���㘬�;�t�p�c����̢�17�7%��مV��"p�s0�`��a��qY���p?�b�Rqb8��#i��c!~d�\*z�g��e����Ϊ]c�7>g�U��]�i���N�C�m��id���a�geV(�)�|����:�@��rr��2�Q{��6��D�\(�"���o�01���5�X��
������4q�+:�����g���[�ج�G����f/7���q�y��0`����)��a偆���>ڲN�A�
�{�XV��<���霘Z�/E�r [®���t9_��A��m��9�l 񍝰���᫿Z�������m��"1�t�{FրS�����z�[��~����O���[�*�E�B������>��h5��� H�"��#9�P{��I�E��̃)2�u�KǼ�8Pl9!��W�oJ �����f�O���n�!�|8~�}C�����j�n�3%�,�x�~ߎ��7��@�CҔ��E2�)���\����e-d����񺭰��z��*yd�z�m ]��0#��2�j�)�f-���x�O�����Њ��_���[�<���6�"��0R�-�l��ʒ��Y�@]�J��m���zG�΃71�Ơ�����g>
�B[w���NE[��E�������_��_�����w�<1(;�E�m��>\т
=��g=UuRI���/����>��Tu�Ff�Ģg�_6��v=�`�C���Q�6���T�p|�^֚}�����Ϲ�r��9�4ؐ�O8mS�m��#��<��¼�u*?-Das��q]��K8���)�G�(�H�����T��ʼ��(C���^�*�pN�e�1�/_Z_��O}��U���o��׬�<�1�Y��8��
<&�}'�e���*h�,��7�B��+�xv.�)�����\�я}(G��.//�'�[Q�§��pp�mOڒ��^4YϢ�!	..=^&��p�uA�]D�p�Jc���W_���h�y����a�|6�N��C�5p��*�T�}
���ƯQ������)��6�O�}�Q(�ںb;N���W���P��S�:c�W�;E�(&^=��6�+%98�d��p������7�O}@)D�X���� �)�վ�f����u�Pc��l:�D�iE9B��zд,��:2��x��p��Zs��m���ʁ���J��������h��5�>��Z�v>|m���y�K���=�sT�b+�8�B�׫��<��;�7��{�=�ͯ����ep<�s��.�[t<yP}F�t���%�(q+{��<`5�2��ꤻl:�F�9:Ÿ��u��Ӏ���mlm2��Oj��+�{����`�C�/gA��:�,^��\v���!i��dͩdS�h?h�١CC����&�[Z���|���fy{ �S^�9&l��
y���!�g��-����ܐC�<X�:���}��g(���^�[�,˃}l(w��e&ǧ\���l_iA�����"Et;�5��^�����Ӟ�� �>�����Ac���R���1�Y'�n��˻�ԭA��n���se��}�_�k��9��W|+��_}7tO~,/�\ú��G'�̡��@X{�zjE��8`��8�J/�nkag�J�J���ۀ?Q񔁎���,�����y.0x҄�Vѭ�U�.?��^ǜ�֋L��ʗX��j��<ŋ�F���ۙ�&q١N�c];�!5\*ώ�������:�b:I9ɜ�8�O֕�j�=��6��b]=ɉ,���υM��u�ɒ>�.����9���K[`袃y:O��i��5�X������nO\8x�ɏ�#�x����ӿ��j5��l]���8��[4�>�,:�eNƳ�bD:�����r����W1b(�r:�̽B��G5�w�-������kp�קH� T\��U���!�����i�� 9�S�={�ڋ��(������4����F�j8��kZ���?7����_1_2m~�����]�=��<R��M$�)��]�2yݮ�to#(x��?��� ����ӯ	`#p�gG�!�M��������� 
��	��U�:��!}�ۊ�ɖ5��nD6����[�j�z�HhȾ�}��E�h��;K'~�ι�[��~V�E�=W>g�i~�c'�������
�:��������ݥP�1�Q�\ |�
������[_�
������^��vi.W ��������N��w��n��X���d�.E��ҩ��l��<�V�j���F�~W&~�˨�%���=�������f��ɑ��YA9�9��=�\~;�swJ���g��k�����-���&9�k���V����Zq�k0���:/8-�e��uO�=�?�+قQt-9H���3����� ��Ϊ.��"�G�����@5�ʹ3
N�r�ȣn"�<WH}���N���7R.��=�@z�`��_^=F�q�>^����>��~΋ �"t9��G�DʙAgZ�����?��O|>��W�rq�#}d�H�C�8j��_zF:OMo��Jcᨲ�����kqZ�Ip�r�i��}�ae��{1΍�[��)����SqD-��ǯ���t�1�~˄��*uVq��6��47�~�/�7���[��v\��9��Q�u�ٜ�J�I����?1�p�]e�ecV呆Xi�|[�Ƃud�%�$!J��+�/%g�Y�t��ς�ϲ�����5\>� ,���_��w�XGNOU(�b
�M�q��5���.[�}�������ก��5Io��^�_�N*�����@KD�TxCVo�tNؘ"ͩ��ҭ�5�9d������͉�׶��~�Q�W�6�W��}d�xbۀo/�C]@��:���b`DT�i�:V���҉�I93r卅]�m_F�$\Gl̆�y���(�,P���rHp�2�(\	�����ٓ���������% ��N1��!~��oR8��mW��+7ZAҺ̤˃r"�c�s�D�	�p|}������z�9oy��|��w~^�'�5T�@��x/J�� y��ud\,����7����k�˻�n���!�K�vybin��;��y\Ґy�L�aaJ��������@��%>gWj^t�<�t"pĿ#���Y8��p��j�g�/x��Ϧ���Z���2(���(�v�WE瑑!j:�t��a'�G�O��º��O���&'��"�`F��u!�u �[�f�u�Bs�k:��ݸ���5v��ǁAg)������ԏ�O�Q��љ%���[ ����_���������K/���2w	�EF}�Ӆ�����g}=���_��܁��jP�IM���H��b�VO�:�-��8�ю�ޔ/F&����ɘy���<�� ����H��m"p��ycj텵Ég�d��gn|�Ҋv���i��o���į��F��gZe]i��i���m�`�?�)���$'E#�@���%��ɧR�=��L�d��4=��S�G5g�,I�M���'_�.�(�U����g��O��� ..rd��hjӋ�-?��$��v��>�w�s
��BJ�2���+S�yCB����H�u���F���y��9x��Fٮ�
�(�V�|&l�8+m21嵍8Ϧ��8�rS���{Jځ�c�{�������X6ʃ����v4�,S�pȭ�4a��$��4�a�R��}��pzz4o\v$N
����{Y[ ��`�qQ���I��{��{�SR������ă��b+J'4Ip����z�B����\�
�.Ghx3��]D5$)���]�'0���(��[�=�I(X��O�{�,��p�J��������|�g��[��:_�P�R��@�pC�o����_x���韂�����q��E)����p��)�*2�0\�IpX�/�]Ƹ�L�!���*�݅��W~U3rv���"�5@�QN��ir�g:sC �`_�Sx���b���3�a��yPt*�!}��3���W�뗑������8H�,��*~kI*�f�:�'è�G�	�̚��@:��� 1�%�y�d�D�g��@*�C��*y(MF��M� ���8O1����H]A;͗��T_[UV��HC�I����i��勉`}�Ӏ{��^�],��h
<�`5|[�z~�W?o~����^�����C
�E~�vo������x�?�E�~	]���E'����Cp�����j������Tj��vkEϩ��5���r�� #cQ��؂kS�iP;$=�zU�o��
�lN�$)��	@�Z3m�MM��\��{ml��a'�7�P[0R.�ω��5�S'�R%�RT�Z$[���X�lD V�n1?�Y�ض��5�rQ�v*�|����`)�и�����k��uW�s�_D�0<���n�������k������\��8C���^r�^ِ 9M�B��u���V���r�����s��#�QpN�;
�qQ���u|7ɐL.�%�,����6h.�c0���7Ӈb#Ň��Yn�>/��C]VT��0�~��hJ���&�]pj=J/:�?+�M�gVI������;����a$M3S�/����J��.q�}�N8��=w�. �(2�Ra�/�= ����L�p�SZp�m 	�PR��!�R:��c!�6���1<
�A�lq�
sy ��&c��m��4����M����)��ZUo\��'�`������F�=��v����5IT[�޾����9�����=(*(���8�]N����U)�����j4&��&�K���e.���b0q|��'.����:��U/��^��u#�˱����g����?�Z����>���30�M���x!x˫s��o8?��^��G�yN����uWIsQn�7i.�}*��כ�ұ��oo�ѹ��)�םT���d�f8�CO7�=u�'�-]�Pxm���4��g�c��9<0���L�y���l�Ks�z�\')w�ȦQ��}~,�q�j����c��$��u��gK'�^��<w&*�'P4���'+�� ��7�O�"�e�r
���*�����
�t�A|����`CK�p�Q��w��k�L)�v��]�Ov�A������>'���ý�c'lXT�g��u{��U�T���_�o{���Ր~��Z}'���z	�y���C��x���w�������6��\�=cߙ-��\��ɫ=Ȝ@|�)�`��~V]��>���vQ�A'e�?Up)�epZd��.Tt��(6��s}�ꚪ�nv&5=s5E'�]L9(�va�*q8̙�F;#�U���,����Ms0�
^����l�=��S0M�ٴ�$W�i�]-����R��b~r!�o�\4�`#�Q[#p�|�f���˳����e��w�����g��x ?|�<�B�nn��˯>���.�pq+|Y�Z�YV��Jg�ze���Q���5a�+T�Đ��E?f���BE�b���j5�[�g҉$	�b�
t��z���]�Ǎ�S*:v��m�n���W`����֓*�uI�4d�ˤ�íWf�>NIf$N�-�LsE��)��z�MiN��|&������\�N���V��/��n�u�.،�įQ�������c�p�k�:�y��U�\�G�E?�"���UE9�L���^��:K4���������
��E�oV&'��������i�V�ۮ}�z`�8������ P}���<���xX��yQ2m�g�n	k[�l0[<�O�������]��k]��K<IVI89�L���a�%}����A�&�Rz��������%�Ws�/q��@h��D��� ���~��^�7�<�\�kT��ң��J`�!���(��7�	>��w�bP zX����a�v}�)�h�� ��$&�	��r��A����7=��ӆ�����ߒ�[@�Ǿ��)!��ZSd��l��/C�m�K���o_���q3����G�/�`��p�̧��T�3�a�򁖟���l:�O�����s���`Yۻ[;#� K��'&�e�h$�9���M�m�	�쩯�L��������.���d �
���ʅ c�9H[�yE��+���Ѿ	��HC4��f�T?��)T։p�yt��<'�P9���:O�B�=H+����$u }D��vj�yHɹ:y]�Pk�иB4���p�:J{�����?����~�렃����p�j�c\�X���-��W?�y�/~.��2��t��28wE�u��F�Zt/tB�X�qYi�u��̘�oP&��Z�����l����1���y��Q!�em'pT�� `_vbG4 �E�-�Ү۰ǻ�mMv�5�F"}���1�U&�I*g��A��C���ܡĝ�{��-0�~v�I4�0��W�m[َ���q9	�Y��K�Y	��<�!g�6{���e8�����뺩�$���>�����<��Z�@�	�oҠ�!�R�>��i���*�Ha�m��;ˇ��t���Ύ���V��g}!
|��*#���[b(v�f����P)`����=�ҫ���������A�0��(�C�N�4G	���dߛp��J%r,O[��Tn��Y�x�d���G"�e��m��4���&p��F�
�a�8���A{<�t���}{���b޾PD���b�G�AK�@RJ�i���S;^�_�"���o����F��MQ|ߋ�����Ł�
¡��+ػ�S̄��m�����є�#���魛DQ��5ƮZ�M'$�FD!˪*=X����j�l� 5�^a�5���3�����br|��p}�������TS�׭��E�������_�_�����j��S��B1�}������^o�/�;�� >����LOylxD?E��	�~wBA m�y�S��T�;
�Y�sn��
6�ܛh7+m�>vr�&Ɠe�9p��k��A�����5�ƅ�x_���;���p#�X{�zi�+~�^���1������.噧Q�s*����:�.j�F#��g� <�(�7�'�@� #���	H{f�v���l1�v�:�,��I��}&�㐲�GE��%��7�"^:�ź�p@:��u �r�l(��*� V�|�j��?{|�K_�~�#C�A߉�+�tF���C���_���������7U.�1���K��PHOii�R���v^DpD=�XD3A*��.ԃن�L�I�7t�3̃�n:Gv�-vx���=���+��a2����;5[�L���dV�P���O�ǣ��4�ϖ�g;�ǽ6��^��aj9�F|T�d:���H��T	�o�N�d/�>K�M>��cR��WZy��7eFIh�]w�N��燄֋�5�t��a��E�ga��������h^�Lp�Xܽ�n��X�
���$��w��՜;˱(��kV���7N�V8ʦ��k�z"&�����Fz��0y��dE�'J@��w�'�C�l���z/A��9ߔ��W7��ڐ���B��ן �[��^�ңZ9,\+�M����9�����a܋4��:m���&q/ &O��_S�vw[nʸ��3���S-L��;��f���K&�E��<W��a�U�{'֗3k��6�m��Rn�r���Sw�C����8 �֙p��a��2��E}R��*/~7�FM|�y�h�ٿ�SD9�v�pD#Р���h�ՒgBQwHsi�Q�-H		��W�Lͱ��*Pv�}?b�2x0w܇��ѳH	���'�;������x9��OƠc��#Z�=���)�n���7�>�#�|z}����D�����zz;':[�#��
������!�Q����C1�c�7?�5Ve�y���_n�����Mvm�p����T�+ds�OaL�M(�`u��'g2tm��㙺�p�O|�O���v�.�#��x2�P>�����xOvo�=g�$oA{	0>��W�1�Wz�vHW��4���<�=��C�]�7�=�_�J$�#NY�l��&�9|���Ө�].�@�o��E��]܆O<~	������_��p;�G�'�J�7A�#���υ���5���eX���.�[D\:�{���rc�kʡ~S�4��w��v�=@K������\?D~�#urf� h��-i��3�篈(�Ƕ],�S���������$��)�[|%��j��3��8o�8�4I�th�ow»��,'�I�E;N��)�+�,SqW�5�����2�(�Ç�N�#��_~#q ��������<�����m�tډ���xGy�,?m�l�?i���e�%&�A1
�:�POܽ,�pWB-ꉤ�1�FǾ���
F,��D��a��l���8䄰��$�T�*,=�������4xz蜔�^������l]T�,������!<�<Œ����`+"�f�j�gc�1���f��$�5u��<���4��-'���f�^mGR�Z;7�M���~q�BFk͸\R,	7�>�rR�L~N��v�G&Ｘ�MJ4��^g3��?���Q�pO��A�͏BU`��1PB�D�����8�N{�N�l�5��h��|W��^}�=��T{�w[n=�e!�s�P����Q��+$���|��J��b��6}0�����oI/�5I�=�>�B���<:l�B(ub�5'�ý�{���N2|����Pݐ�&��~��O�����?}���"n�A�]��� ��S�a�{��{_�m�#?��
���+����a��V:�l��i��ݳ��B�u�����N���8͗7�o�y���/��0GlS��d���('�e�N��aiƜӊD�}��.&߮�3lVo�v��ʝ�|u�3�%7i%�P�B�=3��s��ݫs�:D��u`;=DFl�n=�.���A/���z�:��ZdF+����V�.`���C�9�����u�ꉓ���1虯gH��2�Hy�����oH���mX��y�z�����g/�z��w*���.��x�È޳�z�wNC���dq�������U���}=DǍpE����Ő�/��7��?�Q��/~\�J��/b��G�SصZ4�6ՙ����
r�[���	0�Eա�Ap�M���/��O�G���Aj�M����tⰶU'��~wih^vh�z^��B�d�S�<옸F�Ž�6?ێI�ɸ�D���X��kmX>#�Ct¡�����:v���
IFQ��2��,σ�nl_v��h��[��Nj<P�a��(	F��T��$�O{�����E��A,�{���(Oݺu�di����֩�#�5�H��%��96�`�A�yJ.���&�/Fb��ȩ�v76+Z8���Z����ϛ9�g�D����ȔH��܎sG��E�����a<�N�z�����q���*��./_0%%��q�^�Z��M;8~��xQi������v�]	�?�J{�Pa��DE����aAW�Ѐ� T6-i��q�^�_��@�Kք\o�p�B	i���j�*�/�,����<�t�1�P���g�<�[@l\�_Lt�(��jj���hٶ���E�}�,�<$���{�&������S��6�|�1:H���1q�^��;22y���s{�$��^�4O�v�&׉����;.�<��>�>7�����R(C|1-����$����3��E��x��	��%ς��K/ Xu<��N8T��iW=���~�}�V��u!�#���-Z�=��l��S����ޔ̆aP�jLj>���X,3.7����ոF���� ��<��Y͑��-�7qO�jY�H�W��d^~t���t[H�2&p�é�*����3�a���<��A��{n�^�;זq���?�ߌ\+܂8mNL��~�r�#T�k�ũO���"d���<N:i:�C����^��.B���/ₐ�+�yz_��@(�Σ
���*_�H�����랐��,u�N�;�N��d}ed:h��:L��۟���#F��$��.�{)��}��	�0u��:�\,`5���'<���Nx����p���5��X������O�?��k��?����Sc�P���Z(�t� ��8��h�].+l(J��3/�̡)o���ͤa �HtC��g��0 'd�`e�YM�hћs��3 \�m��܆�D�v��9f��i~�ܦ�V�mӮ?�Tj�7�F�;��ki�('�Qg#��8ST~�;48�a�1��2�Q�${�v�mNC���I���v$�Z�gh��g�$�
{��˔�^�-�S�lߥhͮO�ó�PQ���(�.೾���A�X^D�y�P=s0��὿}9�k���2@�����4����]+�";�=��s#p$�`�hă0����&c�y���o�	p�����s#���j�X���n�q�0�;�۵��"�����?�[Z�[��ߖ��ً9 bTKk�7��!�����q���ݸ�r�W���������;2h�W"|�8P'����Ȣ�28꺤` ��j�;����z��s�9P�#Z՞� Is���{M��w��[̆Vb��@7����w�k޳�:��u`�%�������I>��к��!�E�� �JOBd2�f�)��d���8�T�oޑ��ˣ�6�OXG|�Ŕ���\.�yd؇��v�L�QӳQ0F��e�1�"��_�>�3�~���	���o�۷<��"wf2�����g¿��c?����C\��e�>�y�;�]'��T\N�25�RNs����5o�QI��j�J����3��d�����@G�i�|��C��f��n,���S�j�I~:u��g����;�u��,�/��d`E��Q�턾be!�Ӳo�<�Ӝӓ�ˆv�s��#m|e��6��z�y��x]dvv�(R�>r&��;�7�Q.f:���ӣN���. �bh�#��OI���/U��_:�]�m_�t���ׇ(m��t��=��m�,��{~�̿򊡪UB��ҲH�tXi?��c�_z?��g�p�g��VI��Zn��=R�����N�3�����W3�l
�ub�i ؎7�F��R��@�F�W�;n:��k;�k��C륀]�Џ����?�}����I�)M{պ`�8L�^�9o9@�$�{9S��f�ظ��+w�>aA[J�3l��x�_���<��Jy�Q��=\�t���t/��A��_L��_��9]�ʅ�h=�:9�G�u�//a1�?��F��Wsh�/@n觕��Ҁ��:^`�G�hZ���|+��M8F@����+�J��8c�8́9\oSUf=�2��u �Q(����N�X>Syc(��k[i�r5(�Bwɰ���YkGfl�0�/��X�e� ��o4����W�YjӜ����<�6h�{���)#K
/dhX�Z�#��HX��N0���`��z'@!䦌���i� �O�7<�tj��V��`~����=O�F6�|af�w���\ݯ��e��� ���'0�~��(	���c����r}6�D��W�g8��QU;�c���v^T-U�М���7��E�h��WC_��hk7��h<n��
������]�����/˕����_ű
��`�\�;x�k����;?�q��sCq����8�j��țbp4M����u�)��������3��:�����ȱ< �F��=������b8���7I<��p�{���#v�CCaUP:
�	��K�)��P/%��9�Q�`[�V����F�r%�܈ά��`���N�{���!��*�2|�;v9�E�z��g��!t��k��~òz��t4�9�Ջ
�D�+�2Y9u�0;8��85����m�Ϥ��0F���>Gw[_�g.=���~ ���/���c}�y��5%�u�y�|=��G�?����o��[�9��2D���1��k}�[i��I�`L�a���y�f�����a���pX��u�]X��ОI:���^��FD��6�wFVV�*kw��s�W!�n�4��4���Z�(��p�Я�Y���֯�hT����%e�~
��i�n��ر��)�rt��\Vfq�ѪLcq�v���_Ig'Ւ#��C��E �I0ݢWN�K�ތ�M'A� Α(>�V+p��p�v�#+�pvM/*"Y����PIn��%s`n���&M��n\A�p��z�W�u�\ ��(�v�������Ay�(�"�x�ţ��y���P̢� �<;t�H�uw�S���X�I��pj���iV�Ik-3Ә�(^�q�\)�W	�m�6���0�P�M���S��p/����q���6{���U��u:��
>g�J�;�D���pe	#�kc}_���&\���m��E��6'~�+7,a�Z	�$�3 }	u%���:�����x�I��#��]u��x��XW����3�G'��/	����FF��kYb����
�x	�qc���
��r9Ls�e�`�X0Ćv{1��/�d���?]���x�!�6�;�\�y�G�7T������%�����<���G�d[l;M�:�P��<�-����?��~�{^D�q|�-Ȍ9���&9������84���ޖ���-�ST���8���������j
P�B%9����/,���pꎧ��g7/���p��ӦuG�����X<�T+�y���;�k�n@�l, �A$���ႎ"�Nc��_����ڐ�ʩa�����+I��#)�Z�u��AOp����)�E7�C}�͑'|�'5�F�蒾)�4>�Ggr��Lˑ���|�3崀�B�E/Y��FЧ\�}�ؗ�O-�}�E�h5����‬܍��"���_/��?�qx篼��^q�(i;Ǘ��X%C����/��}��'��~X>��ЇevXJo�z'��	zb�k/�d=�uvi�j�5�����B\i�5��3<�4P��6��";I�d4���e�9nP�@��3�t7��R�Lh�΍���i`�
���;��m�Z�����2���K\y�r'������L����a9�]ٺę�ý ��0~@�i'���?�=�3^iwl@�f\�� �E^�Ҳq������J^�W�%,�1o�{�"[�!������59pXz[���ADbC����Aטc62�\��<���A80�6��
�#ٹ��k��m���Գ�4���YIr�m4u�ȹ�B{�֛��S]�:��Ie�=E����v��M����M��RmfC���X�J��>�i��4�`SZ�1V�|�'�����.����U��4� 	>���-��#����6:<8��E����◸����� ���1�bn�o_�A�T_<�鰯5Ts$E]7�����S�+%��63��K~�B$}s3D��_�rY��b���K��U�=�.Eۈ?�!_�h���\_�E��ox�|�S�g<�)���A`�u����-���$A��	K�hF�?a+|*(��t�o/�d%0y�	m��-��Fw"�|�k�TGb���#�Wc���P�;��%Ûh+r.�kÃ/~�	���� ���<}y�dWU�N$�>�A�v�/?��>�������
�[�6�Y875ፔIZ8č����d�["�]f��:[Wc��s�y�����m{ؽ��m�O94{�Ó�~u}ī�]*K����@݄e�P���A��N�c������)��2�2R�ubӊ�a�Y��	�)����@؂"J�	� #�Ȧ��� ��e'���Ė�����m`��YVV�&�iC,|yͩs�,��!�88��R)�<���{#+��u��X�k|���,L9Ų`H��d����#�5��å� w�ãK����g>�4x������-�X��`�t��A��p;�^�Q����\r�OzG�ҷ�����-��,����u�l�L>� �:�i��4�fԈz�Ǹ?^;�t�~'}(h-��:�U���|��W�Z�����|��%�!�C���4�6��Ý!���1����Q����<�����Tց{Y_d��upiSQJץW�T��=U���]Ҝ�숿1JO���;��Y�?��M�7�{��w[�,��T��v&�%2T�
�S��q�38�7�η;�0�0Rnc����?%m2~��k?����1�ĸ�59wH�K^#�,%-S�\Nu�6yMs���"N'���s�,+�3i[A�)?3�ϤP����(��|�c�"p��8Zt��g��Ђ�/�e�}*ʥ��R$�._����ٞ_u���;1�!�ݻwa�^���E��Q�N�O����S�xHw롷���8\7����7)B��!����E�+��' *�*<� 2j�Մ����G+��|�2���X��o��i�u��H(=��tHm��A�7���_''�#�G�z
ϩ������q��1�L=�U9�ȣ��r�e�`pQ� �2i�&S�]��L���5юw���݌�r��c�]W`�9��+�c��~NpL\k�2#�+�Ls�DA��d6C��X�>��*�����a��׻��;$h�C�n�A4��oi@f}�C��:l�$#l�T��h�95F�1�y~�毂��m�5�ڽnI�0M��	��b��o�-���\ApfX������w��y����6x�3�ݺ��,��F(���{��`G��%@t7:bƷ���!�v���Px��AX/���4i���G˦�!Sz��B���"g@�&��k�A�#:D�X�+�<ܹ탰�^�y�׼ϑ8�>��n�u���|����< >^Os�����]�5OKĕY��T��f�ƀ�|�L�)�<nL���Ł�5�]x�>�X�5��W���>[.��~A��g������\+�ބ�[ƌ!��z�Ħ�z�iC�Z��:��9���cP[s�5T[�����!�����v/8����3�(g9v ��h��
%^�id��"e�}��=`��	��\�y*��FɃl>��8\�7aК�M:��$l@�Ov�G�8BԽ�<��^�*�����I����\,�n�0�>��<v�.��c`t�NDt"���ȃb�Q����Wd���� ��-�"�e��#���#D#���Val�p�V�U%9�'������A���w�������G?����t�����Ѻ�& [�\ �Y�>@gN����N�	�ە��l��g5^P�75GA��~����<���^��^�Z�#��^(�O��6v��\�-9�8S�l�h��������q72��LZ�� �9O�_=o�!1i^���u���y�"�E���Ds������ ��s�T
i1k�����/�y�쫨R��>o�q��A�<�r� ��]0�SZe5g$b�\����s+�/m5�܆v|av���,O(�[�ף D�$�dۥ3R싰���x�S��<�ek�Ko��+�t5f��Lk;���[<B���c#�x�+W�z�JqJ�>�u�1��,7~��Q�P��e�o�)�aЃ��TA���)"�FI2��pK�QX�i�^��	��������7:�N�{O�
	<o}*���I[���m`�B�2�V�u�+/���o(dHh�*C��V$v"O�P����wկ
>T���N$�1�'S�ZT�b��w�.*��F��2+�����T�q������soS{h���N���#�PRy}@^O�@q_��4�ǧ��� �aw�}�|_
��Kj�M	N�%���')$90O�M�uK���z�{�.2�I��w�!#�9�B�5��������������K�$!���-<��,쮓�ClĦ�骑p���ND���a���x�Cʏ��W��gH]#�ˆRX�*�f��4��ᱽUNK��)b�a��7΢�I���7_�j[e��WX�!�W6:�Z�w��q��K^���w����t�L���b�c�����3�ɺ����k
��|
9w��Wٶ��)}:}b���$s�0��o����h��\mD��G&PdH��|6��^ᜥu�5��g�ʍR:n��}���8�$�k�L�g�i��s��@�33�?�o����
���v[�i
X��@���G���5Y���rY'l��f�� l:�/-.��Cr}��`!�$�J��V�:U�"%���/�}��x3<��C7��I;�(�-?�� ��h����D{Р[��Q u�T]�m)�a�~�q0���Jl>
�Z��s�����d�\k�E�����k��ש�[C��eH\��m��k	��ѐ�_���U�y8b��/�m���/�7������ܽ����+^ ٍ�P(�=�f1�����9�r�ye��֦�B\�ԷZ0W��zt� �Sp���=vO{�'�e�
�$;��tN��t*����5/��lk;�s��ɽӴ��)�~͈H)r;ٙi�:�m��\�'ϗdݽ����8�:v�~T�������x��2��]k��(j_<�9�-}c�X\���<n�V<g�q3�$���:�{?���1��5^K���4�,�8%TA�#�z%#�2�����9��O��@�����AZi�R�0��Ӏ�ڸ��t��-Ǔ�n�Ǉ�ب��ܙ;�G)��3��֚7+~����Ǉ��)�� `��`�4������p
�c5�5���p��8�V9��kY�p�����_�~ �2��r`pWgr�6`�}�Ih��;�� ����q�y��eSv��a|��}�:X�]pkoz�K������Ѱ�BE,r]�����<�G�Z����|�S���6{��R=�������I��4�<l�Si΋�X>:�����r���0���h�i�a"��.�U}�I��oz��/���I�
�9Pc�c]<�	犮���0KB����Xq����t`��d��-i�6�����3ZW<�I����LJ���мv����df���rMMֱ϶�7������p�p��s����fp�)9��t��=7�:�}H ��4��`t�R?�H�UE� �6sZ��Rg�.)��w)�by�.E����ܭ�r���Aw����[�;^�Bp�_K�-躠.Y³Ӷj�wYC=B���O���a@�+���i�^�z��.u�	���,G@t���}�ܟalb����IY�|(��d=	��@	���oz><��;���
��"���\Ig�ȱ�']�u�[W��XH55�׌�#7�8�l����.�ߪ�$v?@:/� �	x���;u�(:n�c�%�7�غ�ȴ-��Ta_ޅOלhj�Y}kL����|��?չ�2g��æ��;Ս��:����`doµ6��vZ�	��	E�(eǠYīo,z�&\v�$'|�I���䳵�'k�+��	���&@�2P#�a`C�~�`W����`�b!N�g<���}�=�"����xC�D`���4sC�-\�!�-��ejk��Q��W�R�
5o�1�4��9g���uj��^�SƬ�U7�C��#a���s����|��ik�7�� �9G�Xk���1l8L�N)�����%e̴��[�x�S��mQ2Si��Yh�Y.򪀖.}-�8�
89�v����e/�nx_��5 �p&\/��8���)�Pse�����}�[������u�m2T?�8�	ϒ\:Gg�t�4e��ȡ���U�!���˟�<x�W�w�Xv�%���i��U���c*�F��Ķ��*�\�US��uH�|K��y�����ǆ]����_��:K�2���k&
�"�+~_���\2U��$CN����*_{�a.�5����2dmz��r,�c�NS��):�T]eS����m�:h��a��q��SN�o�,daKBo"L�_��'�}��wG_�����(�ɿ�� I��^�S�,U���$x���L*���!�A���~���'?/}�s��V�S��8B�$;�:O�����J$^��e}阡��r9֌:�����g�.-�g�(����R�l��g�*E>����I��i�j���'=^��g��}�)��w�-���-��mjStK�Mi>�K�u�0��-�ۑ�X�l�}�ڙ��z?�4-pT*�H�$��{v�)2P��*d�Ve�Nݞ�ɉ��n��yM�0���~�=����.��zsr�9�H؛΋�B~�<kD�Ջr=v͵;��c�i�W���#�5]��MbW����#��HQ��x�
��&�ㆱ,mO\�4z��t�p!�j�gA�;�d��L�Z�A�	Ĵb�3F�ಹ����nJ_g!���֜;�8x75V�R��li���ka`� �695��)�UDG�5�����˵!���뎡ܜ�;y�o��7�`R��a*����g��g->3���ߖ���0��ǌ�S�i��ױ~ػ�k�vm�ܵ��S�K�w�Ez�j{��s��gg���x��c[�s��,���4,�1��{Pt�P�ZYـR����ɷ���^���;�67[��x����5���h�H5����܁g?�QpWObN��#��d˥z�4�ɦ��"���!v&M�i�>���bj��o�A6�>{U���C6bD�uvbq������u9/����S��K��,x�����%�"Z�$��A]�J9#�[[kb,���y�9����|ĳK�w����-)ŔZ�n,����oL�Zil�@̏}�BLl�7�,@� ��4�N�i�G�6G^���A��-#�*b�)R޷�6=ۤ��������oY��;��Q�kK���Ǟ��o�s�[_+m�<czG�_�z�:�~k�Z��ܾ�����.�mS������úm����Mz�\���mm�F�Uk�A[�����@mN��?�� ��K�Ơ�"�ܡ��e$��7�R[1*�]�d�3���
8�lXgI����:�s��(�J��e���-�B��I��s�����_�9���B��o�/�'�7������Ε8�����������s~��ՏRg	�8>|q��σ����B�0t3��<O���ylW̜��f�ʮ�����^�v�9u(�
�p�um�_٘I3���+��>*�*���/S�jN����..妼�:}�Vï�[�|~h�o����iu<��T����H��j���siI�M���?S�xW��+!Hݠ���w��ZkW~Ǻmz�9>ۂҋ\�d���n�]�\N�}��J�������܎�ې����^��.u���Y��2I�� ���`��s���u9��v!�����U|�Hy����αMT��Wc�_ �*[�$˼6�"Hr`ng:��
���e�*���4>I�+�-5�J9lUcT_���L�
������M���g��k�i����Ơ�4vm�&��	05!k>!m�k��K�c���x��3���1G��"���m2O��q�D5�B�C�ϛp>��%�eS�d�̹��T
}��g�	R�x �}{]��SH	N���P���I��u�G��>�YB��G�܆�{���Nf�o���D,�e!@z���6��'�!w-��;����߼컨�򗣪�KB:'���q�\��iV���E�o�IC��"f~��%<�\���Z�&�l�����߬G��V v���c��(e��i��}�k��v���j�o./�J+l�j6���}���$cZ��O��Sd��ſz0����o�w�gc2�\�c� l�5�_��]�ۦo��X?���̹m{����Z}���is��M��}{ȃ���������k7�5�(Ö	�{�ghy�D�A�f�h".[a��ցH��΀�='�\�K)U=�&��L	i���p�</`2�7<�aX��$������L�nB�M�g����>����4�>U���C/��9���xlD��_�܄��c��%ͤ�(4��,�q~��K�qK��;���9w��>�x�_+5Ǝ���2q��+՗��ms�zriuH�%H�z
���4������0�0�R�� ��;���Aݕ��?�����m�)����>�p
�@,۳,0����И�?v�k���=ڕ��i��2Z����UˁrB�?����[�9��)��n*M�$�M]g�%-���ӭ8P��:֨����0d;��l"J��_<n�w�}�nmݖ67j�Hs*�jn_�� �?�8��}ճM�1��`�����>ֹR2�(����^��L��o��؄ �a"�C�A�FgD�,��
eC������'��PƬl�dA�M���U֍�*#���d��|��WO<�M��2X�2
h�Ū�{/ތ�s�ZD��FW� �o��1���;2���3P���iܑ�*�t�4�N��3���l�؂��b	���u�>;7�5�/W��kk��C�]�+��g�����%���� ����K�hp�8Y���hg��y��c��yjpHY|۱�F_ا>���C�e��kuj���1tĹ��/��ç`ùIP�^��(��j���g�"=��<;��c�@B�#8�f[Sj��W[!CT]�%�0 G�
Q��p�A�f�=)7�!�^�)Ѫ�<&�ēt�uG�}��خR{e�Pt�b$t�SD:�<����vNjeY��r�=�t��{�����3Z;[(�Sg�E_�9KցP��CYp{c�R�Lm���ؤo��o⸹�˛�B^m�+�M�Ő3����&�	c����曎�"�;W�S
l;�dە2M�Bt�רt។W���r@�i��S:���D����V���Y穮�7�o����z�pd���� 7� �5��8T��?�#q�{��]_;�%\%>�j=)Q�D��@�g�F�#[�Ga�g�Z��<k-�Z>��ՏZ��>S�j880kS�[�Vy�
]�Ɣ��m�x�a t�>ҏ�`ʳ�>����S���BY���![��l�*k���Vu���uT�5��G0�R����)x|�|Ư�k2��R=g����F���qQDQM���(��կ]�|����o|@�2h�?]6��cA�xs�����(H�16��։Lh��Gژ��"ˑ�U���)1�a� �?G�0_��"?����hy1!c���O�|����������HG�(.Z�F�z	�]��i��n/�%���YOőA�#�y��м庍�c�Kk=}z�%,�#��`5;C������yN�S�Ž;�:|sZ����G��m}��т��gS����Ю*���z������O|o�/����;�b'lA���d��Z�L��3S�7�~O��3�U~_3{�Q ǋc��Q�uF��E*����r���e�-
��Ed>��G��3!�nB2rI�Y���>�X]ޅ�����A�����n&#]X�JL��t�9�3��-�i��*Kpf��)����<yECL*��y츇J����|y���~�cp��;<��<�qV ���������im�XW}�lC�e�q�e�����<��oQ��## ���̏��Ti�_�sS��z3�<J��YQ�ѩ���#�l5_#j�oad��_�
�z"|���pA���G���Y�xX�,����P �|�ѵ���C���::q�WҐ`��l?�pv��b.3����1yT��-�ļ�&��Bm�f�$y�Q�Q��G�Q�m-ɱ�*��.������6�o�nk�)pqV!��o�ܭ�+���&�zx`���-G%���kwb�ϛ&"�W�Vv����p����sꃵ�Mm�j&[�6�T>kE�갂u���dv����H4ʠm�~n)��<
�u�'cg ×4 �~Kzu|8�!j�:n#����2��Kâ'Y�lK�L�Hsf�B��K��8�hx�㘮��;�
�^;���+����]��|ct2��m��l�Q0��Y&dR!� bՆ�nX���)�CO�V�c��;�(縿䤁|�8
X���v��i[h�.@�P�2=$K-��������_
wAw�중�'GY7�k��K�ȓ���n5�Va�R�W��tb�ӝ�4��ƱC��>��g="�_���s�i_�sh*��w���&p�ݡm��n:��O�b����irb�WNȎ�/���1��$���%� �p^�U���`_2�����Ϧ��&<;&���z'��l�Ok��#j/�ش���8i{L���� ����Ǧv�Y���)w�5�2,ɞp�a��\Sۨ�!�q��L��WE���%n�}�S�����8���Ni�6F�za_pZ���d�(�Ѩ}k@�����೗_�?��#^������+*H���:)X�N�e,����7�]���h}ţ�b��vB����q$� �g���V���pP�rn�������;�L���~y~�]���A���ci��aSv$�ɓނ:Ou�g��)K�j,����)��h��k?k��yl��9���)_&m��-��tē���R�ܗMo"x�����z��3�E��J'��i��"��<�CO�D]T�7�WL)�?x5" �Q~S���ŴR=��A�Ӌ~��8�7C��.�b��z�sAK�m�� ��p�]�4m�:M?0?����u�J;^��*c �L�#���o���nA�z����1�x��C���l���:�kA��ŗqQ�Gv=J[�HU-�j*\=c�0��2�Dc�]w�ǒ����|r�ut8�Ph+�J�ڴpl0
���Ej`��2O7hp&����S$��#p�+-�8�r��uX�Vń��&��o��{��:����X��h�O� n����=o���T�q!�ئ�9��r��BF#^��uY�Be�ð�IQ�4����B)lb'� ٠�T��`���Ia���y:L�^1��>S��JVt���,��Q�H���� ��)��<,�K�@)pr8��8چ�0�B��z�S}K��J� �wgfQjW��Xc�ə��7�~h�@���<Ti=�6���҄�=��.����%�3-$GF^!��P,*b���W
e���ܰ	! 	�w\7���_hLx�oTrQ�Ř!�;�������z�҂���&�H���������w�����~^����˾��.�˻ɨX��1*�Iظ음�]0��}�>��E4�~-h0�VcZ�`�%��e"�T��o���8P.K���T���oG�ׄ�w'�3ޏ�G>��_����qx��>��mX.�����!�����[��ye^v��}�d�Q���r}�;]x��/�Q���ii�ʚ�z�(5R��:w�s�ʣ-�('��_�U=KķҐ��:8$��~�W��N�:ʀ(��ڛ(V�<�O�c'e�����c��Fh#��]�;��Nn[���2����+	cX�y\Tq���Z{�O��D�Y�G�G�`���Z� ��d<2����	(��i��+�<���l^?z��q4C��s��>�o���A�)�1��.�u8�}A����X]��F�Y�(�f[�^5bf���i�H�a=��+��L2�k��f�¿�ʾ5z���΍��p�r��������c�^�o�u�i�MBL�S�/NҘ�>�@*��,D�DW��e�F%�B���dVE�u�v,���t�q��:π㢇/��������O������+$W�T_��A��Qlʓ^lj!���mE����'=��}\�$��UG��6�
V�i�A�y�����!�-dH?h|S�h�����O��/����?_�XB�\j�t��͈���P�eߥ!;':�^�ɣ��or��ME[`[�E����F� ޓ���k;��x�'B�F&r*��]0��u�<Fsΰ|���7>��٫=�"ОA���e��n�,5��4�2+h������j�؟����z\�K��w2����"��h���\�{S<Π�N���E�3%���yf��5����J�ܞ_��*�,ϡ@ �3>�1r����푗�@�(�+ԲǱ��3�����|��JU�2���ln_ސx\�#Z��7�@���H��ƎF7G��R���x�,�R	�����F;/S�?������*|�Q���EQ~sLaޔgS�(�)Ԧ�m������A����Q_��o�.�%����z�1H�W��^�!-JO�2��+�w�'���E���BLJ®����O�?�~�c_͇yT��~T'lDP,����,��N,�<J٨@E�F�-���!��(�S�	���4Zg!L��/85'e��nq<<��2����J�?�9�q=*ؽS1��Y���I�q�<:�avA�s�v���J2_� ���T�3�V��iXt?��Ր��?�����~��������ׅ+?.���z-4�HW.��O��8�����bɕ>������I��r��1J8�|I-��s`��=Jq��.����t�� �宇w}����g���EX?�X�n���;���ɚ� �k@i�:Q��3Yua�) pɣ�j���!�|
��:$Lq��Tv�rx ���`<[�|He��v��gH�v�͓y9��h��r�H+�R[�Q�
��,��_�Q\��g�Ü$��v��)�o�G�*r��c���u���b�9{�n)�ޤk�ϾZG��b]�@�u�z'J�̸Z\�����۲����ʨ��|͹+�dE�ve�]a�Qq&/<,�%�������e��pM棽@�6r�y�e^�#�pm��D
��1�K���)���,�c?�/�|����5�G)lJo�cy��x��?x�'��>������%�~<���T�zm��w�8���R�HN��$ �z�xd=%#+�7���<��B��;Y<�>��I���"��)�Ri���F��Ґ�+�O�������ʯ�燲�÷c1�v�Hv�5�Q����@d~��w�E��Ta�q�*␃����T��Opy]�u߶06|Q^���Ӝ��0���e��K�#�h�u5r:`ݣQ��ES�Q9T��jֱ�Pg�8��2��M�52��}l_ ����IK&��:?Yq�8T���$�5�֠^~����u:u�"zY�e� ����� ��]�'�bT�-�c�Z�����|�f�Km.�\nЌb�n�0ہC��H�����k<��F�9)4fʊ��A��TNr=��ʢn)a7p�U����kVz�A**Ҁ�I����[c��h��<�Z��Jk���exC���F�Q�G�!��9Ϫ�"���8�2/9��MTg0��\�RA.�7��Dk�M�kw�õ��k�ġ�����eVS�$�%��Ԕ��A��ƕ���c�FʊA��`gR�/ʛ�4��5�]<�X�C���V��H���)G����X�������9�G�{?��φ�>���۷��۷���"�M��u+V�X,�Kb�Ic1�m���Ā��gg�|J�^�(X=��0	�]�D:���:!�l�����p�u��U��$��ِ�0dg��vF|��rb�¸c]aO�Y�s��ud}HXg���Y���ry�y�qx����������A �a�|= ���,+J
�f�A��k�[��,��Ծf�hJ�fM�uU�x�d��PJc���a�a>���fTm2۲���,�P8�3�<���&`���6�W�#t
��$ԌY�sD�|������~��i�LIG��������%n�@��1���k�Y�m�qD�i�$'�1ǻ)za��j�*�o6�9szi�W��M�O�ټ�P���:W���<ĺ�#p�cp�:2�Ua�F9��T��@����o������c�[dCx����C��BH�N�E���x ���Oï��'�E��T���=�����ȭ�pg�{.���\j�2:_/��XW�X�~��E�Π#��hl��H�	z���ѯ==c��^�:Fҏd��}\�Iҋ�H�;����9�>��u])�g/ƌ�����%��`�G}�_�����~���-��g>O<x1�W7�;i<"�8OfJ$��X��Y�:zH�Fβh��G��Pc�g84H&��IPk-����O�������V�5��8βg���9��KG�Ĉ>�	_��uo�S]����mjS�=� Z�%��`��e���:��#D��U��Q[3�H({�K�9��VW�H!�X�֟�+JR��P�:�ѭz��	�x�P���ɩcS}ǆ�)��y��>e�a�#�6��×�[D)�y(j�JC����t׬��e�E��e���BJ����0����1�?�@xMd$��9ǁ���=Ď�	�#���K��Z�7߹_�W���d��[�"�?�N^t�+mv��8,�>�i5�{�f�U�n�י����5�>�j*;-��M2V����C�"��Dwn*�� ����I���)	�⤃��t��H�����.����4N�6�#�4O*z���@
;K�cC���[��=��g���{���e�=e�/�����>!`�r(;��ez�k�' 9+d$�.��吶��p��x��zx��Fp�p�?�2�-���0��
u�� NC�:��|��u�{3��ci��Nh�a�c]�窏%�����9Z�~�g�a]��e�w{q;R�.��7�G�����"ф�B2z�du�nɲ��#��9:�U^�K?������F��=At�Cc�����u�𷫌����;G��p�y�G�x�"0��8�(���'=@�����uV�(��ˡ��K�r%���E?�S�sgeq0�!eX��sf�1:@!�#	�N�y�_�����R�x����@օ$e���*�-���P�@̝�'�cb���AWܐ�%1?RWa}L�4gm#]M��ep�h-�����X��vK���e$0�>�������kN+��u�MV�@����,�U�o�'��ő�2���B��p�m�$�(y���R^���X�����hϠ�D~U�&��
i�iS�`×���ju�;��|	>����|���_����>�7n��X.Q7�p��ċO�{��~u�ܻx-��G*�>K�Y���ʣށr@�Cx��:���KW��g!FHp���n}���Zd�)��['�l�u�T�yr!]�����O��B#����?�
VCG.�Up�/�=r�%M��N��$��B	:���e4��F�9��ȵj��^����F�(�@���){]�ݟ���������|݆ߧ��R�,�ͣ��z34`�{���HBO���m��:�*g���ll�N������s�ͪ��d���r��Jj�_��^K�}��Ź
~��G�,l�����X�#z�~��|,��t�v��7��>;��1
]�WhgG�Vd���(i��l��*�6�:��X����x���z6@��hҁÓA'Oh�|D?�WA�~��#���]�PV��5�TSIX�ؖ֒��P��b��g ��F��ZH��(މM���'I�}6�y��������z�.�w�7��+�d��������V(�F��aWKͫb}iѾO�+�*��~���u�Ķ��q���V07��M�a���q9�ࢌ੿db1�^��u�p��2�2/�lAb&����7�qhd����Ř���C&��"z��NQfaX⼴4B�����z_�k���I{4�����c�'�C�cБ ��|P��p�N��������ǻ!g�.3�.��w�p����<�h�R�5��þq%5]�2�$?e�)2VиJ�?ל�Ƿ���y\���N�p��&�g�e��.9�t��|��\�/��&=����Nn�[h�K��X�h"=�cC]�~��`.�~`"��c�H������ʒN]��N�?88oP4�D�P���k.w].G=�{Q�u0z�h�Z�P� ��Jm��P���ŉ�y-���,n?KC�W��d�X�Ρ��m�4'��2��{�!3��7uI�7��g*��'��T��X!w�>V��sd��]�.\ϋ ��z�o��	P/��$-���kz�����C�2�q3sՉ�5�l��ߤ�X�6����;�:��>�z�� �w�>~�`� ~P(dA� �M&�Ie���=�:Mʸ��K�\��9�N��8�(�%E�tHJ[��4��7��etdXY��%������p���N���`�����}']����^�S:P�~��l�8]�Q��<M
٩�+W��?X�q2.�����I�O>9���:���W1�{c���(�_.S:Q2[�Ÿ�2����A�T0D^j����e
��5�6��~����!t;�+��a���v&�����K�gLu��{M�*��[|
D���a�ml��d�	h/ؤm��&�rN?���g=��S�٤_���:�y��h:�W��C��0�g��ma�q�#m��\#k;I$L }�.䎖�Ty6���8�Q�[Su�ķ}tJ�{�[';nh�w1pEO�R$h]l�F��#D�X޺H��Q�ς���Hl�v����Y����Io3
�q���o�
U��{m�6O�����Dn3A<�hAE�8T�'�]3H��k�QOM�m����砲iOT뚹�NQ���)���0�\V���X*���0[�QV�8y�i�<���7f�\�L��B1̏咗��Rq�mT6	�)Z���J\h�ᩄU>��Fs�p	�.��2�Q�]�H��a������F���8R�s)XQ������ v��i�@�Ҁ�jxr�I�;�r2]0�[л��(҆�o'�h"ś�8?�7�@�ASOG�ElC5�"�V���|u�Z�9;�d���[M&����K��!�mG{�6�Q"�������1��p�t� ��wb���B��c�}ս}��;�߻�z���X�i��N-���F`E�V�FY���qLr�1a�N�>�^6�!�P��
0�� O� `���1 m[��K��YY!W�7(<g����N���/�+��MFjB�7�6NO��,�����!]�w��"D��c�e�����g�k�fbs���=�����.�Y���f='�ul��:�c��H݇Yjr��{:�пP/�K�G8@�!;k$_R/[�±$;����1j�Uq�{5��?9�Y�b�TEN8�HZ�X´��i�>+T-\;����
��_Dz?���Y�@�Y'O��@�D��:�	��y�}�����Y+����"�=��rT�.p�@k�P�w�N92W}E`(_�`��Aume�m��vlCۆ���7�_�N�^z�ej��Mce�Q;���$�*;��F�Kk~j�>��k}�ԏ�oI�0sF6Q-���|f�#�>aG1���Ζ�5º_B���"Pޜ��c<Ȯ�u���R� 9�N�捛��;�#p����ӟ�B}�3��G�=Zt[�M�w���g�}I-f��?�����$���B�M���
-� Ƭ�+L�5�H�'���m�Ѱ4 �,J�}�m�����W���NnhXm��jP�B�w� �� �������-I}X���s��;�0�	3&����ĐX�N�a�HX�� �(�b)�)R�9�|N�(R��R�LB8q�b0b�y�<2Ø����w�9{u�Z������k�������kuWW��~]��[�:�WH�� s�%��R��X�׎�0�wFw�w(0ҧ�Fv�ee�&�|ǣ��uH��p�F�gۣ�ƅl3$���lsD@WTh���JPS���%$�E]��B�@����ל���c�F�5�G�w�C|I����<�W�d=�y�E��*��T�/n;���i���	I�Hصd��#=���ꉵy�Yi��!�8rQ]�y�R�ĸ��:��<1JY��0-:V5eR���Qw������_�!���0��i�ȣp~r�{�ϟ��G�����w������m��i9��
��=:md�<��fў����8�	��Ŵb��(��P.t���#C�mkji;.F�>�]��fХ��Q���,f�$*�������=�Z���h\�c�b�t���,����w�]t��P{fӑvM�Rۤh���d��6}�|�S��j�3U��2�r�X��ڳ9���[g^_��=~^�,u* t�L��N�����|=m)M9K`Y��|&�Y�>����{�g����/ +R�Q�B�Bp�'�Dկs��)'�ߴ�Ye�Q(
a���ځ5j���s����.� �(��,��O�"3�]x�r�)��M	�	��@`}%Әl(n���;hS�;5(�ƅ��8�]�C���j�a��!��wp	%w܃&���;:y� 9HϺ`�0�Eѡ�A�ZZH0$Dq��X��,g�]>	�p�*�+�8�T���>��!ʐ�;�⊏���Acxj��=M7�u����c�M9n8����)��|�]-������hl�R���1Q���~����1 9��Xix,�Q�F�&-���[ ���Θ�Ŏ�Ś���[< �%ˣ_v�LRo�x��y��]} ��"��9Gg`�/pR�n�JQ���ށ���I�;Z��EI�������ry�쿍'h��vdH:x���+r� 5�n�4��P"�n|������'�7�'oP��S�F�1�-D壓D*�d3��ry�촞��E8���W��{��!t����������Tp�J������4Ak\S�2���%�m�� ����X�=��9Ġ�>/r���S��p���i ey���@\��[l�)g��t+\y��[x�:q���앇K�3S���:���Ey�@RI�>c�'y�k�k��\[PT 16ng�'�㱇�ϟ���]0��kRW[KF���W����D�<Of7٢�@���My���y�׏��C��)���i0�7��L�z�ɎS�~u�1��`|-|.Y~/C�<�L�<�5\7�#��������<�G^��*<� �Mʗuƍ��gЬ����P���.`�}p�ԗ��x&�,��!��'�ǘZ�\o7�v��iU͢�*��xT��|T/F�#~�g��9�&C@v&��5�:P�����g��+sL4S�ވ?J��y('��4��ü�\с��-1+�$Qe��v8�r��&f<�m�(�D��o�1���Xz�nk,R���p�K�U���Z�1rI�� ��g�K͸4�K�D��/�/�fK[`'\߄q	w��촗��^�nI��<�t�2�w���/�݋^�S�D����Sَ(M�҃����/!kp�
�ʇ[�7V�ި:y;3wˏ@��a�A���=�A����'b:�^߅�yN%GfM��n��z��i��m~��3R��&8d��"F,�ux�YI��wJ��sڶ.`m�H���}J�7�-� �H:�w�(�ߘߴi�ʁ�i�������S�r��^�����$S�6+�n�^;-Kg]g���l  �^��������|�p�K�Q��=�6ާO,�9�]��],R��<�Vv�Ԕs;qa��>Y^e!���N�_Kk�kv�R������5���o۴<|{	6n�\���d��,�C%�\V���mmK��~��zV��V>k�\j(�k�h������<ΤcY%�[m����B������oܭț2!����HE ]'7-��%�S8�S���H��D�9�"k������
���2�;�	5�$OŔ	��b�+�����G��զ�����"��<�Hg28��S8��=1�N�K;m�����y4*O�� R[ȮM|2��U�j��Iyjw�՞y|��ś�kJ����Gm�f��j�u-�S�~�m�|,i��Wg�<�����Óm.[&Ե
��\�_nA��22�=��Á����i��E^�8X�� I����%LQZy"�R�[��9����x.�/��a��l�i�2���X��Է���1��D�w��d�A6w��H��9f�%��_;�������N�$^,R�.�Xa��|�i��+�ĹJgI��wr|�� 9�DY4y����}�cΧ�r�.���%w���JO� gΠ2B^��n2��?��6�O��2�mS�#%�]�:����=��r-��<��6-'�;*ϵ+�	m*t�����L�ѻ�J��3OG�a��)O���5֦i���M�6�5yk�S��4����!/S�������05��>����_����v�T۫�Z"�|�ڃ�s�64����
�ř
78��;�x{e(��|BEb�?:zx��Q	ۑ<��nK{LsX���d�C(ڪ+�2Q	gG>�WD�W9:�J�Aֳ���`��$��cǟ�@���H�Ȏ�c��a�D���q�*1��(Z��嗂q��TՍ'��O��w5����w��ӓJ��w��Hc�m2��;����OV�2TOvu	i��3�\�eO,D���j�ۃ��
�Tr�E2P��y�AƯ��q���3ae�9�����^�5Br�˕����<�
��eXZ^���oX�%�i��ʾ���{�9"��	���
$�<��jqjiش�d��?�ޜ~6�o*?Kl����x�䚒y���Z�jv͔���S��t�=hM��+�Z}Nŏ�߮J�Rֽ�l�v��g�kژ%�'w�w�{��bZ� N>
I�qrZJ�3�0�����o�K��+���`�n��:pX1�Sp�lG�Lma)�ki��<�d�{S��gזi�-{2��z>Bf�
E�<�
�ޠ���r��Q�!cu�@9U��@q�Jck~��-Ě3��#I� ���29g�+0B6v�16_ҹF��Y|x���ʗLS���C]��v� 5.+ IF �&$ 01`���>a �(��<��v&ۇ��6,K��.� �c�����H�p y�	OLe�Ն�GI=.qÌ<M�櫗�:��s���S�+䣉s��R벚လ;�G�x0�E�����
Ƽ���������T��Fc�s���jW�7:�b�,!��-:�Z���P��/9O�����l9�@%,�������ד����%ac�Xk�����=hm{��p�[��%�{|P&k��l�%2n��\�b]������y��íuf�si��xs���W-m7P�s��Z��!�;�2,��F@{��8���[A��V�4�/��L�\��EEa�CF:k�JJ�0}�n�v������2C��1��-����Ot����Ar`��-�6�%_7�J`�`ޕ��b*�V�l�\_t�E�wt��eH�t��y�E�3���L�c��F�|�2.
��V ��xbR��p�
�+�ݱ������R��O�>NJ������T�gj�'�Qz�4��b�:�����΢���3�/N{Mvy������ĦX+��O=�z��k�ݛ����u�sd���j��g�-�u�$oS�TN�B:�Nf�Q��н�����C� ���!�1p!~�����I�nHg�G�%̼ڻ��X���+���I�1ޟ�u��K�d�M���b�̦&��0�࿱^l��/��JsI굼��yE����|�M#<p�����F|����iQ�u��C�A���uch�Ns%c���m���$���(�/*���2�'>JJ��c`�N�c�W���KK�{E:
���u�x/��2ȅ��6���oF$Q
�~��G�^kP�ɠ�A׫��sL?3#py�s0�V��oi��*�
I�0c�E���y(?3�9���&����˲��~]�Mך3pw�]��\� 8Ǥ1!�~�x�q�s'�k�H��iΝ^�.yE�f/�|I{�[m�%�O���<K��xo�E��3o�&Yn^�.\Q��o70=���fm<?�J�e�^:g�y˃����5�o�i@���:J�E �@�FS�_Ѳ)��+��H�\G���p:	aU`��yA"pa�(�B#� -�e���g��dS�nW��kVDSo2N��7i��v0L�9�B�OZ��@��&*hc�C�Y�F
R/��c�T]�y"�-
=q� $���H�]�W��;�^T
��7n��z5g
��ɶ1�Y��F/) 
���}<nCX��6�LP���|�Vw�Vw6�F~i��%�רǳ��1���a�Ǹ������(����1eRh�9=Q�aY�E�ɉj�GE�$�Q3y����@�|5�F{M:z����hvE#�+%�F��%xg��x�z��N��e^+*!��䢭IF.�S�Et�U:s�Æ@�L��Ve��v������D�ъ�E�d�O��)�]g���\����!� �w�)�� ���z�s�X�9�ז(E�%:�d��*^yz�P%�Y��c�9*����m}Ƴ�m���m����k��q���}���Zl2 �}�Y6(�ka���h\]k��+�f�4j�0t��5���.�Ν|�,�h>gB_q��[�>,��DW]t�0��Yyt�Š��
e0+A� ��n�/��1P�8��Bล�c�z��N�F�y���W|�Zˈ�f6�ɉ py*�&?gok�_�M�֑��;dgQ�ܷs]�ɣ�w2㊗�Gj²ٶ�o�z O5�����桝�p�������P����>l��oZۯ��}/�)�n��w���d��(`[�?C(ƶ�;�$��Y}������:����a�<������S��y����z"�D^�n;�
b� ��f ,����խ���y�,�.�O�W�
]�9�\ ��P���i�&t� �'�p1�mRפ&�(��6oE=��b������7��G����]]u�7�oT�c:�3�w��m�rA���ӍJ�>^��U'��i�K�ͼs9w2�W�sG��p���r�#��a׀%Sr��,ɇ�6�
�h�e}N_j���;�Ζʱt��T�^�g��o�@ce������0����I�u�J��x���$�U['E8��=��;�7�A�|.���X8�Fk�!o����4:����Q�$'�`��+�ϭR��)�-�RA1�*k*sJ�O W[C���T�� ��L���27�`L��辑�E�_��]�J�A~	A*� +��HJ�!��oѮT}f����L���_S~K��ñl��5��5;��>���@u�׫��	sz�\��S:O1]�����������@�K��KP� �'2kSx:=���h�,�)>S6�=m���{���Y�@�%�s��>v�KK�K޻aGƷX�7���9�Β�̔ǖ!��H��g�.��:$m�!Oǘ���K��3F困F8��^�E�+d�2��xȈo<�F�4� �3��[ 5dYK���C����Y���\b��p1'"�Eo	���z��'$#��6����,�'�TFC�!s�v��(X��x]0�+,�2�x��q�!�-�Q\�I�_.+�9rB�z�P��B�3t9�vF�0<��|В�%L�+(@7�9�!B(���[Dh�)�z|�|;'�OǴ��/:AQ�Z'�$M�W�a�xb�X47Rw�}U�	1=!ֹ���c"jlű��z���|�2�);}���Ey�m�yM�cc���R���h�M~��pK֊ja<�q��'O��T�)�b�B���Tz�*�L��yn��>��N�^��?ȇŗc�L����L>����W,���q)��S��	�R�io��9�p�k;/q��~�g�(��4ʣd餵<�;�L>�T�2f�si	��t�8���<R�`�S�X6a�v���Dy7�j�(����<��)rxiJ%#��,�Ki�I'pf*O50r�>mZ�0s2ɸS�L�&�f�<��i���ҥ��X�(���2����~T@�< �d��d[dP����ҫP�d���x�,r���
p���mX�d�DzY��4l�#� �[q�w�)� wJIs���"YX�h��q�&l$v5 �3O�*U����6��P�<�ᄅ'߉2�.�A����X��q"8�T���*�@���S�2�bO	`�ϋ����
d�=>{��V�U��ҷ��J�=9r￰�g-�I�a�ϭul�[v�{:����^v�>��W$��<���h�v�$^���Q��7�ᗤ��o�?�º��@�oݧk�ZZnٞ�Um&�SC�>^c�]H�ֳ�Ώ�7k�!p\���r���);{���2eV������bE��OC�l�o�m���M�}^��e��D=����l��Q�ec`������k?n�d��(^��O4g�YoQ�A!�gva;I�'�h��J���,�뭡R���BN�u���u?��}���=����;4�_�<���/����iЌ�s��e������b�>�:``���}��|����j�"����L��Y9��	/Ål�?��Px�-�Wr��Fq���50�V�X��z��[h�N]��[���7H��Sն�T��x�aÄ�E��XEn�H��'Ѧ� ��S.��M����@6�Nr4U�x}jh{�v��ǝ�*uo�Oa��vذ�����F��a��撉�6%�+Y��L���,ʶX��}>@ra�%{v�s;е?Mg8p$�<x6�c�T��WV$�s�I�)0tɻ-a�ʵ$~���h�R�{����{wn۝z��/�3m���k�8��v-�P�n�(=���z�����z���[Z�tdJ��l4�F���H3�T�a�7aQ��5 Q���Q�yC#�7�i����}'��4آ�0UP�E�WP�:��ƿ, e��d�rJ�b���I'��L(���r&$�B�����5��j+���\���p�F�*Z��4<g"�y1m?l(�k:
�=}/�{/}j���D�5|��t��Qs�؃�;��G�5�'(*8�X�[�����P�}f+Fꑊp/F���+Jm5��3N�4�x&��eE�ˬNG���c�"I�/2'�[TMH�ڃֳy�3%�DîV��Dq�+ܐF���^\���1�4�����8���i��3�6m"�w����K�F�#��������b�a�v56���SN����"�|_[ԔϽ86nM�)�s❢YgZ9��8sy�K���Y� <}:d�ϒ:S�3��˟����|�w�Ad*�)D�I�9�D���ʁ�<�����-{�O�g��������t>��-�3+�V�x�&��?�� �Gz��<���s��֏�$F��֥Q��j}��E����8R�p�V�"��ŵ�@�F�5ZG[�Q��7f	|���
�Ji�������P�!+>B�5 �Ay�q���2�Ĺ,�%æ����N�����plxށ��w�svz���L!��z��U�ʩ`�dfm�~����
�����Ѳ'��3@2�p�A���iC�rL��OU�:Uvv�y- �2��r��4@�*���૷'��P�qy`_�^I��_<� �}8����Q�F����ҒE�9�;^���/3�n�?��m��x��!+
��*��~����d褣���G�!'� ���-����ס!z\𠼦������B�	��=�,@5��l.�`�o�{�nwi����ü��,S�S˓ز���w"*�(�9�gY�k�8�t'�۠�7�u`i4OC���T;|����=���ڕ�.����Y��9��p��.��x2�M�Y�#�-ѷ��W�G%�^^�򱄏f	�2����YRg�P�N��jQx*WL$&���3��Ȉu��]_�xg--�fjm�V�^�ܼTc��2ӧ`�>��c�<��jޮN,C�u4�)0��'��kF��糆���";�	f�op��Ӗ�J^s^i��D0_-�L�1z�?T��!ήF\�_sw�R�TCmԨ�c�R��[RM>�)9|�4�n��N��A}�zJ�$2 �c�x%� ��@m���Q�1��Ƈس:��ك� �z����$\�5��U�b[���h��3eU��x`�09�l08b9 =0x��8���T?����Ĺ� �[lP����'�+�H�H�$��O� c*� TܠeT�Ѕ��-�)�X��w�u}� /A�ڲ�;:{j �i�bpx[�'����5 ��d��ɇ�3�<��T6;[�+(�|�no'Ȓx��l}��1���4j��|��a����gk�)����I�l;�rގ��`g���f]���,+������<o�� �^b����-�����^:�CY"���¾a;���{�Jk�����@z5�N�Q�S�O�t��1X/v,&'d�S^ǘ���sd�jc#wb</����o5���,��I	���<�.T4�TG|!�7Q��E!Z�4@�gQ<�za��֑JY���ݲD��I��a�;�=�/�_FaLRtpyh��;jw���� ���cb��G��7��b���IAE#����tEA�X[�	 ��̀�����(*��T��/��dxv�
�K��-��|��"/�P��|8�g#�k6��WL9fXy��N^>j�l�a�d�n.���oYj*��|�������H�j�u`੹�-ڢ��|eg�gJ!��OM�3�Ӗ+���h��4�fj�%����piL�ôBw�����8_v.��6"��'#����
���3հ����=����טW.i���"�_!��pi�G�F�5�z?1��fl5ͣ�`N�Qb.ֲ�M��V*zV�_�ĝ�REo���N�(<�hVoP�FG� �T��֠��W��H���g~) 
�piل�c� �bʆ�Z�͙�3�B�����ĕ�+ �K��i�~��p����2Bfe5<m����z�J�tđ��"+����lQ���Du�Q�6ˎ݋������TOC.[�z|T F}C��[ٞC�e�?��ڨQ��Py�E�{,fN>m�ظ��%
F/:��Z^n��NXNl��D���ư��u��6��S��T��:�A��n�'a2�}��G�/2���,������&/`���A\@�+3��I�۱y���8罥B^,���<�CQ���l{�P���J/������:k��f��!SA�i��p�Z�i࢛Xd,`^]
��Ʊ.��[�2���δ��M�ff/$˝�t"��Uק�<��Qv����O'�:�O��9�N%���ԁ�.T�HcLt�8=C>J|1�)<����̇�+�RK�m>�ȑ�D(ۑ(�)��%x�u��?�g^�Z+Ü���NuZ��P���~b%p����2���Nyx���B�1���|�:	���"Dc�SN=��Q(~��]EۘkW����"��)�Os1�N���!96�������ͭ�mR��W�U��a��y��W��v���G��V�n�P��q!z���G��Q�F�S��[��Vc��t�W�v�9^Q��WXغ���ۇ2����-�(�!Z\)"A�h�g�R�CBTr�?C����u�GiyB�#�9�,Th�A�嘴���>&��E�L0���A�)4&�q�s�}��,+�-F� Ծ��lJ�xD���mM� � ���W�5ҧ�ɀ�/@�7&Q����m(�B��B!�L~WV2t�����0u�%Ʀ=桩]w�y�)N�t5��W��X��G�h������~��i����f���K��m<������k�Ii�'����g��7�F�*02��6	�+ˇp��j��c�}�'����]n��\	)�ą�g��8.�Щ/!]{>�;`��z��.jIr��u�AO+:e�F�h��N �K]�m�eF�YZ�R�(>�]^���y� A$��#!�������,���$�˻�k��8 �ϏB.�6�MKJ�X��3�� )u�`Ƣ��:��9���@�4�������/*|,���G(ƫ�����| ��R�M�&��=�=�a���-'�X�N��tX��N>O	N�3�V%M��Nbk�hs[����Ś\r��(��Q�g�����:�N�7p�H��b!�5~8|�z��
���X�ۇ�.TVR#+h�G;�'9�4ޜâC\8>y=�Q�F�5r(����5_�� z��F�2J���%G�`*]Q+�<�Ω����ROߟ�$*�B��#���Y�%erT���>����r��F��>����]�.��p1p�r���(r;��E����2�V� 9�D�=�@�IuT���
l�)�.h`B֬�2R<̧2ޢ�F���p �'5��%����^�=/��Tfj�j�	��C{��>��x�:�5�{�d�F��Arqn5�}W�|��+:��*�e%�� Y�Ȏ8j�T� �_|�K�T�WJ
ȋ��oUV(*F�|98o�EW_��zD|�Y~z��ե���d�C~;>m�{ҵ�rq/R�r��'��.��Q"d�J%d��3:��y������EZ���H؈�a��9�AԘ�N�5�����<�R^f9S��ZZ˹���#y��ū!�i\���
�!�fv!f�R33�LUaa�L�+���gɻJZS|��U�:�5��M��7Uw��t؅i�g+mn���W�cU�[�7��3XH,nv#̍l�r�B{-L�锧0'��|Y�𒧓lq��t��ڝ���ƅ��s2�P��PG,hԨQ�{'S����[�w6���c�#'�Vr�s!e�Sq ���QE-J>ʝj�$�Q��$���4��u���/;R�,S�Ѷ�y�8Ȟw��~��5O���c<��]����cG�)9`Dt��!�&y��
�9@Q&��/V�̑����Ɏ.�l"�T��
٬,9�	Aw���oW5�^0A��LX�>n�^'��LnE���x�Oq
K夙�~��:�nC�Z~����	�Q�H��l�F��y�<��a�*���,�;t)�=�<H����ځһٚ�k�[N��	D����|�'Tٹ8�Y��vG�+O(G�)�apRG��8�;�����bmx:�G��/�=t�0�;!��Ś��I������E9x���R3�6� b�n/��+�.m�fe�a(��{:db�'
R",�4�d�)�
�
/��S�CJB{�VK��y�sM��&��m41� ��t��W�lv���5j��<8<�}�p�zHV�j1շ-�\R>ޕGۉ�&�'��*b��Y�R�>UqxG�øb�=�q�j緲52��lԨ�=�c��|�ޛ��E�̓!]-q<={��c����%�UK5c�쪦E-���Ӈ�I���s�`͗g��x4n׍G�n��9���$�IN�Ncݧ;2y��DB@1��*�.��h=%>p+�OSL�'5:<)��v�F2@��|��vc~���2���q�]�������
�q�ހgOa�r��'��]	.\��b%�X��+A8c�z�U�3J�T�fg��(��T'u�f �������JE��1U���?y�h�{z�w@W �L&;X��0!�숾k�]�{�^��U?u\�8�7S�~K�C��.�$�����6�t�x<D�<�|�O��;��-k�`�s�-G��ｴ�F��zt���|��WE4^`��9��)kS���v;�)r��E +\�js�%�;�������v�ǠG G�p�I�爆��Ak�r�=&���){Xg��Wb���'$�,C���'{���zN�8��/��4{����=�#O6��a[WUW�C�/P���&v����g+A>F��x1UvK�M�i*��>� W�Á�}L&��C�����&�b�,؂Yj	�i/,�d��[M�����竦�����-�����ɘ�^s����`kԨQ����8��s��A
0��|�8�Wy.8g��N�U��5���B�9م��Y�ʀ��]�|�7<������V�6?Z~5j�h%Y��Q�q1�&u�|�ؗR�]3�M#����9m�0p��ݏ�+�eٚ�T��T������_,cf\*f�U�
i,�T--��[��)#)�㯀W��{��/���`z�w��������� ��	>����o|����k otp<zq��,�p�7���;�s;%�/2�Z)�9���V��*����IƢ����y*/Cl]����&a�N�����}���D�Uԏ� ��_�~�r�~D��<�Q�LG�4���KP��a<���X�Q�RD������.'x�1���`$?�@y;���saYwhԨ��K|��uǧ\��]����2���>t����Gsl����S�C0{��oz��
�$� �-ɵvm/h�z�j��l�Z��:[/Վ,K��!�B�7ⱇwN<�}3��|Y����y�|������g�ӧpp�_�����)�����xL��WP���\%y��6�#DϽ�A�<�OQZ���s�P&hʜ�=��Cx��
%�
��0�vǎĚl�j�;��e5U��Լ��(��#��e�n[�l��c+au�P�bp
��n�Y�:M��b\��/x���!���A:h��#�F���$��H=�3�E��{q�E�:8�{�K$�n:�A�6���+���2��
I[���WZ��,nԨQ���y���g��s '���y^]��4�W}�}�ܙ c}��T	�  "eXB�J�*�F��P
�oÙck\v�����/���߁�}ϻ�������g������롃p�����o~����c��8|�{��g�~��x�: w���A(ʤh��4�{�+Ĵ ��K��_�&rC@��	�t�F`8��Oo+�_U�W ^aU��D��+%�Z�0��8jB��-�y��-I.�LI2�١e_]� ,����Iw5_4jԨ���E�ͼ�����J��O����O�����uF'��z��	��O�mE��!j�5�o��|]t�A�C��z��~G�~x����N߿���ɯ�������_���E�^���p]d������~����O����8����}�=����|r��zi mC>�OoTX��S����R��a�@�	�P�:����{m.�%c��B����^4g�9k2����6����έ�dD%V1µM?��~�X��&iy���̯F��'�a��$��,�a���^3��8l�%εpm*Bչf�`���aZ����_mjńۨQ�F�L�:�cʳ�ܴ$P�SO�8Gf���\�A�{�*&������fJ�\��c��~�5uD{��L���xn����D��K�FC^���(ñ�8��6��} �������ć�� v����fx��#_��5�����;���q�L�l������CZ�pt@��8��c����V����Zr E`�sJ`5��BI�>E#?ϯ�.�{��K�> Z�j�/U�N<x`[	O�;�\b\ i�9��O��ᤡ�.��8�q�e��5j���T�e�����Q�O3ؓ.����ײK�+��~�E�\ZC��
KZ���f�8@,�>1���U_�%G��g��{ң{N1��Ë �{����ʷ��~�w������/^�̡$�{��n�#���#_�5�_���?��߆�����9�y���h�҂�3X9EAD�e��払�SeV�B���x�9�߈q �g��B^��%gc�	�nm�VH6�[����tB��Q7�I
�6.��K`&�.GT;��y��՝�,i�q�eT��7f���b-�s|\����2��ӍnC�u�kB+�N��J������S�gMͥ3�_!_�xI2^�2m��k�y�(Z1��j]�/�����D��߃y�	[�?�n���ݷ�R蠏/�s�`=�5jԨ���:�c���,�^���hT������*h����<��hw`7K� qt)��I@:�X�
x�@����L��(kf��j�|��ma��g���@�w�={�G��E����|�W |��C�s&�+R'�/D��7ބ��/~������ٟ���t}
��u�p�R��xP�GS�fe�ho�g�<��kKW�SC�(*O�He��,d��o��1��H!+�^"��cJ�d�=`{A9x���~l�9��D$�
L3�
`&gqXQ��]�T6r`��B�=j%4+��tQ*vb�E�.�&e������mԨQ#1���IyM����<�@�̓��k:�F�vi��\��8��?�Х��^o㦳!Y4	�6�F:���Z�l�HpY�'ݝ� �D�����E�E�ɱ�k+�����M�;-S��I�co��y��o����w�������1�\4�+%��'�����{�?���K�ċ��?=K��C�C����	-��$��Z���b�K6�,�%�'̾S���1�&*z�TU�N#�8)N鴶^��5el��EG�.8G�:?,���0yl{�|�Ğ����R�!r8�'��3iٯb�}jW�����Yk[wG�15j���uKA�9��=�R�3�'p�k���G���\pM��=W9pX���ߕTx5�ei�p�=Wqh%��`�5j�y`��<la��x���4�3�q�����K�iE�S0��r�s%M���5}�Y��5���i��6
�l%�(�F.���lk([��;�~X(-��{��Q�D���t/�� 8t��;�6|Ç>���^��S2�{a�˥O�b� ot�K���g�ߏ������k��8F��.#���J��{���M��a�^��*AAX�%/��e������TI����K ��L���	D��2�2T@?��q���U�G��ؒx�~�@0��Xl�`Ĺ�n4;o���A���pj�hW��l/���Iͩ|��u�Q���\Д���5j�Hӽ�Os �8Ĭ-��d���s��R̪/j���~$�>6�uܸ�na��D�A�
�0&[�ԁ7�p�J l�꧰G���/��	}�C�I��Su"�E��Y��:E�g�R����_��o����}�68j��Sǘ�ˬ�������?�A����=�_|��g��p<e� �6���;���eOe$mO�څ:x�<`QjR!�2� ��c߬�T�c{�
�}�����rBKh�-�	&�-(=�lP�Z�aB�oQQ�-���Қ%�
���R�#�ѱm�>L$��^����������v���6�6\ �ԇ�G�G{}��m�-Lɪ��Z�[N'��q�R��Kq�?GKO�Y�gi>���ȸ�$�K�[���F2��q�OceNrY:����ei���.c����G۱+��V̦8T�X�u|ͣ������oԨQ�G#k$X�#�:����g��8.���=��o�h�� �.�u
_&ٶ��R�ï���o����r�`�UA}�Q8�k�	���_�v����J��y;��Q! �g���0�U�~/���[�7�֏������N��2x��-���~�i ,?�,�'�T���R"�t^>1B����	\h��W��`�d�.V�e(V�M�'�V#E�փg��b��=�Pq��x�t\����r9P�*50�@��4�t��6�mt����5j�t��Ӕ\C���t�`ޡ6������;٣��E��C�Pk8�c�������B��
�e�d�tNC�33t�n�N;����x�{��w���u �߁�a	�U	ȫz0>;�l�?��~���~
~����(]�ޑ�C��ҕ�(�<WF�;Qo��+&sY��9�U]���*�����F�����i ���P!)�Ue�YK#�x����a���\�:�9x���l�Wޡ#�I�L�A-%k#N����k�1Q��)�05-�0�I�k�8;���B��Z�F�E�nO
���ڰ���0����KdYB����)ז���-h�xW��h�QM�P��r��"؍�K��x�����t�ށ#���a�5jԨ�*��txI|�2��=>p��>�(���'6��F;��WV�c4r<Ģ��"m�<�nz��i������sz�n��� _��k����G���ӎ)��L�
k�t��v�)|����o�������[�D��:�0��*��J���Mgl8�/b� \U!����EQdМtH�p֋�-%�ŉ.K#����V��5V�����SgI4�T�PyzGc�=S��6������5jtCz8G3!*��ԁ�ëHy��W��u�Rs4��:���,<
{gp\��0�+@\\�������!~�V�S9D���>�%_|2w� |E$��ȫ�4D�2���]�����>�I��l㠓H��@4����3�R�b2�D��'���H��S�>��
v|���X�1�#p-�k�lY�ë�]'�R�g��-��9��6"ހr���D�>��oSќ����Ζ�
�L��>B+��8�Fg9�d�,�-O��:��ѭNG��Rq�?M�P^Α�x�;5fܣdO�J�J�Β��r��O��!a���tk�+�Uꆴ��a��F��eN؏�֍bn�� �^%�ݵ��yǼ�[GmԨѫE��l��3�_.��Ksר\&�ǣ}w���K���ړŭ`,�W��|v�}z/�3y�hS���M��,�$e� X�q}w�wp�����zx���X�uؕ���91��6���~1�s���_�9��|-w���8�$ �o2�`��{t���^�}pe��U
� E�\��n�|'4`�ԣ<�ÑSR&�9����
�Ӿ� �|9�MIgS.�� *�#Gq��=������ tp�C���JEo��5j�r�9cS����ƺͲ�h��`��Wut�+`a}����Q �����\��+pa[E:�TQ]�� ����Jr��ة^�O!@y%ڐ�`QO͸�����K�O��:����362r�uY7;�H���?��~�:��+-#^�(���jH��Ss���s������s�z[�s�La�?�)-b��,Ke �d��F�7+s�O�	㳋(j,MTc�r��pN4IN?$�+s@�[��vud������f�G�LqUZXͯ�����2�ѥIa��ug����J?]NmƓ�3A�:�o�B�\��b���9- L+�s �6�(�du=1B���KT*ڢ<g�s��n j�F�nIk@���ԐF��c� �D`VHWS$�6�3�P!��t�&�������#���gw2&O��̿kA���}�&/f~�	�%�ڿ>N-R\<��0ΊL֣���H?AU"��r: ��1��?���}���o`Sg4K�����e�.p�\��K�����pG��L4);A�<�¿ؼ���́.�ހ�)Q�t�Z=Ի�C��ԊjG���Mfi %s4��	SZ?��w�~}՜�#���X��zi��zm��䙈��tO�p<xpb؇��t����rX���"d��sD�ߍ5jt�c��O�����馪��.M���w��ٺQ���'���Zٸ�4sW$�ajK�W=���HgR��\�A}�U�ԽP���C�U8A�<J'KI�8�2
���>����}���������ئ�� 'X<mW��2��1:�Gxϻ߄/z��p|�3�����L�O���ޔ���d�I��(�[�G� �`�?/lav�x�D�V�*���l,ފ��=,3[�D0�+��I(h��~�&� �Ө�͡c�dvNuz$����.�A^�;�;����\��0?w�l�4����f�A�N�1M���z�p�'Sq��f��>6�_~q�fN�'�TM�~��M]�-�+����d�����g;Ա��њJH�=� ���d�����:1��i�k��[Эn2�Flr�yQ��(g��'�Y<�"��֒CVjҨ]�p��P�<�5j�rS�ycO�DA ]y���b�p,���8)���+Z��q+rU��xs�Լ��ِ�y;��1�6<o��9Tn�a��N�@e�*~��+xBv�He����8)����/�O�뤡�Qo�Ձ�f�0yq���y9i�)��~��T&J� ��PH^��>��� ���y�l��a_��Q߱ %/��W�FЖB�{��_H*���J{�A��5��מ��Z���|�*��k��G�[В�o�5�������6؊��p���L�~����k3@ٶt�g���
�����cr�`n������Iv�\��T�B(�K�'mL齔�!�8Cܷ_�����>}�Nc��r�޴wa����8�̥���=� b< ��9]'�cɥN%3`�	��w�/� [H#e��KQ��1}�e5�jHS.����"�qDS�p~w���� 7���%�����6Z��ƴ�����nTȱ��s[�p��5j���%����{ t�Hģ+����cb��f� |���e S�L~V������b?n;�#F�<M�4=�\��iNH��ըQ�FS�lR����$p����%Hd��{z5��z�ɷ�ޭ嵦���ڮ�5��J�;�/���2��&�q�E{���iY2���Hd(}rn7)�i���}������OÇ��@��������g}����'�
p8��B9�ɓ�ΰr�j�.���1j|0�)]7�9E�e0��K ӖO�|�X#K�}���IU�����$���uZ�K|!y�u�WT�
�hV�G�GrN���y��;��#Wb�F�==.����ӥ���f~�s��*��Xj���X�fWN�l��+v O�6�C�w�y���:�du0�EFG���Q������~�k������ݳg'#��r��b�G��n�h���|>������a<u���o��cG����Љ~�ӛ��)�^n�BQ_ ��NU�6.���c�<�9���"�Ĳ��S���
慫�[N��0SHY���8��d�W<��8���!�-��Ca8���.I��g�IU�5��S5jԨN��\��Q̇A�	w�۳��q��]_��<oo�����8��o�.u�p���B���3o��h��5z��cw���v^�A��>�7��$AN���qCv�y�qz�u_"2?�g�R�	w�r?���g��8.v��jP��<'0�r�R�!�<�$���>DxW��/�?�����B8�/x����./<F���_��o�O��?���g с�/��|�������B>�Y8oT�D�j�Y�g��:. e�����&,8;�6�R�sE!�㼑s��{L�i��e�<b�q�է;����k]�ӨQ�F����v��ފ ^n�Duq�	���Z/$H��S�y���6�P6�Y����3\0~:��s
0p����fb���G�^z����߁O��[������c�m2������30�=����_�O����ӻG�uI)�d����:I.�>P��,�62$�,�	�uT�r��+T��11�Iخ�%�X'��&d�
f�(�x����l�j������i-������v��M5�_���]��գ�;�}*�ik�h-�Q�W�ΘN���,O���)9P���{W�/:��e���o�v*#!���J�I���Ͼ�qf�Μ%e�y�·���l�i�F���-�2�]�[?�;�.�Km|���y[���a�<BqG�B;|����ݽbd��lM;p������lJ:�wD�8-�Î�;{�qDٰ.
��N�섏EX�	����܋QEN�8����~�g~>���_��/�����P��	��������O��φ�7����hڑA���TC[	��Ae)��iޢ�$[��Fq�(=2��G�;�rx,�(#`~�ҕ2V�&h����XH�ěթ/n��]��Ǒ_4-O�����b@�o�5r6�O}�4t{����,'��6;�	a���Y�u`��(�F�5�g��]}��fF��:�b���VJ([^t�t�]��bZ���۔�t���fc��mZC�K����ʭmQ�!È����U.H�7*&f�WcU��t<=E���� ������?�/�k#l=8�����.s�<}|�ӟ����ݛo$(${m>j�O��r�%�pS���ԩ0L���?��7q��b
�cY)��j�Lt�Z�I���m#�l��+�+��z/n.�T�/�.k3�rv�Ls�(IU�z�����a%c�\��ݶbͺ8�^Q�P�[Y\�5�F�^yZ{���a]
wY���z�8-�AZ.x#H�S��5�13k�/9v��q�+_����ދ��w��2�0gm����bԕZ����5�si��N#��nԨQ�[�G�5'[HV�Rv��Ҡ���#2�u�	c`�.��~���i%u��c>�<ۓ nE8WXǌ���_Sʛ�xW�5``��dLJ�X�:1���w{%C9�#=�w ��*X
��Ut�E��A��;�v���~���Nm�8|��>�i������������w?;�Ȁ�B 2���p�����?��>8�R�	̔H�bVe>��Q(��7�^����\�4Z+����<̅�5�:�0|d>,���	�1��;0afH64���`J{�5�K�8qM�7���v!�(�q����U���>��uy�`��Q<��Di<KSj� W�3�9��3���{q@lԨQ�{���F�D�<�b��E�U�C�B�CG����2�]IQ���7p��q-oξٚ����Y';V$d�¥��>Յ�T�;=�VO�����)�ر�U49@@U^��ӟ��扇���������|��/�����������Ԟ����x����?��s�o���_���C|6���)���I�^ebc���R�	v~.�y�G�]EiJ"߱����Ʃ0���1�=ߠwz&��*�����8F�O#o ��B��ԝrB��q����&\�� �W�'�N���EUv�a��۟R�~������8;)1ls�(�S�_�KҕcQm�Q�F��\����Q�f����(���}��u�4t�C�����O7?�P�A��޺�U����SY_>rh�*R��L��$�sV�ƺ㕜դ�܇��O��t�M͑�Q�F� 'S��;���8�I~��6a8���\�݆Dv)盥�ݖ$и5�>���A�I�d<A�L��"�R�$?Ҩh��l���x�U	���@	w�����x�����_����{�ܟ����= Ǔ��bP�P�;}>��/����O���ȏ��TڧמF=��ʻ�)E�����)�N���N4�q�"�`�e
�$a��~�XS�����B�'~/Ƞ�1�(���du�K똷<I�f VG<D���E{���h?�K�+�5jtO��8��Om%(]��i�u"�9yx9��e���F�ĎZ;��S<�� �\<�U�K��U[��̳�SR�a��㲻we�yx��d�8�~�E��Ϗ�����������7���O�NLv��1�*�ӿ�'���]�+���o�ү���g��qC�h�8�F*8�(J���g��[P9P��O����jV���B�l˳f�����ޡQ2��,�?���6y̖�]�f����4;G���/稸���Ø˶�rzC�OEJ�r��1��XՌ�J�C帋ڗ훍5j����I���P9B�R2~~��B<�S�u��u��ܵ�Mxd�@vw�=�2>D���f��?���jNr���۱o�5�&y��@��-c��&]:V�2?;,.�̶օWή�4�S��2$7Y� ��&�I.2��u��t��:���N��W)P�� <�Q�C�w���������,��o��[�(��|=���'xm8q��|�����o����~���3�A0o�6*�� 1t�݇�2��( �����f9<����8DQ��"��2�*�L·%�9�&���y����B���'��5YZ���^~�hx�?s%ݝ�D��q�Z����j#6jԨѣ�O�*��6�sm�}d0���"X{��zv�q�tR��-���
<W6�V���EZ��#B������Ѝ�/^��矃�������2��o�6��W}9�	�ў{�ᓟ��c��������W��p|ﻡ{F�p�w�@2,X����o*|��Rp{z1^�"���Of�66��B���J�2��?�	y�K�g�E2g�D�Q�<��>��J�躈̝R�Q������K�KY.ɋҸ��Z�^���+��5j4Ez�~�C8�Nm擻������&��Vw �.A���|а�_����`���H��JI��K���縻�Z;#5j��v���vP���wI��2/�]��T�|\����>,s=��6�D3x-�_�1������H�F1�^.ה2��Euȟt+� �jHG�
ȳ������w�����_��C��?�w�[�ȇ����ۿ�����4�������������4:����\H%��ӣ� �&�s��0���&r��&�T�U�i{]kU7�}\�!B���	&���*tǹ)i�|F���x������FSoo�n�M��Ӹ�󆢏F����{N5j����~��On����D��s��/сp'��&�[�]��nثN�W|Y	]�QI�ڈ�p���!�r�ݍ�����=9�r�U�%6��`��y��c �$a���Y<�~���ݯ���?�5���J����0�L����}���	��O~
�~v��]����aL'$�히�ە�j 闀��_)��/	A�[���b�_�����:%_�n��F�B�#U���f.�[Y�N��p�Z��d	OU-�}���l�<���Y�)~����ɴm����?�i��m��?i���RkW�5����4��� T;qv_{'��U9#��j
F=͋�a�ٍ=&�-ߖ<E�8�!w^��M+�~S|�gͣz���䁣���m�|��tg���;�;�~Mg�7��8.�hڨQ�W�����y��s�MN�/��b�8�#�c̹1��M����g/������d.�W����q՛��r�m��(�W�\]�Ob�gx�s��a�{pj=d�����!��NN@�#��!����N��w��/z~歷���/B�s�O��^��;�ӳ�G�����_./n�|�f,ߙ)
�N-|t��,��R� H��΍��H�+�Vs�� kE�`�`���l�cYj�m�� ̅`��ݦh N������	���{]2��=vl�zk+Y'h�=���V�.�
.��<�P~�rO �;�gB�,����a�N��'����3v�\�ظS�D�=5j��t��z�xj'�u��g!�H�z�N@�n�-4n�B]8���!W���(�K�8s�i��� B��B�R+��!�&�f��K�3/m]��~��Y���Z��S6;2nX������ށ�pz���0�5�S�>���ħ���7�ٳ���d��:<;�8d�~8}}+:��'�z);�<���ho�6������.��SF�� �Ņ�E���:�5xY�Iu�P6 2,�Y5T��d��ִ�Q(='IO�u������^"A���,E/���k9�a��]������t&�^��v�c/a���h��'�a��F�5ZD���pc؅�ʖujo-z.�ܺ�8�[;���f����0�y��u�jsǞ���/
]�$�sQ�6����∬��lC�8+�
W�T��Ȋ���L�9e��<|��;�&Pm j�F���5c��q�fxy&`z�q�#���A�HbD�	�p�	�0E��]`��u
g��g�X���EO����!�0�x�N*�����5`��� �%�>��a�����r(%��Bt)�����t���ز���c�:/"��奜7�5u�~���OAI'��ǔ9��)y��FxU�u@~H�5$3~L�DM�+�Krf#nЙea֦�q`w�Ƞ)������1��XqmO��S��W>��!)/�a�l�b?�=l������\i}ш�g7:���>���g�]�F�=2yq.�N?��L���	8gG�Ob��c���]ү:��Ja��+/h��Z����֧za{эQ��s�¨B�[ ;qr2 B%fB��y���
�=�Êñ�Z.�N��~܌#>Ⱦ���I�p�cjDO'kf�pC���ɸ9�B>{��g�h�C�P�����.7�t
�Ș(r֟��#-Q*g,[iWU���5��P�6N��rקBF�DX���^�fR����Y{G��{EǱ2��d�ͻLqz��i��˲���kU�i���ҷ�̆dN9�֦��aJ���*���o��[F̙�k��(��'נ5j�h!-���,�Xc��g���8���x7��'iBƑ��y�4�����/3�79p�ck^��J!U�VẄ�����
Z���_	7W�Kk�"O��q�htY���]��D������0�!����ȁ�P�5���"��7�2ځxG��X ��������S�g�.�{�7n��u���)���l�z�!��A}�BXO��*��.GC��q��T�~�/�hc^�rIy��{r:�y[{c,x�¢���	eɎ6����uH�/���4��O\�^������['�cT2��.���8�VK�ܷ��knq����h^��Z�(<Q� ����9�S���wJ�.�v},�^����Q��w�6�=�eߞ��l[����e'��}Wn�z%h��.�^k��� ��������l0�ꤞ�x���T�J�Ĝ�� #t�t#��[)�����p��`C��脥���m��WE��w�Kڱ'��+���5���'hp�h��f �'�L��w�JVm4@l]K�	7�h��� �Q9�u+�p�
am�Wi�}0�'o�s�&B��&�5�.P�˱5j�h������ƾkЮ��dS6#��� �=�R�8
����d nI[�/
��ث=[���ѸW�z�]p�l��~�;Q�;R}ϴ�n�e�7M��	���ey���ƌ��;/=��Y�_�#Q�Ƽc-h�l0�#̐WF7�q��^��0a��(SK�� �����"�N���c�1��@�W�WG�w
�e3�4#�,��i��.h�Ѳo�α�I��$�>�w�ۄ�0	�f�~��:_��9�"g�IeC�,����Y�Si�!K�5�={nR㬐�6�_�`����t�tS�L�>�cCQE�myHos��?9|�Fq�m���^=?�}ѨQ��S��}�q�dP�C/�fk,'_���B�������3r��W�$I��3�.�a���=���O�����k��7'ڂ�:�਑��k��BV������N�:�R`v��R�b5/��^2V֤x�5�$4��BrVQ���+���j�J:��.�ǉ����A�0݊��l��Y��_T��嶔n����z�م�������Hz^�1��~����V�FM!jԨQ&o�����,gl���I���8f&�I���"�Cu���#�}#m�B���3$�O����kTX��.�`i�}l�|���qN����7��fO�X8�X>a�X��F�#Yg�R_����7֌9Kg�k�#�<�u(?>V�E��$
����0?��P�Y���=���+���
[�Z
k°z�Y h��%C����s3���]�/zWG��pQul��}G�6W݁۵�"��J�[�t��~���()��%2��4,�b���.�!��M�%Ј/���>�`2E2����g���ih�<?x�2���;[V�T���m��H�Ӈ/i�Y}�:\R�-O�`qdt<��&��<憋<Aԧ �|�GL��ǲ�W�!e�����~7�{?R��}�u�Fףk�k�ڳݯ��7]z,��jqAI$O��+Bqأ���r>�j�����hkg�)>m:�$�y�dqs;��.j	�?�c�]��G��T"�-ʼa[�ۓ�k�7�����7��(��⿠6��S�����)�B�ـ�Z��\���v\��c$�Rb�V��c�9NeP�~��U���쥉(�?�
q8[�Z�	,���9$��k����?Π(���$�o,܍T����O+�ӊ��a
J�)�G�Q5jt	�cMȃP�ut�/Z����추�\��c��]�p)��H�[�2O�qy,���[Ҷ+TƂ0��}�
�UX[���Q�p����بwY/K���:qȰu��r'x�Ns���<N�p_��޺������e���)�������O����-��μO������@�@�tq1�[���"��N��0�N�;nȪ��#(+��aȅl�a���4�a��ʚ��W�%�A��Ϣb�>p�#�9�eBe�,R<���IR��
2�
��� ��:�yW���ԙv
�xʻ�eL����o%���7*�$��(=r����o��}Of�f��C~>ʭt���XɅ�r��}V���r�A�.��OP3Z&�{t�{�3'���N�����ݳ�S��1��L�(tl��:��}�q��'p��y%�<��0�J,�~,:ꍅ��8��۴�9�Ê����y7�yßW�o�[��e�F�h��	ݮ��=���z��}{NZ4e:iM�{���j���x�'�c3Lѥ6�L�P򽦴��qN��+�}�UP��&�����;`S���� n��%D6���,���j���#
=�J?e�]�O~6�.�?��4�R Ra�%��qX8i�\ݗ�'��m�36�Qӵ�u|ҧ�[,��Dm��ޅ�8?�^}�m�M^��Ŷ�,�Z%�4�3�ךc��I�;J8~n���.>yx=겵]=|�6>��� ���@cyD�-
����+��r�v�fjr����g�֒%�0�+�j`�4�z�=��u���	;Y�W8�D{#c��5j4��ۈ:9��+����s�#ֳ�&)��xW�|��Tbb���0�N?^���xR� �I����2vZ��y��Q���A3���i�	B�L�n��8�sהf#�%�����T�{d�;��	0�T���%3%����MTg��=�Ng�wp獭6�N��&Ұh\�E[Z�\I��h���*�-��d�7�g	�c
��Q��P� ���6�L�R#����d1��¢R+ �@KXG"�K]f��i
��HEo�!�D�b��M�#���M:��<�'�H�$�TF��6g&ԕ�<�KM�n	dr)E ���ZBr���q� ؔ�Vǒ������.�����K�K���*�W"o5�O�,�vfl��	��1�F�{j^�{A�U!O�����G�a]�&��ݛ�F[�f�̵�-�69���0o3�{�7s��p!���S�"�)�#�%��[�Z��e�(���d�6Odm&���<�J�4XR��w���)R,��b碈�6�In�߫/�S��M��Q�>��V��)/�V)L=��+����9�+�<�,*4��nl�/�����d;��:$�$�
�r�6��b��(7��/T]�MzճW�^�ۣCݫ@N�v��	ǻ9�����odJs��EqV��,2a&T`5%�2��5zt��?�3��mQ�=��F*��ż���kq�d�#����yY'yܩ�k����8����=s7��*��D���7�:�6~�FeO�Xґ�%�7�UӔ���nؙ@{dq�<�uvϕ&Ļg���]Us��gXY�K`$3�Hp�[d]Fe�I��ۡ�;�PA�;�zF�N��u}~�༁p^��lC�D���y%�K8O�Ө��) x+�V<)B�ЎJD�B�;��Q����6 �P_�	]lY0�ST'��=jI���E�@�-�$'�^�,#�eޤ�,��9�8X�X+�Ӯ;ೢ�곭�ڂ�*�fn�V��9��N�PJ�4b�\���C��9Gu5=7�i,�/j@/idSaVt�)qR�mtU�fSؔVͦY�lmz�,b�� )9_"��bf�X2�-Ck�9����Ѣev�Щ����qH:��變�JAC}-H�PC��VQ������`�@���H�[~�~^��I�E^��r�-��N��� O���W:��_U�>ȡ,�V tt�qT!�t^��P��*��٠��(��>�]��
��t�5`S �E*[��\�]�qW�1\���k��-����ǉF��ǉ���w��zi�O�;6S;���W�E9I{c4jԨ�Hx�����V�ťl=*cefl��U��;A�y�����A�h�2���� ���h�X�+��dC�ղ���4ow�5Iv<	�{�O5j�h-u��N2Z�G�e8�1����i���ڭ$��/���$82,�\D�>���m&�@1'	ڔL�������h�q���b%uG&8ajG��o�!f@�����%gP˩� .�5S�W�D's�t��(��#��v7\��w �ߌ9�J�(�A� X�A;�H#�L����7�*��5VYX�d� �U�;��-�εI=�O)H/%|5I�H?�j�"�!��7(�����_�&l�Y�רQ�W���P��6�e�Xb�xc��������@����t��o!w1�H�^��Y����R��Ҧ�B�6O�?�6Ȧ�}!��)�K�ճw0=�C�O�r>�o`�by�����Rd��AXք�p=�#28�I Y�2H����ߥl]i�� ��D&���c/l+�Ρ�	Nv�c�`_/]f!9fRiڶs�!�b�������;�aO\�f�㉷�w�e��W���q#L�?�~�Q�F/)�t��?����;�J�f=z��u^�ߥnYV��$��/��W�h-*�|Z�Xj��K����P���A6�Xf��;�NsC	���S����?�J�TX�n�6��-��Ү�'V��w��;m�5�O�'l}dWmw����FBOyu"T�90#S^���� ���"R�`N��N<N2�؝8<O CL<�i,�8�{|Ej�y��w�������f`+���H|�
T<�;�PW �4�"�*�<j�Y��¢��3�OrА�$�����Œ�"P��"\@3غ����T��Bdl6a��^b��%��
 �6!�^�HL�ߢ���1���Q���;�끀��b���[��չ�VM��_�Dۨ�5:�T[�$yN��zP	�E�9�^�fKm�\B�縫kbJ�;�C�۠Ηu��| ��>�zP�`��l�F�	�� ���c��+֞� me��Tǎ��uB������>��a�<@�wF'a]k0I��Z�.m�	���@��
g淶0�	Y�m2�l3�:+�&��o!MTEϦ��xe��<:���X�ꦣ/HG��Jdr��.�ۄs+��u�d�/ضQ\��OLQI�l��K�EQ��+��(�:і�ud��=a��Y��IF��5�=��iCz�2E���,�k�s�To����x�h .�%w�)��a~�ܖ��iݭ��ªdT�޳>�H�.( �SrAu#�f#����!�0��\'�5j��"�<-��캍}^?���O�@N|���K��0f�q�<F�=
���� �(�[�4'�;��Ӡ�rZˠ�Ӵځ��XG���J��f}��4�(lY1Yg埾�4��Eh�5��T���E��>��be)Ң?94jԨ�<y�Z͉�#oAlIz^��̌�y-Vm��2����?���	��t���T]-2�yl"E L�94��^7�t
V-�r�:�ܴ(��s/�w�e.̾װ*��:>>x\�b�|���<�̍�MgM�����5^ax��c���_�5�*��K&F.�R�*{��EE_2s:�9�U2�;�<��L���Q��yV������C��t��UKPu��	���,��g�}�
ljf��b�k`!��Ggu�.�XG�)]y�4K'��\�s�=o�!��v����$og����^\ �Hy{���S�Yz�sj�F�.K�5�J��>>�[ �y	pr��1�K�Δ�Mo�l�<��Ru��B���O�n6PN�D�>/�aN�h�0`Ԣ�Hm\��+���J�c�A��Ž.ᒢ���6�m�~����%/�M�Mɞ!͟��QŦ��Q�H�� RySJ*7Kg�8N�<�K��H��d��-�mM>e��?F��f����X�Y��L�<F~1&b}��vtFr�Y�{�6�Ġz�2�5'�ykۯ�9���w��W�SX��z�����3���Y��I��׶CCX��H��i����W˓���C��Wisʩ��n_�5ZCY�	G]�K���TWb~r]�nJ�$�\��eE�89;��.n���DSB7o^m:����J ���4���)~:2��+��ϣ�H�3^����H<�'��M�_�U|_�Q�F@5��y)�mR��U~Z���<o!А�� g��(C#v�=,���m����)y�G��6Z��/�~����U93)1d��+u��e�ֵ}-\ۿB^�D�*R����"��}��K�B�c����"�]%c?2g�z��m#d�d���������� `e����#/�S��w(��P4T���=�+�Bm 4)A�s,fZ@J�!�c�uY���鹽ȅ��$.��1��^
H�Ҹ�P-4��;ٮi��ݛ�;u����* /X�_5jt�M������ǉ"}�F2oh��\�d�.��;&9�l!y�g�%�(becՓ&}cSW�#����	Q��`�ෙ-��iC�;��t�:,��ه��l]��	��]ggה���$�C���Y=/2~��/��$���#�"J�G؜d�`{�Q�ތ��$z��6���"�w�-(˄Z^�QYۦ}�<�p�*�-&N����3�V��{��[u�k9��+!��7�&�9��5P�n�Xm���mq�pY�M�mLa^�GY��P�EM,�ɺQ�F��[��Z�B?�m<=m�H
��x��,�7�� �d&қ0?��N�PWI��ɁC'�t��~�y�M=�[��)�{�7���e���N0�s�e׊��nw�_�o�3)ם5vc�-�C�F��4u�a���#`�hY�5c��Xj�؝�N���<��q�9)���Ɛ��{�ln�d\�{6���H V�x�CC<�26;�,���,ֶ�:[��9�����'6{ )N��)���Ѷ$#�e[�ɎCHA� �G~��'��	��	�����%��"+b��,Jg��n�I���û��]+�j�U����>���s�jX�jM�j���3ŎE}�l���0[��5�J�����Q�C�- �@s�IPj�̑�����Y3[��@��ٱ�Si Ev*��4풋�-C��T�q& ��7��S��2Ss���o�w�.f����,=6"�8/ G�8�Z��Z�l �<_:(��-�C,���zE�*ZsO
��sj�8�g����)��r�x� �,S]�����_��q�8�-���}�3������\{�s�����g�8��f�9��3��voji�˹ y�i_}V��&����I�8���{��і���ņ�]	( h葵Z �gͫuBt���J�	�������JKA��=!��7Ef�`�ڒ1D��!h�R&�n����]���a�)�#��ȍ+��蘆�3��5��z&noɄA�"OB��`��_�u@�;l٠���vT{Il*�h���)"��:��c&���e��ќ���-��6O���<�z�u��ChZ��ٝ��q���W����/M�|��~�V��-�pq��~�mY[	*�rW���nG�p�ߖu0�i�P�  ��IDAT�t$ĉ��N��_b+��ȦC�"#����]�H���R�'�#��"��[.F��}ߵ���L�f��� �)�a�l���Z`;�n�������&�:.RDh�֑[#9w��)6�j,L9/�lp�h�iv�ٝ[^j:�. 8qSu���ušqe �ԭʶ�E��G�r��-D�؀�E��R���uo�~��g0H��y�9�|�ہNC���REߍ��4�b��g�����zֵZ���Q~Vi;��rf��0O��;�@�!��3��l�h	r��N�d� ?�u�<�#s��8�U�3rDz.��^�<���+�)݊�U���+V����T���[��ѡH�plj��ӳ(���� Y�DM�}<L��@��Uwue���?"C�lИO�1�(���6v�l�L�4y�@�;�E�����L�� ���ʹ@�:��� ��,׮�|��Y�$�+����u|��N��O`'�v9"�H՛D�����,C��+�?=^��w�Ze�0 8���X#�a�n��h����
�҂d�K�Q��F��#��<o�����l7p�rGA�ɺ��?�,�g�X5�)�S��Fñ�&1r&���@���
����Ӊ��J|2[rt��C���Bm��`9]:k�+K�NU��r��~r�S�g��e`z����� �S�{�?���Ŏ�5Ol�"0��s,>[��]; Am�������L�� �����Y�Ai�)������H'� �L+�c�ל�+!XƓ|yɼ?����Ϊ]��֛Kh��|���n������8��E��i�gk[֗b��	,����X����q��C}�A=�bW�I7���&|Yi�K���d�:_��?B�ܝ�D�aÎ���ݴ�M���Џ�j���Ch�D�����;ڽ���ϭ��}�3����͕p_*5�n��s�a��v� w3l�e��D5��;�߹�V��]��|ҷa���ڔ~����=_K�����RY>�sa>�Ϝ��&@�O0J�\�X~X��Mx�VP�bUn!p@�Wuv�k�Fm�U�U�,7�B�ir^���EF<��`���7��Aޭ'�_yo�A���4�]�D�����f1�cR���:I�:�b���{���n�zݕ�Q�ŜV�˙8�L��� (h��
�Z�G��:3�����?e�H��J���к4�ξ��y��#�6�*�����0E�w��җ���(2�O�Ḇ�@v��h@�:#��H�;ů����R~7m95�=���FY�q('�w�������A"��x�dqɷTP�x�N�M��뜂:	_�Fc�7E0L�J�'n���f��3��4��(������#zV~�mJ/DG<֯���dZ��6����\+q�Mf���]�2��N�"c��N8�ޔ�S&�J�w�&��g�g�h�YW��E���TaV���&!�5:�F���X'ܑA�,	8��I/d��������Pg)HOe�����&}��;���8�Pf=�rY��r���B�8����hڼ�;}~��C�p��6��y;����N�K�y��߯o�r�� __���PU�(t�׀�D��Ƞ6<�Y3���#�������n����L�,"]�yҷ���sD�3k�iHt�H���c�#���#���~�b��!�?H�L����ґ�9�~�y����#l4���6QG�d�融������VwM�����ڿ��[�U�.��77x�5�.b��f��NJMAZy�k�1D٤�w:��m>�I�o��#B�����m�˦`�Y{
���9�oF�.B�Y��>�-�݆���>���f]���Pos���|����#g~�m3n��Ԙ�y6�q�+�&�(H��[�yS�Σ���M������`j-�^��p� �\����l���;qE����즂����VԦ�����lu��]�t���9A��ٹE�Z9��˽�ݩ�λU����EWqpɕډ���ղU���K��qq��R�ε�:	� �:s��7���c��>�t�jb(�q
�9̦8�)���^�^B;�>^�w������k�Fx�c�/|�{�����0���k��~��_��-X_��w���3Ev~PS��� ��TYӬ�~�
9�yHs�K��1�n��}���`�����g��ulCip ���:��q�nǸ��������/r/�=U���UY{�]D�PA���L�Te�DYQT�:by��
p$cE6���Q�ҫ��5��]�E[ܮ@���h|k?�a���0m*�Eإ˯�s8�D�b�<���z�nxǸ<����g<�qW�]{� 8�9���������~V�-���oz�e<��`/���w^_�>��+���q�Q����˯���$Ӄ�����M�����j�6_(�/���z���Um!�� ;��3) ���"�������㉷�����g�U��/~>���p���9p��b�(��"i��;B�M�Eϐm��ߣ�-��\Ʋ�M�jX&;d S&�>q��q��ˉ���X@�~�,8��͞���dI����.�<��Ѿ���O� ��d�D� w�{��<v�9�a�{�F�P 4�%�)2���@69�)3���d6�*�@�������ɂ6�г�����V��cM�)�c�1��LiOe��`Kɳs��u�~��z����Ї�n�}��u���W��E���zuK&n
�0�PK[�2����^ s��x���u�g�m�¹ʮ�o���8J����*E�PT�@o��Il���!�m����H�ƃEK������uJ�=j�߫�>���6����ܵ�]�l}��<Wn��(�A�$�}���[��5��dR���^�����������q/@���3N�a�zK��;��K���сfZb�t,Pr6��������_��
����%䭘]���~~�3����𻯼
kX�܋��;��w�a��ԅ6�S��p���\�����ѫW���%<vt�rn\�W���b�8�K���g��7]��z����HC� ���S���[�����NW'�����_�	_�֋���í��M�0�3�$e��A���85;q.7�Z�N�$/?ݸ�V���n��wZ�G�'=ww�l��'�f��.�D�FK��Pm�����j�."%�.�$MsZƭ�S+�;�]>��~��.Z��M�����[Î{�J8��p��*G�/`��V���l;G#.ċ	�5ԛ�ΥǈxreN�[��M��EǴ��z;�w5gB�k ���:ME�3�ud`F�h�@�Z;%����;�G�6=�@�����|�'�W~���C�<}7�5�f���������o�&��O�sxv���I��)Т�]����b����u+�s�$H�g���9K��k�F��ʢm�+���<zt�2�;\��ˣH�m�\�<)�hw�{������6CO�@�\���f�Hm�sk�w^��<��K��o�/��̶�#�<}����"�l ��vU�*��I!��~UZ�f��6[Lz/���̶Vs<uS���%H�^�u����޵�[��Kh;�g}ѓ1.���D�ٶg]���v�;�P���a������}�7l�3q�^��~����`���+�@���lۂv�E�l��7��^�6�UO�u;�i᣾7���$��2pL~orT�0��G�e�D�ʘFb��E_�[�vP�Z�
T.n�eT�<��t�,��~�9ٹ�Q��7[}��;���m.P�2:*A>mE�������Ӻ{��2�o�m�k,�h�g�Bv��޿ ���!N���>Mf�9_8C�Mg�AF�[��h!�99w�?��������iyv���#��d�����S�?��`�^�A���8 ���}�����������7^\td0�w`J=�,�-��S����8�� �4��� �/~/��_�<��p�h���z|p��Y����#���Hjs\B�?t@t$O*ŋ�5����������H��yr
��_����~��g!>t�¢�;I?�	�ѓ^��.�5-�����RK�r��y�Fԓ�w�[5��-���eҬ}a�Bm�l+�~��vgna_lt�oƑ�U�|�>�Q�Ї�{�cVf��i��ҙ��:G����F�2uM7�=��r��� �.�)8���7���[~�	�{[�`���^���ɗ�$7���Yo��;T����_r��.���XO���R�tE�l�w�ް�t>�q�U����K���J��S8��O��!�����=?<����c�ă������w��i����_���Uκ�t�Pp�j�
�f�'�>���ѯy��hS�W\��������_�Q��3�= ǣ��d��C�Ƕ�}%JJ�y����t,+��lˈ��ӳ͔��`�6�����6���M��~����� Ͽ�:ݸ���Kǆ�r����Z�����Տ>N�i_� b���k��/_};���i������a��v@���>�p(/���VN�e��k@�Y�8�����wC�w�Ս���v��^��-�nc�pC8��˭�bh�I�}֟�������%����:;��/��6�?�\�q�*��ҕ�o%Od�)�f�"���.�NB�ַ���2pLj�V�>\���.�}�([Rjl�EMK(�51+�9%����f����ϕ����rQ7�1Nh�.������V����X;9'u�L���,�}������{E~6��{��8��
a���#5�ޔ�c�N�M�N�gǇ
}y�O���УW�����Y�;�m�}��� HJN�'\F�e�h9%����Kq|�K�Dc?�;-�f�vfm��8���`��u#缸x�A+���8(��H~��@|[2�|��%��/���Y���u�pS+��W���z�����F����-OO����N�����p��r�j]\sh.�����0��G>_|������;�]3c ��x�{��W��D	蔚[���˯�?�;~�����qH�+uV�:L��{�V�(Um~z`�;֌k��.�P�S�+��� ��G�O���ާ�����������z�L�)�	v��p���E Vcx���nlef��(,ެ�P�t��S��� ύ}�i�eo!��H'�~l���p������Q��,B�d/;��V�7"d.����G����CZ����Yp��M�Q�g��L��|&8�;Ҭٟ�=S�~?>sA��1��Qg�s�pA��p�ܯ0��ts�𑋫��-�s�̧;���N!���Sx�V���/����\���$'z�R�:Vw�v+����ٟ.ځ�g)��(��ee�d1�ր����{�;P*���V���+�n�����6,j��QH�:�ȓ��?��M���g��'�u���s$70t�]�Ï~�����~��/�-@)�Bu)�?lKבZY�E����l���K��+𡷾�ÿ���3O?�izbMv�1�a�_�Ud{Ŵ�>�Km�G���>3��	;|e��8��������߀�6��?��ڭ��,�)P�>4����nǕx*
�_�ڶk���"����D�V��9P�ѵ_K��Wo�.�>*���ʳ�eܯ��2V����x!,ف����WOoF�tE���0�&�;�zC�9�a+����o��p��fg}�'������2ٲcl��7G�W�U9R��u����~���o1�t!e+#�x7�Y2�m�nB�!�/�`G��BKo� g��,.Y�vM�6�|����T���xe�?����D�ٽ)�F�=�ɼu�Ŏ�x��,^����|��p����ڇ�YT&�k�0���e`�{
�ٵP��B^���m�Ҥ-�+�|��g�ã��6� ޡ|��p����)�c��FS:�^]��SY��B��d������:�눃>��Q!�tv�C>�������$<r�:��*�9;��/�
��u�~���~���a�R���؂S]��F��׀���ր1�������	���8�@.�0r�R�)*h�C:L��4�ȹ�Җ ���BD��`���ix�	����/�s���� aA��Ʒ<u��m�K'����E9g��R���٧�vSz�RҶ�8�y~�7Q��@x�3{��\�E�;�W֋������=_�ee0L�����W&�OyVyE�����i8��)G����z�T n��p�l��<����#�<��� 5'��e/y=�t<ԠT����뒡���vu�6�م���X�%�d ��y[���""E믏C!5��,�5���/	g��׹�@�:m��:{(o���������)��/��_���{��Zq��>�����>��w�~��`8�sh��m{��7� =�<����0�m�N����W������|����
�Gr��c�OЂ�O�숝*�:v���;j�.�1��t�_����O�j8����_���᱋�f���~��+�b$����։���|.����X����"��ӗ�DG�����4�Ϛu��;�#�{�1��Z�x|ʦ�@��e{>X�i�D�eD���3�aY�L�v�]����ZA2u��!�OS��y�rks�.�gӦ�� �!���7�$�5��#rY֯7/R�2��i�k9� m�ob~>gl���OִĮ����Y(��/�&�����Mg�����݋�¢t|۱��OY1e@���IE���s����� PgZe�p��ꝷ5�g��7f���b�3�D8k�'��$��9�Ž�`�{�n�U�ߟg��ue�o1Ԋ�`;E�S�Q�\U N��ۮG�mR��#J+�u��!�|�{ 摒y�}�U5�#���}���@X�)�xb�S��su�C��c�#W��~��Eϸ�]��ZmE���P��DCngjW�G����ix0mñM+�')N���#�G�cPj���K�ҁe�
�(�]w 9
(˚fy�]�>����%������9Us�(�Q��߈�94}z?��pT�2�a/�x��ԡ���9u��⹩��j� �Cۭ�� M�ٮ/w䔶C�.��7XP��s)�#Nw�����
w*�� 8��U�f,�p��3?鞧2��s� ��I����y��D p{q�n�A�R�P���:�E^;}�g�����g�,f:U�k)u��T���/����
����I�e�@>�I�N�7�Ín����+�𕫔�B6�u�������N�w?�68�?�A
Qr�Y��	u�Qvk��9�M��S�0篁�F��?���|דcyk�4(ǥt�$�	g���{<Xf����+$�y�����Q�.V�g�%���}Ս��ï�s�k��2��ň�>g%��st��hR�pvG��i���R�Ȳ!@����]��w�#\GW.����7��߻<8n�X��b13�g�#^�vY��f����`��S;���w9`C�on�:�jY�ty�`3���<ū^��{|^�fo�.7	���V7q��`m+�i|3u��s���wo=op��8�P�%��l)�l��!�j�����&E��fe���(gʂ3���� �O��Y`b@M��bUF��A�8�P8��!� ��s%����)9���V����X��E:�P����߸��4p"�^gXc���Y)OD����^O?�{:Q��NNCM#����3�Lq��,��I�;�q���i�_ �y|~�~���s�+P10;��%\=>&n::h����M#��;8�F
�HU�؍��p�����E���7ANo��I�ue�e�Tǜ׵���;pyn�:WN��#��ǜ��#o{�y�Q�ԋ/Mّ{�.���х=���VI�c�2�#��W<^�	��e*}�ͪ �_��-�0X��%�����^��#�N�<�n:�&���i5l!��Oܻ�Hl�ۖ-cێ��If� ���|�j�bNq���u����~�5C��#�S10���Qڼ�3\U`p��2��A5C���Y����j��z�oظ>��+U���j,��k�����:=����g�}o}Bʼ]E^Q�/y���49�Dp�\�����+[TN�S�ykx�;�}����q�ǹP]�K��x!9���#$�0b6oa�ԘT���k9pC���u������w?�Ux{Bg	ɾi9JEZJ^��X��ڶ-��ƽ)�{�.��7�gn���Z���SXcwz�>��9CP��3�N/Ѩ,����#��mNe,����o�µ@4#�
�����|FA��B�p�7��
hz�ƶ�>+��C��ᘎ{Һ��t[+�|�.[ݝA��=\�^����q��9ܒ��u�~���I�ci����"�}`E��\Y����4� B96�G;A��	zS�������@�p�Ɖ��_�� �PP3yg���;�|�E��>1T�wk��I���"N�ڸ�mf_]Y��l��m+}V�m �����p�s�дR�łSqT��mek��;E��B�9炪�����X�::��t,�*��i�7X�����|��'(��&����w��I�!��+xyuJ�,:U�Tn1u06n:O!;Z���ࡣ�!n�RB�����M,<"-T� I��>5Ü���S��5?o�HPm�QOgE?r��|6�}�%X�#_���lh�Pɷ��t�K~��fX}�%wr��έ�0Ee�t9����������@�7��9�����._ �v�Y�9L�L�Wȴ�|� �/�뭀������6]�]��Q;2���CP�p�;��A%�j�ԋ�T������)�N���[�^��?`:�J��E��>�R���؂^?+��Rƫ�	�yP,��֢�Q�|��M=�����7��N9-|���	��	��pV�׿�ðLe%C#��!�R��o	����IL�Mg=�nU���&�b�a�s�� �ᔲo�{!��*Z��o��}?v�,����C1��G8=?]� _�~6	G�~�3�G�^�WV'd��rb��ǹ
�����V�6�)�V���Ů��0�����ֿ݃�>錰���׿��U�jJcw��7�A)�$C�k�5 �3_Sc+=/Y(AX�����0{#o��j즼B�x.�J��lF��Lmϴ6?A*[`S6�}i����RF�̋(� �/L7i��N�73]/*3�Nx�x(E,�h��&��d[�)[��W�}VPb4�?���T�(𑏁)���OX�2�����G��B&�������]}F�@
�����AG  *l��(T���O�/fg+��LJ���D()�珝)0��L�����U����c@�j>��V'p�\�2a���mj!^fØ.�j����S;�E��ϋN�C��7�I�f;5-ՙ�>��0o�]�i��Nh-K�������~�$BN	��-�΢$;�*_6�93 ���U�l:���pFh4J�U���՜��A�����,�5�Ȋ�:�y;s��1W�Zn�(� �.Tu��/B?����w��y�=z��c��Ɂ��Wn·o�}ʎ�ܠ�_��se�窽K����ַހ��
����X�.c�E��������o?�`�P�!�Gq��cх�Јd�f��x}�/�O?�?��8����~�	�����U�w6���K��n[����s�Q��ӷw�!O淬0Gv���j� �̧ۦ�pΟt�����v���0�DAwE����M��	3�wڝ��Ʌ�3�� �>�'ح�p�<��<��@�	�=�?\b�qOﺛC��q��E�X��2�7t�K�p���U/j��y�OyY���ㅱ�M�岢B�qI=)�7�7r¨��G�k�:�<�(O��~��k�MX�@E�Bj����Nq����#JM�xUj_�ZF���]�G�
t��pe4�l
ux�R�"Eg�&z1$����������D���uo��[/ւ��(H���������o
pI�)*�K߻�i����ֈ�a��(أ������F@�#��\����W �P�'�/"M�!��FI�V��!<�ezF7��H�v����ք�֍�]6��;�u� o����[�/}��~�;`��X�Z��� �+�v�&�P ��M"4;o#�(	�a^3^P�PA�m��J�A�l����Fz�����;�̶Z�)m7��{/�ԉ_f	(�#_�,��K�X��́�C�z�բ�<'K�HЇ�#=g��,�yN ��5j;r�y�{�V�˾p���R�E�s���j��8w?����	^��=���m��4��3��/*�g���Ӄ��t#�a�l����\~G̗=��/��DB���l8R��@�(T���/1	���A��.t�cJ���,jQ5r��(�T�wP�(�h�dF�:+���JD>����y��+�~Ѣ�{w�'mb�	u�gҋ*�"���� �b���^���r�,:l4�AR��hJ�'���2B#�>:�y�9H)�@�Ǖ�$U���P���͊jP�I�!���C�DN{�t$����J�$�l��!�;Ҹ-��r
z�2Xg�g�&d(�?+U��̍��sʭ��U9�[���L� �a`��zo����?�!�j�pJ-d��?ϙڗ�w��O�)�p�&��K��.����6�y�Q�B��}L���� ��d:��u������팑 ���FAǷ�!�mޓ��,�w���:Sr�Y 	�>�k~��C��N5��HAƫf��p4f��]?������5�K�Y�c��D�(�P2��'�E����;�I��	uW���,Z�2	V����í�Ф0���x�d�9HQ�0�n�s��N��vS�KggyoRnU�ؒ޶����,6͝�1p�����+���/��T����N�j]˕�J����GZ���2��J>�~t���bU�ٹ��^d���{��3���h�)g��5P�Ċ�*��nWm;�F��v���uߜ峱C�ɣ�u�飡�'�7���9���������7��(<��[!�b�_H� �tL�ԕ��v�~�_���kX��`��Z������9���@�a�|�U89�ˣģ �M�㋴�Ma���K��-z7/�d�2�4�j��g�F�����2�c��~��Cu��� 2��!�nL��m*��Go(>
ۥA;�[>W̶L�VC�q�|q1 �xy�}s-�=(<яWڵݳ|�G��)ωxh΍v���^�L��ŸrQ�K�@h�"=�6���f�\���]��"o7�E-m��	D:/�ƌ���5�o�ܼ������z�M��P\v��{�ot������k�zU%M��7ꍷ�ìs_�����.���_���eGe�>sbϳ�u%�#�:�#̰9nr��Ai���Մ6��8(��!���E"J+�׆'#GH쌧�S&>�P���J�|�h�0Ң��] �Y�n%@�b�?��z�
����bȈ��K�V4��=a���	�C�v��ԏ��p��xfz�o�Z�v'�7j�l�o���z���Ed�y�7�0��9���Y8-/�FV`�1�8�<��s3^�\��r�{F�D^��%OU����JpN���5n?�4 i�k�W`������Zȏ��C>�|��{�{{t�<p�
���� �|	���7���pHn̾+{��P�ۙ�j{jg�[������ ���CU֋C9���X�f%��ce���?Y��c.9	��#,mn#��aU�xC�U>k��Gn��-������_2��Q��@����*��<tQ�)�寢�3e,�Unlen�${i0���އ��̢��"�6L�G7�q��R����W�b@!gk
��B�oh<�;����v���Ҽe;Jg�ӿ2)g�-вi�� ��P�J�q.n�37X��3�����l�p߼>�R�o�NDĢ�lG�߁���P���r#ǿ���qIN,vzJ;H�Bp|u��/�0]�;L�+s��IC���n��Q�>��u�#\��6�kk��5�+4��m�i�Q��H���@��e����a�+X�G_N`�_��_x���9�Li~�8	Z����`A�t/�N��3����7N��/�<�$�Gg����2A.:�
���6$��.`'rF�^~)�"�&fhE�<k��Axe1@xl�yܷ����9�����	�y��T�Cm��a��Ӎ�+O2jh&�j�hw�ֶ]���R��b��{��`h��`�ll�y�S��2$ِ�Br�?����2^EAR����VCl)�@Xn+�)�!g�P�v����+-`���P��Q;�}���B9�Dg*�D������?���/�g���c~.����yҊ�-����MdL�X)ñᐞ�� �>$V�����bk8>3<�m�B:S�"��7]	�.3-��@ת&=�ctU�}�9[ +��{��r�-+�b�u9gGK������n�(Qܘ�gz���(c!3��х��8!U2�G�Z-IqzI�7}�YgpX�����(�s�I��]wx��g�Y����"�,�����(.�8�y����y�I�$� ���Ȅ.Ew��f�GQ|e�:P]���J'��N�8��澤H��4�*��ʴ�U��u{1�gA������h�xwk��Ι(I�iЙ� �,y�J�� D��._b�Дw�C��pz�:;+�K�<B5<��ݬ^m����Y5�.J
6����~���������̒]_9��wd���<�<|�߀p�e$E,�����O�G�B25���0) d�4���p봃+I7
�(J�*�Nvh�-ʅI�l��|�i��V&�y�"�I�uJ�m��@��T��#8>�8C���!�w9�+��+��_h�v�:���ac���!��49���h��@�I�Aqv{޷r������:�~������á�=�ү�C�uu98�e[kO��y~Ъ�I�F��T����.��硳�݈��UD=���x��Y,b�|G��^w,���(�F�%v'l���S٥;dŞ�ƭ(���
���{3Rue�W�m�(j7)��ut��|I���?�yyF�T �-�?9��Ӕ�th�;�n<y�5�e��9��rMek%�A�PIV���+������
"�+�Ƒ��z�ot����"�A��|���Ϝ�"Dx�-��z��?��;����c���߯�����p��c�#L ��|8�w����5�@ǁ��������y��x#��Hˆ���h6�Cj�/���^���]���G�'d�6;%���s@����n\�r]�9���q�6d�6�v?����� Ծ��P�?8�������!��1=Nۨa�6Rڋa��V#b.TD \P��B�k�T�����OA� �o%��e(��Ό���a�|���b.�E��u%O41ʛ�����z�˻�%�*���r�nP���qr�cs�D��K��<SF����nl���g�uk̪+���D]h�&pY:�v{� l[����.�������1��˥�s��:
�]s��dB5��t� �}M��M����������4�~��!
�L��DI�h�b邍XQ(h$�p%˿$^Nq��E���Q9�D�hK4��}��tփFE� S �s��`��6vƙHM��eGu?��ق�O�>�Oڹ+a�ȢzvK1gCRv
����Z�����A'�W(F:A���TFo��.T3ODYW�K?<�
dU�(~ט��\�~�0�J_��P�a�1
���Ɓ;��G�Dr����ڦ~X�V?��p�mS(��x���ۙ1kЙ�����7upl�GA�RN9��J�1V�Ң:��ܮ�Slӌ�Y4|慠�s^拐�#��a`���'�"9�4�"�<��X�IJD!���#�jϬ5��2�c ��$�N�]?j��L���w�,���P��-q�2,L��h>6L.��W�i)+2���q��w6t��ҋl#�@�j/�R;^f��vD.χz^��֕8EF�G����1R@0y����hN�9��<�4..[D�$�<�G��L��@�{���4�N�H��e���9 e����/�K�,��q�W'nk�W��Ckm�	^�G&�)y����>���/|>����Q�b^/�G���\��s�_���S9�9d�����"x�-=�c!gL��FN��s�����؜�E�~|gU��8��7����Ф਒��1��!�����w�}���U�����`4\��-��l:[�Vu���*����m��κ}������[EDXT
�is��6)ڬ�a�/��?�e��3�<�������T��KZo�Q2��,�`��hŞEG�o�3E灬%������H7���v�1�Lϯ~���Ap�j��6���͵Y�˖�G�Â������a�~l���pAk~p������w*���]+����]h�)�Q��i� 4-���(�sbҟf[RFk|\�h�5>Sڳ~�d���؏z��k~��E�_����ui�J��r�Rp44�S�l�3����|��u�x���(�p�W�+���� <յAeI��̛:.c���q$�G�c�J:QZ؍���.�� ��$+�v	 8���Wt|��X>������}qBo�V�`nG��>�ug�*��N	?h
}X�^n�%����`�5(ǎm]Ş�F�c�t,Pd��=��Ç�qp����8�QA�x��5�o��)�+��y�tǳ6��[g�,�Yp��u�W�^�ZX��~�����h�A8�	�xH��p�.�%o�[��m5��_#�Ћ�A����lm�!��9X��L	¥V��ګMKe'��6�&�D`�P�F���`zO6���Tx���P�q0?)
[���|Z��J�n�mvΝ�9�9��}FD���B��bl�,�?z�iEs|�y&�/*ڔ#~%��)|�M�oR~�7� ��]�$�5��J7�^Y����g0}vȚ�^eRU7�2z�`�t�;�T&�����4��1{s�Yp]�ٴ�b}/��؛��V�ԁ�:���	~$H~�j� k3WX�mt����2�P�Q2����5��F�D��A�]�� �5���Z��d��-��"���6Jy���1�<���.J5$
��F�֠�B_�F2+�q4
֫�R�A�F��kU�5&��x�|�̜:��P���lDŒޅ#�._�t�K���<Q�u\��9�d�:�x����d��d�Z3j��H���/r�o���	�K+VWa̻]�V-��o�$�eU��g���f��Wd}������Teo�fp��0N�i�Y(�o7A²�D�d:(���58%LqX�̵�;��8;����7����<0.FI�9�5���BA3b��3�����h����h׵�ӕO����#_�o��)��p]�n���ٰ�軧W*��:����g8#͐��냵��FQ���g��!�\.��!Ggj[s	���脤���TW/N��́Ǻ���]v�tp:��t�&�N:'l�\=�����C�0���q�8(� ��Bf��
�'wQJ.%�C�-�����ȴ��:]�y��/;�$�*��F����)���o ��`�^=��(��\�|=~��#x����y���v�J'=�e'�믿����X_�E��%�@ �D�?��)��=���@;E���}������G��~r�[�*M,P�/y�=���&|��,9��h��Ћ��I����|-;/��cy��C��3�~�x˵+ ��kq,�bK��yW?�ˋ�3�B`�� �������b��^ᶨ���"��Y3�pW]������Mi�,G��t^,,�ů���>���n����U*�8�N7Q!��y^.�N�P���O��y���0��)�2�+�Yn�R^z���iA��{�v�i�ɼb�N\-j&����$�9�y'r��P~	6�c�(c\��lW��:��:�׵t�z]��rKꝳv�a��oqct��� �w[?�=�{��M�1J����q״�~�'����n(th�^C����܏�]XҌk�b����;}G�s��o��B3`�E��W�3��i�k�ǫ��*�G{�^�(pQа�8����|?����*7����ϗ�_�Ω�,�z� �g�Jk5����)�<�kU�>I�g<A�ϋ�:
eC
��G��TېD�~��]>ҁt���t=��ݔuMJ�BM�A�v,�=� ��6���Z`P!X�`��(iD+����������n��{ӻS�[�O��6xN$� ���~p
��y;\M��)zIw�=W=��O>���K_�|�;�@�еd���W��E%��+Kō��IC�9�d���g�	_���{�z�����s`*3ۜ�"�VG=|�K���'�|�J?����/:X�Vp��vΐ�IC�ͳ���S���.\9���õ��a��p(�/�\��U:�h��Ay_�V�~W#���׉j���P�� h?��;ir9P�Ҥ���&:S6-"�g�(�) �i:I��w�g9T7,
m�Ѻq���W6��)v�>q����d��+���Jv�c"�����!��8���̧j�4*hՉ���O%l���yu��"p=_�j��o���M~Q�\�/�6���e�=2ȩ2��d��A��YW�SO��Uޯ[�M9ɃH�f�ەYkOx1�/��S�Ϣ�CꖠZ��Ė)m�g��\Fg~��U�I={p��	�wPY�UQRa�����B��ο��P�y��H��F5stgZ�ee$�yj�Ӌ��nH$5E��ѩށA�(�Rq ��欫�wF�	1�
O��j�H��-؃�D��G��[Ժ��E�k�b����bIV�g���"�|꒬7�\BQ�@�h��u�rf����&[$����2�$V� V���Z��h�𡋕P��2~ʝ��d}��9:�.*�+G��Qzn�(�l�m¤��0�h?h��-
(B�~�H9��N�����2�!��%Q� Z���1f��Np�cf;(:M�_��}����u|
j[�<O�7�u(�ô5��
j�H�������M��7�]*��A3�\�!�9�:j[!a��A�d�>~��౓cL:�����Ɂq�tT.b�ٞ�M'M[�6�k�4 j?k�����;�`z�N��ʦ;:�<o74=�	V��P���x��1.\Y�Y��݉#2[wP�s�#��a�}�x���T�ݾ�A3p�������?���`q������f'a�
=��6��O�||I����7�����Gౣ���4�>>�����j����������+W��"�r��Qne���	�-F���YV�9����i֥�#.~����~:��H��}YJ�����39&�Q��"oK�txi�T�B1�3su9dW�j(�ld�2T������$h�ZA�������&�k��0���Z�&�d�,��7���Ŕ~������ʕ6Yό)-7��R�fn>j�8�J�Z�����,��x��B�q����M�	��t:�O���ꣅΈ\tK�^����Nt������9Vt�Z/���P�CyS.�y�[8rTϗ�vxh谅~ț
��a7V
,��F?�V�6����e˾����^�a��̯��3o�z۲eߚ]�i���j��������"�_@���S����iQ��Fl���(uŶ�T�o�j�΁�!8�ΩRÜ�'�W�����*���+�Qmg?�l�ȸ0?�y�����O~��Ej���kj��G���_/<��C"R���P��9kA�S;싮	#�f�X�[7vb��ʀ�^T�s<��k�'e�Wu��)ԩ5qT�k�W�F��Ԡ�E���պ�R�e\�+c�>���g{�x�_�x����F��p2��5��ȶI�V����ǪN�<L�):R�T�%|����/����� *\���:	J����ٛ��W���>���ay������=,"٦ ��d'Yt�x��V�H*�ۮ-����_������q�1�r����Xt�F�7=P�$'�&J����BB�y���Zϔ��_	�oT�|� �f9FS��;�*'�V�:���K`=���Mr�獭C ]w�;d�������t�:���n���\�'���ꬋF/�n��k/-�nFh���p��j��\]�Ge�%ve�K�f�F>S_�^mX_S=OU]�� J�!Gt�'�����s;����x�l��/����u�>�sϚ��1z�;�#�F;<4hc�@��T�to)� g	M����d4��B?ty�h��]d��ct?d��W'E�j\��,��<�����,�+$�kAD:���h羨�,N?1���CG�8>Y3G�rKĠ�a!/
G3O:Ub�>?͓�u�,E�P��w~�3�~�6����l�[?쾍�Õ/G-n�:��k�(m�)NQp�������E!��N��(>�~�}l�(�8�|��_�w�	��k����r\�m�8��ɏo(�����+�S�z��11���:V�������m:�����&� ���s���1
���_��S|Z�_;��4���k�� �����p����a�Z$:2*������?GE\~n0^)��Adt��֘R�"��9��;Y�N�;k嵝:�j�g7�����L���,ط��n[P�V��"٪rCf��ݹ��S@��@p���Ar,_ه�^�Z��{`�c�rM=�.����0^�N�CO>G݂��rt�I[��|�_�o��*_�\ؼ�4Z���;�����]��)h�;߁�~��#�Ðw����N��8�.;BN/���%«G�Ǉ��rD�"�q�;R�^x�l*9Ed�a�3@��:�_��K/���SX�Go�fݠ�q��ˮ���B�u5Cf}(�W�ϲh��E�b<�KM�LI�በ�"�Y��֜h�l|'p\���;���P$#�3`:���E� �l���u
"��p����:-���qi�^�������r��&;<�@�s�OZ���B���-���iiT��e"�Ne��#9���R��>�K"CD��^q��\ә��	:��O�q��g`k�V`�	Zw�(nlt��Qړ~�mSCԊl�uO�W��=7,��<�a���[uX��k?��U�@YO����}�iM�*�� J[[�[{��oo�ע�P��ڛ�vZa��9[�7ƉO{�g�
��=�.	P���/��9eu5�jB��7��r�ոb�6�G�G��]��P���\8���s��B�,����E�X��x��`�}e<�]��,NǲNb�!����o%=(��,��2�V�Z?p~��3�l<(��8���EHM|��*E
^F�<�tlǊ����J��.���Tt�F����k�n�·5��;�e�a"��[+���}�E�xPξ�u�V�d��M-n�ֵ��!�����`}�����?�_����GG9`�[�^�~�t�[�ؕ�}7�����q^.��ಇ���CJR¬_9y�����Ũߥ���+o܂o��.��u�&PBUʾH&��ve�̙EFe61���A��8�m�1>>b)qZa���p�q_V+�'�~�z�3ǧ��py�܊3��o�ӈ+3p@�z�C�qPv[!_�Ћ�|A���n$�k��R�C7�N�6j��o�H��`�v����K�H�󂮑�V|���{s��M��禺��JdL���3�������ws��?k?΂�M��6n��v��
���>�lj�e�Y��y�
s�4t��� =%־���s<��(Cw�x��5��nM��e�IW
��Uɿ?�L��j�d}e��8#P6ܖ���p������L8F�`��c}�t��٬U�ƤP_"��؏
�h�tKX�S�\�*�sH�.U�9a:S��C,�> ��
��6Յ#��38e&p�S������3�,� �:�ί�Y��]jR?c�H�3�����w�9e�P��r�~PC˜N6��FJU�8+ڈ�6�L�NÈ���S�ˢo�
ڎ��EF�q��N�B!X��,ەU�Kh������u>Ԁ�-�?^���!h�����Q�2}�F�6Vu��E�(���Ew�h@�?�[��5-�R�+GQ�v���R�O��?y]?����Q���%�#����=>ȸ"|N�N
���'h����4be���J˥��d"<����^uTC��w��yG�i�W^�v�C�W��6 gKZ�V~�:԰��j��ݝ�0Ų���|Z/�7��m-�	�TPZ������e�c2���nW��n+[��E�.Q�2 4����uo]��lR��Ft罦�:�|�����Q/I2~�[6Yā G��GZ��?��,Sf
�
n����]�]iܢǭު�*�2;I����7ƹ�;��3���<������;�qi�s{"��G����,S���d�h֫��"9_IW��f=���eZ��?���
�u�n@;+1��=�]�i $x�Ӑ�LA�E��ܯ��Y��{^Z﷾���}�2ps�ɨ��9(�}�����\��]�صM	%�UtO_C��n�8�]��Z�g�R�[�Wp�NYjRP����,|�%cޙځ����I}b̛ܦ�L�,i-�#�^��2.��c����(�d�1����l�ʧmPy~n[��-2�K�B���n?�� x�е@��gJ�Ulé��YC��=W8v�d���xٶ�.>� �iUeB@���a]�ˌ`k��
�j�k�6��c�o߶� bW�f-�x��hOa̔3��](�j�v5f��ngB�BC�-_�d�T���;�N���r�ơX4�v��Ts$8��t�Z�Zv���L	�7(q&���By�1}������K�>b����u� v��]�:X!='OF^�	���B�HJ���N�%���55�$����\���[���� x�c��2Ά�pщ˃:8�2�6/E��*�3ƨ�$7���B���}`F~�+|\ń�u��Ǹz��j(*�¶1i�9�LR�Sl���~�^�(ćz�er�0Ý����'��K��|��_8Z^Ƈs@E`�޵g"[(� 0|���n���s!s��Ͻ _|�k�����dqǏԆ�#�������8��O�Z�
�s�r�d|ƞЂ�W}�>���G!g�鎎շ��d��>��{Ԁ_!�FB#��z׸�e�r��y%0�q��:�<é��� S����i������'h�tV�O߿����
&��h� a9�%�J��TүNV�5PF��{����.�眔MA����$����<���@�d��u��R&&<���Xh�B�9Jk@<n�!��)��ط`/?k�_.l�1�v�Z����']������������Y)��0ɒ�2��^y��u~~.`(du��Q�OMO�l�k�w]kC�B��.�|5��N�!��c�t�u�}�v�@����f/�{�g�d���[ׅ���{p�*��p�fg�[���3b��u�[.�� ד�hNI�l�kx�����?����{�u�IJ̕�rH�N�;�#l������Ku�n<V.R���%�PO+R�3��GpI���jc�ђ�}���=gmdN_خ~���<�#[�F�quu�e��Q�r�Tg���. �(�\'Y4�\ˋ@��噱f�V*�su���'n�?�𪌲����8rN\ap�����t���0�����5�����s��a2������8��u����~����	�U��k��R٧+%-�8�9eA��n�Z��SZ�����6��P���Tp4@E�<���;Od��0���?�f�	���$�-�L��d����HAh�T�iws��8��, %e �G�Wo�zq��D��o��02�t#�*]:n�Z�P6Am�Ǔ�,�HO���}�����	87�0�~�?�zwW%GΓ�.�9���ݒF�ey���\�-K�~��<'+��O��Q(��5ah!��㾃�}�o���WY��ZG��^�~IzKrdJ`�����`���}��Y�U9.�?�O���7^��^�Q,�yq>�z��1x����9%xΜ��xŠGщ�Љ�湓��J|�
�����빮�����ܑ����#���c钩�f�'%������rOM��V 	s�8��m��w�x�)E~ZʙM�Hց��7X�>?�c,�Ϯ������&�x#�< ����k�J����BA��ҹ�$�ʀ���u���r �i����w��O��^{n�܄Я!�Д���QJ<�&��u
atE��'�J;:_�N�S@z^�̧�����]e�ӂ��{�?сK�4� ��OO�Z�@u��~��s$+b]t�B�UqW
��'�
[	'ϩ�p,G�!,��s�zk{��Y��C��
��x&Tux�EԞJOn�:�+�m,���%S��۷>�:Z��5V�{���.�����3�En�ԁή,&�.�/},l���W���ZwZR������U�\?����O�z"OKY&w\���Ø�*�`Ψ�s�������J�����]��:��E��py��X��%O^�?�����^�kȁ���!�o��_�	���[�LJ�+��K�V�e�|OCu�g+�_,��EZԣyJ]�9��w�R�GLߪȒ)k�^���bU���L��U�����|��5�Q_y��u8^�S�ƅ�WT�xt_����ӓ�{���t|��K̟u.����>�=��Uo��O��'͍��qN�<�`�����>���R��������z�+���Xb�6M����;�Q�&���ֱ���:�"ڣ\DI@i�W�w8X]�:鮶�Q�O1�*�g,��	��`���N��Ne�RV��Lux��K�ld.����~й@j3N~o~�!�\c9I���d�P9���|�������������)8y�&t�N��8���I�i�E���*58��u���6��tє妶US�4���A�k9~g�����f��#�Q�kd=S�� ����Ѳ%>!�5�IG��B�"�Y�r��|/pcsf��S�.���gV�:9�X�F�^�V1^�	>��ߏ�f�t.�p�BN�qP߯����mmD�p��k}�h=ұ]�Y0� ��*2U�b�|�jo[e������O�7��߮7;;��=��	�s|�ۜǰ�p
Z��.���_�
6�:．W�ݩ߮�����	���|���X��c+[����}�G;��;�v���/��%e=�r�GQ�[�z.�

��M��&�������P�?�~H�b��^��E��������(�l���2_C{~�����ф�E�K�S�����ӀF�����'0J��b:��A��8q_k�GX��2/��2���\`�ӻK���� \�r4������y|��u\�~�?0��Ϗ���g�A��!X"��쟁������"@�F��@�|7<�jI�hM����x��? ����_}=�����]&�D�}B�d��7�/@&$e.U�(��@{e�t�J���܎X����ʰaN�m#�ʲ���.� 4��*}�
�>�2דb�^L혫k�z��;g���J���B����e�=�w�`��k�UN׻X5k���}�8�PG���z�ў��������V3�9mt��y�F�Ʉ�m3q<�c�;����;���㌋�;k���<#j�!½8=(p�={T��H�,���?���<��X����4�6���]��ND��;�Be�P;7[����q?	l ���BHʓn�<�t����.o���I���h�D����)&����?$�:���ZÃGx����d<�B�c�:��͛��W^��rI礧I�]�դI_嚍�(�+�KB�_ݨ�?��w��?���������h�MK��y�c�õ��kɀ����d8��ݬb8g��Y5:ʺ�ܮ�ɗ�:T���h����b/�k�Q�L�.�K������״�iih��vs~U��:b���0�c� ,m}��������t.%�
�-n�5Q�n�k	��W�#we	�l�?��w�Cϼn�1�6ɮ	�Ѯ��E��W�W���*�i�R�m;�y~R=�4�������� R���P�k�>\N����mZ����:��<��|cv�d�r���n�a��M��lnCs�ϰ��u�Q�Y�ٕ����q{h?Cp�5�w�j;:[�m�#6�*^7�Z%���!'s���S����C���E��.��(!k^&�G/n�Pʡ�ɡ=dǭ�=W9s;�{!/@�le鈽��垼�m����ޫ2���T��<�[���-���мPȋXH,� A� 4@tc\T�Y���1�h_L�!�ʔ�y"�z�Q�;atӞO�������I.��{��!�c7��t��l�Ń�Ҥݘ�{��珂qH�I^�
�����Y�(��|=��8F�wz�E�������c�0�l �s9��8'��o܀�oB�� �����ȇ,��/
ڰ ��.�Bx���6��� �ݎh�6
�c�5/��C����j���N<�_�>K��7�XP�-���� c��+?����,��
�:�٠\�0�s�M�D;��e
���w���ӓ� ޺�j��	-������͐ˎ�Ly��[f���DӗX4.d�F��/�2_q6;z~V^d9N*��I�I�i�<�u�� �|L�[h>���lp�E�ȋ�*%��N|$ܯN��L&'lau��lYDG�`�Ƶ�#d
���w�@��
dUj���[~^Z_��n����]{T{�Z�v�  Ө�82O�@�ƃbG}5�_O=���jf���^��!������:�tX?�}_�S��ćmz�R���}A� �cp��!��U0�dN�F�h8�vY_�Ʒ�����#��1��(���v��R�` �@��l��b�O)'b�3� &A�Y��MA�AW}E"9[��Ӱ�����/���`�r6��~���'�����k��w^����t\dST
[0X�����M����L8������2�'����뗰�zF��c��:IPbJi��=E+	Q\�'��h�M��4܄蜢,_�Y
�עčiH����f�V���Rìқmr�'�����c��P��6A���}�Hj��1�:��v�Ϣh��u�[�lc���s-����v�M��M`C8�����GWu?��sCa�:���]�?�ưs9���Sh]m�'-�_($)L��,kB9}U�N��M�Vⴍ�Rh�nb-ě�b`ћ�j�M�m�}ʥ��;Q�ߚz��l5�8_��,� �g������iSr�|lʐ"@���)Uk~gū<M���TCpf����a@,���e��6���(��ly�D�  �Fz���k�Y�'zִ�,y���nTZ�1�W�ܸv���E�.󒬦�������5�zd�?�-"O�� ���H<TM�x����1��Y)�:*��]�=�u��{�'��'��1O��Ϸ\[��n	/�s���q��B��Fr��Q��BO-Y�2�\�i���qO_S�l ��j
cAFS�懱$.slC�׋&�@2�\��]~gA���=k�vˉ�[BՎ��2@�jps
��h�\J�z����!$99�w�,������\���)����|gI]#6R�r��ߴ��hFos(�R� ;%���kC��f�>�&p4$r�2���|u��n:�wa��s�N�\6�N.l�}uX�	y���Lu�VQ���9���"[�*�j�N6��YN���u��r<a����<n����M�7!������/��	����g[��R�l]<�?Fv?Ux�놌ʴ.�O��`�$Z+5[ݸP+�#�ˋO�|r�e5^����Ѣ����nmz��h�G�1�A�5�w_���ϡ�$��"to�>J�g�N>�U�`#At�Y���P��R�s��Th����U�h.�Y�W�B�IX��O�={���p 9M6��N����b�������?&��|
����\��R�t��:��⇩ܤ��Y���~�Ex���ѫ7�����,8f������JL��/ryi�I����;�oR�r<�*�����Wd;���c���h�#�q��]�8O���Ѫ��V�n�����F��~вt��8^0��ferLt�V�p�P�R���*".`��#p��#X]]��$���8���	�����Y�u �l.9V�+�er�����U^ז�țy#�Y��bZt�=H��y�=��]  �t��/��dGa�߲~�m�˂���b��Z� �H�K9?�eȲg�Jf� ��q��e`\M���Btp�Dg'z�7��Ut�K!>���08W��+�.ռ���3�^�ۿW��c�3u�����5xL��*������������`��3�*~7�כ�S����N~hs����Q�a2K���S��;m���e� ����Y*hy�&�h��&�zfR���kۙ�d����4L��fj���N����N�Vt�yY�C�L�{?���C�3�D{6��u�8H�Ȑ��e�S���ǵ�eX��� W�=��oc���+Rv-�A�M����@���j����Etӝ�H��s=�h��Hrdѐ��H��E`��;�4���5��Z�\B�J�y�����`�����J}jav,r8���BܗU(�3��\

4�7�ZTű����w�l]���6#��\�T�,�F�˥��Z���d�
�|�X�c�:��`JQ��?ⴍ3~��2����U�g�;a҄�-\Z߸�Z�Ʈ|G�����~ܯ �'�D�0���Z��D��4�|���:_�>�`��f�G.+����pǯM�ME���y~7������e��8$�.L��EU�/�#�(�6��52>�R;.�\����d<�PZb�����3��r1�K�H����Q��]��ج�����TV�M���I��;�Mp�P�2g��k.T����&�Uw�2*�	�o��ŵRlk/�9�aN��v�g�7�vC%��ڨ��s�B�ʉ���M���W��"D�Z$�+�ȻΨ�pPH ���L�D2]���Z,�c�CG����\��Ed���1\���؉��٬r��G���絤O�s�鍮[�d�ϣ��돴�8�Ȯ=�8�hF�<�F����@�h�S%��=%q렟BK���.Pˏ��%���|p��?AɉnBs��+��C=^�wE[�%��Hp�V��yF�InE�Hf[!��@��4�̻a�z���\�5!�!Z {&u�
 �>���e8T��Ur,듒}����~�fu�(�%7G���Z�������#�0釶E�Ȋ�^:l0����T�������~��6AS�Ug��=�G�RפN�]eG����m{zÞ����C�w�:J�.<e7����]��A�m�]Q_���i_'<9�Z�����M6��6�ӎ3\��9-��-��@�r��a�Cu"��#����H���G�c8=��	��8]�˾A�DK�(�|���u
�E���u��Sj���p�:ĎE�v���xGk��Z��ʞ�b���m�����%�v�&w��>�2��D���$=�w�[�M��9wsu
/�q+O`�?^X�']<�MC?Px��/2�n��;)u���5<��w��w��Hv'��m�l��?�����5���(Y�8�D� ���Iݵ���{��r<@�djF��4��	�^$�����VW��������nϵ����n���ey/h}�y'�<#�u���{� � �Ŀ"� #}��)��@Yӿ~ř�OJ�g���s�R�cr��n3`���E���z�w����&� �ݶ�֤3zZ�5:~y���'��U������FCmk�3����7��"C�Um7�O�D�~���t�~a�Ut`�F�e��2@���.H�l�k��)�3LFI_� MY���FT[ͣ���0�O���3�DR�6%ȮŇ�
��e>Zew�w����Z���\��A�(�QY���o���*z��#�=l�����m�U�z�s�}���̌fF� $$ !�d@b�@�!���	���R�$UI�RI�rQ��M�8@�$2���DBF҈���������4��w�ٻ��{}{��g�Ͻ��Κy���wVw�^���ի��b[�7�R9����\H3�'4��eM���<���ј���Dg������D�~�-R�Ժ�tҢ�� ��������zT����t��Ʒ��~�5DJ�ř�0\6*q���(9��%�ץ��7'��>ؖ��`g
r�}�.�,<6�]c��8�3��2Q8[�`E�i�{A�W;�x
k]���Z��g�O��������f�K��u���y �F"�w�!�HT�r[ ��b��Tp{Ђ@�4�p��fDq:���z�'�rr�h�}��#�I�����?�X��_�Fȗ��;��y��
�5v�^���㡺�;Yy��B�A]{Nemb����}1T��-��:4H��$b��%�@՞ʷ�{~I���$�ν���y{�5`J��[�sA�,��_�4ă�1��q�$$�rH��� �>GT~R$�F�֘<mT%#-
0t8�h8�Y����Ij�dt�c���[��yf�)oN��#k`+�O��]��i��!�)���
/v�xܙ�N����?z�V2���5�ˢ���(?��ţ�-�Aj:��=i�J*�Z�+]�G�L�+�-�>��.������Q�r~%����h��Њ=u*k�	ʨ��Н4�EG��Q8 j���'�]�5�����A@?s���⼁jo���6Eŀ�xF�+8�Ǝ�_E�YP	�O�t�������4.�F��=␨�˱��_Y�z�#p
�9�c������Ͻ�����G���E�j�!�G���*jr�2.���*�A"��I@��J��Yf*��Y��;��C�*�3�{@�#opu�2�2O�!r`����� ���A[��Ѧd�Lsˋ�6�(�*c�Wk0�o��\�+ZeA�&��2�״��W��or�(]��,��v4���d����r��/�a��e��eꩲ�2�s�` O0'Zst��n��7�v]�s��-�i;��S���C�9���P	������� %:S<o�gOr���6��N���I�'�%�J �yèi8�\�����$��5�&	)0�:���v�U�M�S�x�?^-��3��f9��uٙ^��YtE�N>�m�6ϻ6� ��|s���e"�/��C;ť4"�a2����@��vx6�+���,i�^��o���o��t��O���������O�U�F�Yt��=<q�<z��h$�;�[W�ұ9)49KU}�;������=%�M5?pp���=���N�+/���n�n��$�tE��'1�`��E�t��4����	�����ډ~D>��K�E�Nm�fN3������y��9��'<�����kq['��BG
�̞� �d����k�FƓ�
�p���J@�mlp���y�k�ϡMv�/��gs�v�y�΅��[��U �4'�4�Vge�֐�'wG���[r�I�1\�Y�Scr�`Z[��y�˃�:�ڙ�ruIW�Eh������W2�S?���B�i�Qs)�[W*\m��w6�P� �h�����2��܊���U	$$�h;,-�Ԏ*�jG��]^=��MI� ���U�@�zD�)�u�%�@�^�YL\�NC�G�����pi�e}M�C��K;*BF�9Χp���)>�kE6�]����M=�l$�dxMo$�p;�]��^l��v��_{���'�������Y������Gc��,Zs�5��8�Et$wr=��4����(
L{.9��֙B=-5���DY�^�D>d������CI^��Uc�Db{}�a��u�vq��8�$_)��낉��O_�ȹ��kT0=2���h�$bHe��ĀeifK�K�嵦6���D�R�������#�2�]��
�h��m������;W�UN㊸�i�no�幁:�`�t�̳��(�q��_Cu�۳��֥��x�ju���x�ތ��0��_��W���-�S���� ,�E�©����:��@d��e�e��"���EV��WW����Y�6��ݚ-*K;��b�)!��T�?�x��?2����V0p��fBI��1�^,���4N��ӃU�}o���'e��-K���fq���P��P���(({Q�����^w��N�Wn��p���nf�x�'0��#!��1v�s2��"���l�P:9A�x8����p}M�Y�T��x�����t��tyR8a,�vc��R�U��i��t��oR�$\��<t=J� ��<<F��Ƀ&�^d����B���)N�Esԩ$�Li��І����G�K?Gik��Vͱ��E赲ڀI�N���Mߣ�`xR�Wދ�@k"C����yPa���i�ک���dV5��{2���f��:��CK����+�x��C��X&����rݤ��E���X�~72:C�I�e|Ju�S��:�H7��6y�.{�Zy�'˗�(�zN�ccև�K���*Y�ٌJ�(��&<}�kD�T5ky��u��7!�C�Kr_8�Ӣ�NCg:��k��k.y�64��qU���Yy�H,!e��t�u�>,��j��l�N~r�� �%9�:n�xM�!��>�j�،�����-8k'ռy��޴aY�����vv*���i;�QQz}�QG�c�'�:O���� 4���"';穯h�)���ْ.�WBd ���?&r�
-�}�[��Nwr��щe��Q��Er�m��(�������0ɣ
 =�ciė@;���OLD�N��l�24���l�Ѝ5�#�=�iF�xΩa!$j�yD���MP��Z���cH�ŚE���wU��wD�!�nU��O㓣b���sܿi�5�m˺D��t���X���m1�y��3��)۴S�t*���0�2K�x\���ԫP#S=;��g�r.y�!���Nq����>҈�4�Ʀ�ӗs�
�)rQ;|���M��s�|��Xi��߈��r��p9���r�\�</G#Uf�׬���r�_7���\�,J㉖U}�������9#��偆xQ*/��A���
t0F����9#���~ؒ�Fz�v��b�����tJb��Ё�����_(�u����&���`�����j�9<w�ڤ~ �LR~��
lz��@u���oO�K6�)j�Ӷ�Զ=�� 6� �^�@�3���t-J� �(�rd�.ս,zd�����+|��Jr���S4O�E�g �H��0K�ʂ
�'�EO�Z��'�1,�G<�Gv��S4|�@�{\vJ�{��p�GlD����G�:*,���*�2T���ʷ(�$8 ��c���=�ӆ&��N��vh��x_Z%%9��8�$9:�<��w"����m, ���(O\D�^�9�t��|e� �;|ʔ;���G^��y���K��|�'g�E�i��M�P޻�[�O;�C�|Y��ץ�iQ2ֱ�O��Z�
0�/q��<����Fӡ;�C���?��6c���ƘH���Wg+$m���R�����4Ȣ���>�X�KyignL�\y�e� ��('bLB2���jhL�M\3���D,��K��Q��%;�1�k����|'
y�$X��c!��=�G��qc�t�jK�[���!r��s�'(��2�f�cU)r�$!R���zk0X�	�=ړ�qM�p��fn'�d����g$�^m�;�lJ'2r��@�u��Mt��x���da҉D���	gCZ�S+)�D�&�xԿx��#�>���3(��t�p]�ɓ'046�AR��,E����y8�0���l�$��4G9(ѯ�B�	_ѵh�Z��aZ���J�FY�k��U�ݗk�?g�م��Xp!Ì�t�&'vn9���Q����!�E�?�K�k}���K�%@S.Ӛ�~"��.ǫ4R�؈�\��h;R���#��)0c��ne��A���N�`�����f�i�M��<��4�۴�bR�L�Hu�5��c�-r|��Lj��Y_`D5�:B{P��U����)�G�E�����pwc�Wfm�z�k��p��eww�A��^?���ޤ���R�j��i���܆Ʒ-ѻ(ߤ!љ�B��D��A^ˈ� �����-<�.��a.~ɻZŃ�4HH�	�!��Dã'i�PZp����ɨ��+�����8�|��<3����g�4�,�]㶰���o���(���s6����S��}�{V�28���
�϶.�4�6�RH�t�t�.��W@�0��	�Ä�JX$C}�^��<��V�j6���'*/[��9��2dq��w(��͌Y�q�* /�2��t,�nN%v8��y���8����է���ܥ��s���3m�Pz�m��6�M.9R��u���G�R�W�N57-\{���(���ډy�eq��\�E%!�k'Ec4'��)���?%Yб���,6�Z��U�#���j0v�1�7fL��i^�dL[��b�dy �������P������'��Vܶ�����>�;3*��jG�j�	�ge��N������\12���!p5(���-6h��'�ғ�Hɰ�^�-&a�a;ȚA�S�i:+��x�����EI�еsކ�B=f�ԣtY�2}��Ri��	�5ZeN!�%�J���@�հ/͊��3ʍ|��[�{r@$beG�u>��hpwV�7���e���U2��s�A���]J�g�Pr����t"��K�A���0B8�d{V��4N@�����]8����݀v�
�BG�@cƶl~�64x\�<��@Q�I>��?��=�SG�=E�s,���}d:�-$:��Sk�{���1�H�>��$=o���,��<#��&9q�^�}17���JS���%�����'�����(Z�����7��q⃅;M���Ж�d[��e
�����(�(E��s�5x�)(>6������Ӳ����dc����JRY|�t�6�A|蓽Yqp��T�64�y���V��RH5
!iN���)M�ΓbrZ����y�}/���r�_mi��aؚ�7/ї��y�ζ��X�s��� k����u�;���-L�� ^Gl��3A+>	���Ј�I���:��g��7�F��Y�-��aT�1���&1z��ܹ�č�b�~�w�`Crĥv �o�e�Je|�q�P������{IgiX����K�vw>ʐ���ڴ�����O��dLATmt����������U�~$��i�_G��Y��h�f�E�2�N��>��đ6x�Y"��Q!y$�]��Ӣ���W����މ]8u��":��$ec���Y�vvfp�i �W7i¦�hL�R?;5�ğZ�m'��J�I%���"g/2"Viø�F�t�bj|5?�]��L�{��QrxA)zei�1UP�~��g�j	'����*p�|c�)�^T�#g�����#�l<Zhɑ��@��y�g4���N)��Q��.Eg�� .1C[�* їL)��^+��ZY��N$Z�P���2M�s�����]9�V��V?�13pُ"�/�W_�5h�Л���̡:%�M(#)�gމ��٢.��ҧM\�B�z�q�E�M�trE��(�"��}������ŕ �о$V��eCK���=�[��1p%^�!$��7H�AL=	~
��A:�;�O塳�%��HBqi�����hqQW�7�!��'/v���ᵑF�q��u����n�I�O�mf�c}�e�|�b�?�N�"��Hva��u���0���ڳ�;�j���ږi���%���_lST��p[9t$Ǿ��-�P����C8�P��W��jT"z�(�Xn�Y���|v��8�2N��Gf�ͽ��:k���T��c^d�E06���t>=RG��\�@|F1yNz?�0h���Z���_����_�������F�mJ�&܈��.4(n`�갔������-\I`m!I,����=�.9�^s���)����/*�^9��=��&��J��}��&�%�B��Hѱ����z�?:��s�:0,#CẬ>���1Q�>REX�I��d�<�]����Mǐ0��q!�Px��<5�h�|K*L2܉�M:yh�4�+xh�9;͡&�:��E�lg�C!�� ����p(04�i���W�P��ԏ7υwx�*.�qxUB�>@��(6(]�*Q��$3x���(|;	���g��2r(�N��ko��=�ȟC�x�,�3��*��ڞ�8��/A1l��dqK�-f�$�`?1N�9_��:VΦ6C�6��hi�K1ְ�H
4P�J�ω@��T{�+�u��@���6x��A>�l����:q���ί?���bX�Uë{���
*��<��)��~��X�ב_�Kp��`/m���o�o����}�����5A��fM8=w����� 8���*olG�s��|����B܍�'^K#nzQ��%!>�n�Ȼ� ��{/�4�GgZ���F�G��Hx�9i���:�Kn]�\��qR��a���<�ʁ���S6��x2^Nk�^Kb�.V�A�<[c6UwiM,֟����H��$����Z9�TY�J�č�0�n��y�����
�eay��G*�"

-J;\��^�V��ۙ]?�s��X'��h��ЅFɒcΐ�#t���}rXH_��4Aȶ��-L��95���'�s�@�J�X�N��-�i�
�#��)X� ���Nޕ�ӫ4��/������ĺ[�4x�M�ʫz�:��,ɦuZbPG
o<:��v�&��2�Em3o�Lw�%�,+{`-�hy���D���]�I�NRit���͂�{�+EŌy��r��m�c~���h�Jʽ��Bw4��u��5���A_}�twz�R�Kq�(?wt~���p����pv�"�Ա��F\YG,Pm���'�~�����-�<.^��U7��=sǮN�S� ��^Ȯ�
����y�̉�0�o\�.i��{�LӔ��3k���Hy�tz$�]��q�H�
R�KU��礃H��}k�_��1�/1]Q:T��-Jr���6��1��&+���v�d,�Q�)HCY�7-�_/�|5������J ����b_�#T�g�j'���D[؊��5�F_`{#�L��PuUk�E��R����3�5.���P٥>9��-l����u(@�J�����d��BߴL9 U��&�a[[������	�����ՆOB� �v���QNJzG�zͣ,`�t�c��CV�_al
v��['�`!\8r`��,�Bx�eش�D�$L��A�{Ћr��~ˊ7�ʉ]jz\;�nd�E��i� 3"����N[��`F�l�
<�8�8H�/�la[�mXē��
��٢�x`5G�?�ɂ�:�		�	J"#�6f	^gĄ�,�q9%�{_;%-�E��b����T��OS֑R}G�c��AڰS4�P���רQ
o�-Ʉt��sB2$M�OjՆ1�)��<�``Lj2�^�������{
~�1���c�P�>!�TN���[_���/D�` 	F�&ދ^��hp�����(�	�4�D�N�I`ӕ۠#�<���;	�z7]��T,�f��^�7p�}���K�+�C��F���N�W�E�P׷ X�AMVu���+����F�_ʳ�N:���K�M]�~rRN�����O%��P��-��&�'�>���\���!̜Hav���?����8Ѧ�up��\�,��5E�9]j$�	�v��߮�yC<�"U5�a5g�=�X$s���ȏ
Φ�~2�17���:VI�r�*z��6S��J�#��|w�Bֳ�o�.�RI��4�G}"W�Ҳ����7P��ٸ�*�PrT�ke=�Țx��
�ʁay�۪`G[@��ʕ�yt/�2*���`4	,<� i#Y�ɖ����ix�e�\E���˯ޤ+[�S`=[�A��Z�y��w|���^Z�Q���5n8s�����w�e셺m�f��t��Ґ�1đ@�HVp���f�q�!��&^�B8�p��)���!��8-+n��_��8����x�I��t��m1d�k�)E����������x�q����X��1;�Q;.��Qe��\�)3;'����T��<���t�O"��y�:}f*�	�t�d��Qt��T�x�Ⱥ�ʤ��߶�z7Dk�e�[%�e�Ud��m?C��&L��r�����zA��J�P+�@9+�]m�x�`��D-�zc�FF�x��CIh�舐�ߕL���u~��P%Ad�Q_y�d���6TH��_ޕb���%L�1be���Ş"c�ʉ7C�5Zj�J'?J�~e��1�6�4ٮ.���p�`����~�����i1ƍZ��  \zN�80F�I��C�������qGa�F[�����7e�3&��%� 1���S��	��20l���Ț'���y26�5=^K~�l���2܁�7�-�ˍJ�沂�W��8�E��~��	�jő`����s������Kʸln$� 	^���¹�=x���aww7�T �&�����%��	���t������.�X������B=��� �q�/�3�����:�Ӯ�T�ޕԗl�D�Ȱ����,~�T"~RtV��rz`��Ʒ��NGFA��[ޛ��Yj����6��:��\���}͌ʐ�9��x(aSƸ�7�z�[Gm�Z�>
YNL��/��_�î�I٤Tu��r��z
�����K�L�;�):����ʠv��Տ�+�ߕNL�����)�(�ְ��-,�Ӝ�6��6Z�t�-'zZ�����������[4h�p�a��(j��Ā-L;��/ �ޚ��:�B�i���$:��������x��8���$������S�>��'^"rW����^��u'$���K�?���}Z�`�]l������o��g��؃6\��,�6F٬��~��,��{�!��v���{h����y0o�x����xPN�=xֵ7������'�����/�	�v��M��C:p���	A=��qI���"Q-��V����/j ���t�Sm��h��X��}Hg��%��}_�k�\7��4D�b��\��M�-,���e;0Ww����B���4ę֪��}��w2
����F'[Zo�d����/����M�����TxA��SHU�#�^\�ʢ�ѕ��mGտh�ThD�{@�	�6��<�H����r�5�(�!�Э}�m���I�qΞf��E�r���J��8t��b ?�������%Z��`�maW��|C���x��cmK�~�O�e#�����p�!S�l��^��Ӹ�3g#�O'���!���N��� 7[��5!���O�����
��O��h�[���Z�	���*O0��K���(a��T��3�i�G�2�$c�A������f�7��ٿ�^���%y!V�E�!Zn�<|Ʃs������}���Y77`v⻹k�����).�8hae�2�b�P��y7ߚ6|6��x���V^p��].�,�g��������`7�ܫ�:�P{MIC�8��L�җ����T�2:p�g�C�����(�m-o���S�B7B*�X���|��oP��)t��A�c�7���)m�8Z#�tՁ�$Yx/�.��N���,�:�F�h�7��NE�i��L�9l,vޠJq>؇B�\��ͅ��6�E�o��:��A��0�f[��tXvތ��������K�B�*��G ���^�]Re���������V� �`�2@{R�𶓾���ċj[�)��N/\��jt�f�ޓա4���zU�q|W�ik�)I�#�i�!��n��}��.�8辌�M�9�j���'����ę��e�"nh�=*�	�B�����N���ŋp�7��t�����+�ẝ8!D���Ӹ�����a�G}ǡ�w#��햳'��7b��)� @������?�u�;�ە�����iM�4���e�8z@�/ɮr����x�D�C�Y�!t�Q�̸gB�v��Z�AG!���Y�[�V���,�̈��)�$��@�U����O�E9��}�7�*�+�!���d� 5c=�:�p	Ju����r�lj)<j�zl���[z��$�R��~���o)˓�}��v�����ڎ�dk��[#҉�؆d��!��Q�}Vr��BR����Y��wɴ�Р�\�Q��R8p��th7e�7�D��Nd��(�"�VIHA�E��9N�$���ϟ� �
�\.�� 9��y5q�-l�h`��1d��?��^2	J�A�[�����ď+��V��#���$���3��0�ڸJ�Q�I�)R%<�X�Y� `��^L����/���s�ɵb���l��ވ����֠��g	�����B-.�\�{ �E����2�Kܟ(�v�W�*�!�E]�'�|'�? {.�54���9��u�1�ǿ���$|�ɧ�=1r�h�`,l��&Z��1�<����xz/H%�<�0o��3�*ռ�-.��G_�<��/�N���\Q��=`�xR&��w��wqm�� IZvZ��z�Ȉ��̽=s�N��iZ4Ұ#�2[
*�$x�y�b9٬��i �)�43jz��
^l�,�3��r���"Qbw����mH>�:��e��OU�ؕ�T`�љ4�)xi���Z-�TR�|Ў�وq��~$��P��NL8)M;��|����u0�f��]�N�&������C2ʢ|[���06�������Q�O2����z&�	L�>��bob�p�8��O�����2U��t@M��a����ǴSˎ�QL�'��s	D��� ��G����7����;��i��F���Q/�$����YUJ��Ծ�r��ED�F�v��_N@4N�����$�?q����Cp��s)�wt��
��60���7� ���>�w�?w`�����,:M���a��<'<��؁�s�e����#^�����)?�����^�ï�kv� .�O�rT��܉�5*�pq�=�D�j.\o�Q>�|	��8�����Q�lN�ˊ>�K���ۅ��{@���>X�<�\U�5��1��¾���Qҋ��3</uѥzYP��C��[��S#=-룠Ak��t؄�L����|�y��Z��H����9��^���Z�z�幵G�]^���c�2�m�67�S3Ԏ)8_��B��l��d��bza�<���kG�z�5N�1ʎ�F;�W�ު�?E݌MUh�%~G�h���[�c�N0�HEv-ń�PASGWF��qB�r��h2�u�Ã5"p	R�H	&9�Vh`�Xw�^T�!��n&z�iR��>�?���f��Abt�4�!\�[�:��6�R���(:d��P�lZ���mj�)�Gڿ�cSW�K=����8-�mpm��J@w�d<r�r��������Zm��o��E�S�'�s-`�2�E�N�D!"�-_�k&ذa#9{��O�Qg"�*�ٚ����s��QO�5!�����M������@�,�i���̘Ŀ���ǗO0y5�P�ͥ8>��3p�CگPI�6��{�S�g�r\�����I��az�G��㛞��m����o��;�t�ÎG���ҝ�L��y�'�E�b�K�ј��u)!�F
�[��8�8x�s����WÙ�,m(G����#e��X��w�+a*�eJQq���RK����P �F2C]�6l@5���.�>�8�i+K��h������\�暾ל��DU�K��1*T�?��y�A�G�K��?$8�Ӵ!@2�s����։^���T���_��J� �{Z.�@Af�a��d"O�ҩa�Gו�y�&=+�� �C���A�L�w��֥����!��#��G�_J��oV@O|�/D'-�i='~Xv��=�#;�ڐɱ΁�FU_^��A�e��_�'Vl��-ͼ�B�9�A<�Ӥ+,�,Z�q6�%<�cB�̛��,�:=?��m�Z��\f�@�W�Opɢj`f}(�z~ s`A���С c�������\�x�k��A���/��(8$i���.�g��2��9�ߴ}9S�?�Z��>	?����ݟ�"|������`��0��0��>�!k�QFI�G��l�e-2̞tMI�����*�:=������/������ �w�ݴ�J����/£�?���U�7_.����O���u�{�s#�F���Y��Q8����ZVaE��٦}wnR.��D=�cѼ��֏�ˀd�ς�H��_�Am9hDt?�5(���/O>�(D=i��d����
I�q�� �~��.��Ïٮ��z_��_������D���Qrm=�
�ϸV�^���ԋ�M�����0'�v�t�fQ��p��`���z���2�5!�a8nb>�3��+���Tf�ߓM7�9&�K6���Q��p�?� �D!�[m��,����oў�G��,ҾMH;��z�'����ce�Ek"���L�rprY� ���q�� �&���4�HI���9Mp��| �ð�&%�А�͆b.�q�r��69y���O� M���_�Tp��iWVKyp��3l]���{�`h���ȇq��#.#t5�KF��gdO���(��(`���)[F�/{��3��Q�[J<0o#��͞REC����Q��SN%�k@���G"�l=��]��^���枼���ڙ�@�HJ���ш�T7"D4�%��^�?�S.O)��U��CT����y������-�t��No9�3v�f��+�;�y<�����\�+8���ϻ�3��H��\��EԞ�B��L)M�.%m�R������m���o�o³N��w��Qn1���g'�����ů��S9V�s�g���p\S�Vҿz�2]�#r���%�0��6���<�T��7ὪN�#�FvW@�y�m}�v��g�����N�p�G6m�Ӽ=���Ml%:+:r����'*mX���:��@�7�M1(,�G}#N�`�P�^S$�����3��&�;*�b[X�5��Q���߆&Eo���l�:���a�ҋ�8|�6���$�g��2�&_*�C�d�OҪ]{��*��D2����}	���o6鸱LYn����;�+gF�=�U���CI��B�����7Ԣ��[�J�b��Ԫ�9QQ<�i����Y���6��:=%\-��{�o?{���}���u:J(#:�H��^=�i��/��o�?��_�O<�4��+����N��H�2���8=9�����i�'G����1�o���?~�o�(���}'ԝ�)jIa�s,�Q���>���ۿ ���E�ި#+Ec�	:^KW%� ����<�� ��t%ӢG��]m�f�Qt���I��9�)�F��u>�26�PN��<�|�d9��AJ\V��U`H���['`;�z�x����j���~g)�TzvDG��������9b3Ӵ������o��m=�@��+C�����6�c;T��l�Sھ�+�耝��`�08��L�L��|gue\A�$�%�K� yB*��Mμ��-�b>J�d0�Ϡo[�z@(/_��U�㳶���q��^�za�(e��g��+air9g'Ϣ�^�B�$��W���}��4h��2�G)�E���P��C��5�'Fە�ں�Z
/�I�w��oa	p�`.ZTy�=�q,ͩI�u�m�z:)/���l#F���f,��+�,����!'�V�����(i�$�\�����t �a��6='�F����#\�Ds) �&��N����h'J�,�YzEO����!�� q�
�����x�����H|�hi+[<����=�*�/~����	xû�	�OW1�p8�4��C��4�FƳ�q(.]1�yt2�!jq�����٦����|���u�!�p��M�zhZnR��]�qL��~���Ǡ:���?K�:nT2��Q�d��C
�6bB���lP{(���>2�Wm�������Ⱦ�bz�3�k=�/���$]iȠY"@�WE�n,�x���@�2�:��q��5�*a�@S�q[��|�gS����Qr�,]�lP��T�Őo�2o���MU댽��'{"���)�-la�P��M�/F�E`=ĩ��>�����6�]�'����u���:��~2�����i�^�jq���>,��	Q��Ǳ\�u�`U�d���c�<S�Ï�h�n���V0`D��w� ��(�`$5�X�J�Wz�cS��H��V����v&!�X�h�}_���A��oxv�h�v=�W� ~����n��ۮ�~�g_����=wA{��u�y���6�x�S�c�$gP#��ۤ��g�1��߇g�����k�_�"�=�H`�Y!B���\r�w�����#��V��V��#�I�Q&k�� |,�A	�54��_!E:Lh/�� r��;TĽ��z7�]2nD���y�L�Πd�R�K�,���e��Y�/��¦ �9��,�HEID�B�	�=#~��&i'u$�C�*���[��@-�S�=�]�<D]���w�`��X3%
Ǡ=`"l*��3X�0kMV�z��+�e��X�9�P��Q2Ƞ ��V��C�S�x��CH��EApJ�-l_J�"x��E�����Y9��z�oj��e��t�C��Wt/�� ,���zt�Rs�� G�۬�D����C��V䝞�"Hy�P��F'؇qw$��@�qRW�}70� ����1�4e�=��7)�,�����_�LXV �dq�u��8�z��Ey߳lǌ�����&eȥ�ff��ޒg{��Z�/���e�ha�b��e�(�*֍�I(5Ѩ��҉2dyYK����:g���iR��R_	��������<E�!|��L6�>�� t�U'v�>�I�����ןh�$��pČ7Lp'6>�p�S^�C���;���w�W�컝t�,D���~�`v��bhaV�^��$�'H'ӂA��p�߁�x���_����ɮ�y
wL��$]�~Dy(�@��ܟ���?�1���f;.Sh#��X�we�|�/�]�Q����2GN��D*�g%�i�*A���m4���s���ãa�����i�����z�� o4�l<�9qӀllW��eZ�x*��	�����wQ�r֏Y�SYj�+�nG��sI�\z.�zd�tH���y(E(Fv[8F@:A����_܂�ԏJz�P�c�|f��Ѻ���G[���q��q/Lנ���1�0���1��g�B_N��ḳQ�H���>%���-����#z6���GN�,�Y��\x��r�kD귚WY�Qt���V�����^b�@�'�0���:����o����|�7<u�*�7��(�I�	�s���t��������o�w�x��yܩY�����Bu�K7�j�ō���%�Ьޥ�]�Ë�]�ͫ�/	�����+;�I�=����"��+%������N�_������(Gj]*Ob`� �Y�1Oe�t�6�$���.��T�SA�9��+�����9M���LuL���V/��s!Pl@���RQz������0�W���#FA�Fb��n������'��z~!z��YU��N���øSo�� ݑ��ZF��(��6Z��UxeBU�����D!crCI~Z(`��pލ�A��pa=�������Mѓ�y�B��I_����^Ӈ��-��Y;�Ԣ��Z�b]ŔM�I��8XB�_m�ml�`ؒ���8ԢHW4�_"F:�d���I(H���e9��"u$��D���ϥ�w�=��R%A -��M#؏N�8�Sp��G��"�.���3���cCz`�Lu��}C����ƻ�����v�a�?a`A�ͩR����R�R6^��+���6$�&��Np��4��%�\���2y��Hu(6����j3�=ֳ�~�p_������:y����� �K�@���?=�d$2����(�J�%�~���T�>p�/�ׯ�[&)��Z�ve岃 ��d�
R��_����|��W�7�:X+y]�S��\������o{�������߃?��C���S�s�D4$Κ64c�x�@"e��5G+g{���SO�w��4�������_{�����CB�\�P.���C��,��> յ�t�H��Z˕dv�d�Fb2� ��I8=W�A+�G��+��3Fސ\WR}t
�0��̕��䕎5(%L�I%�E\%Դ�E+-�.��!2稲jX�Z$-y��ϻ^���=�҇87�{A�\��!��ҝ��CZ�����^�Qt�LdZ�72^f�l4˻'�i Q�N����<ΙG�=)��Ry�������(}�S�_d4��
����,�%���-70�(oX^��n���u�b�R;}o�Lv���'��5�VȓG�f�R6�tj��n#Jt-T�9�Mi���D���J>JN�+5�8R�&"n�'��?V�?�)=� �s��b��T4����$'�{��.z��r��T@�&IF�q�.L9�+Y�Q�m#UM��EEmO� �tT�YG�o��O�O~���i�:]v:����)b��5�1��sx�3����w~�m�7������s�Lt���43�CG</���:�V�S�����>\7߇����/�ď����4��}�0����{Qc�<;�~�
w�?מ>��;��ā��FD�
K{��
�Vr������.�#||W����o�h�:9���G+"*M��^B<5#|o�'z�~#:��	:��Ζ�ֺR�C�Wl�� ���\��#�n���_X7�C{"}��tK�<Z�:Qw��ϙWc��4�$�����8=����(75E��g	!r�3Hx��h�"'��w��s�[��ri�.;8
�r�޹��h*��N���EĠ�14y��6���A��ɒ��K<�3_�<�&�L��^ٯ�������&`��s&\R�X�
�.3��\��
c�S�=�)��2b�ɝ�<q��]jJf/����l����f�-���_��C({Y�����V�eW�M��95���r2
=I��a4se��yż���������A��-2�R�}���Nl��[��N�k�B��J�>iͬ2e�[���-���G"M�J����(����bq�P;�Z��|m�᠞�o��pۋ�7�>�����.��*x@�/fm�|ޭ����f�ӏ~~�}��|�I�z�C��8mpA���7��v��p��n�	^�=�?���\f�n�9��;\�h�8̰!�}��-������]���^��N}�9���k� ��b�$��R㒡;ؖ���n}4��S߭��X�H�Q�"=�.7m�3���$+P�|�dY)_;/-cr�:������DCF���)��8l�ڨ��>��Y�5q<�i���ֺ>�����Ua�VD��e��hn���Ӈ7[�����ed��݂���c�+=̀�Z{]Z�AM��G�A�ې�S�òp/�^��ҡ%�Q%���zS�<ے4L�����:�9���"^���ޝ�u���.-���$j�����F�k��W~9o@��z��C�Mrvp��ŝБ�l��O}������_�-YT��y���8o"��]�d=;;���^����[��p�'���#�>��.��Nt����̶��북���̽��oz����n{ɷ�5�Y�>F*`�ˉ���c�:���}	��C�k��M��ʃU�?���N��<1(L쯤k�Â��!i�5��з]�Vu�D���$�E�
Uʲ��S���u�@�8T�
�<�^%���N�Om�n��lE�ED��6Ǐ��A�L�&z�6}h�ީ,�˼Z���`UFG�͝�=�˅�5�ӱCbt�o��
�wr�}�M���a�*���ֵ�#��p�BA�st��*��9��P���8}'�˛��͙��^��ek��k=_F�u�!�P�J�����^���7+�+���١�WԦ�j�ѹ�?B���p%A�|��=.Ԧ�آe�G�7�=���к`xa��N������o<H��-O<�@J�D=�v�E�5~;C�E9e'j���Q>m8�*Bh/�R�y�.��*��U㠮j�5@�S���~����?������1�p%$��v`@��7s���i���^����|���k_��~�N�����ǟ��.����݃���Ͻ�&�����}�M���]מ<��P��6���2�j��M��ǟ�윾FN}a�ۧ�
Rt>N-*�xo$EuHC�1R?���64�QY�2���R�$[���7�<:o䆜q��uS�\izՔ<�ޱ8:�b躤����ƹx�q��d���<�_`}�����*9��i �-��M�������;�R���˜�����<�2 mō�*���$h��PN���`5��j<�y+�����PZ��H"'Y�d�- ��7{3׮�"���XZk)�;���q\�33<h}Jk��y.)�k��T1�at���l�dnʞ�/�N�i�
����[�~��o><疛W��BN)T����1������lx�߹~������_�˻���~|�<|��y���j�����ۃo��i�;���O���|#<���N:	.�;�l�Go
����J�H�/��w����{�_��gΡk��d���	#�F��-����S^6��rf�
[r���Z��N<v�{T�p��&�?�T:\��N��Ӵ)�FJ�
[G�Kdz�C�ؖ���b1 �r�Ibx��ɦ#9���3�sz���dN�[���0�r�Q?��Kș��Y��Ъ�|�c��_�k�Æ�tma��b��X��[.ˋ�'�O�\QS��_���������ɻ\��iY)T��)aT:y��F1l�^�-\ٰ*���o��ԥ�W��(o������K*Ha��7[��ղ�T	����+m�W�p����w��x	=�������1�r�/5/W8���R�3]�)E��&LZa<y�uqër��']DZ��E���|���X 	��������r1�϶���V]�pq���^��[���=\s���cP�k�CC���é����t#<��[�5/}y���y{ �	'�:vO���l;љ��0�d<i��9��o��X���[���|+<ލ�Ύ�zV��^9o��Q� 9���X�6d4%��i�)]ܨ����RXV�N�t�O��I@�j:��<��~ܼ����Y������d�4{�v�.�"�I=��Sn�88#İ�-y�m�+�L�͹^��(�yy�W����*��x��[V���T��|V���J�G){na��*�:V��CӍ�x�V�u+vm4���.�H�d��<�x��Vo_��H��3���-!8�0���C��̦uYgd;�^���ӛ�ճ��5D��0+�@Y�q$��MNq���5*q���h#E�u�^��Q��������sp�^G��Jrs�I����6������j�����M�/���E�������~��.m�`w�$��+8�'YH��!�F�c~�~�w��@�f?�ٻ��wp͹�P�\�QT��X��\n'{����u%�*ʃ�9u^nv��#���0�c=3�)��*<e�J�e{q��t:֡5��2����0/�5qTg��Wslae��%�K$R�~�k�$���s*��~d���x��=��^�����F=�;�]:��� ���a�/�v�7�|���d���+�ܹș�/�w���KC����Ý���t�XR�6Į�����eO�,�ߐ\L9z�6���|���sN% �s) �bѽ��|?lE�"��q�k+�x[�5֌����gI֓|.��Z��<�)&��Ӗ��	:%/m���9_)HbPH��l\���&І�~���F��{6� 7��(�
�]G{w�g��8 >�<B(	�ǅ[J�赌�)�W��uZ9c����ڑ3^:-9vR�b�쓢ZE���GB�=H^��}�c�t��E�0�u�꣩g]�9��8�'����+��?�s{'�RD�x�4�=�� �
F�m\t�p�
�v�B�v/��	�d��a�#��r�غB�چ�&�P(��_�p����o}'���/�5O?�RoJ�(�0g{(=k3y+�F���u���ྵSE%Y"PB�^W2��m�!3��S3�g2���^�-���}��6�N�Hz��@q�B�|y�i��
��\�{��%��	���X3����9��Iq��e���DĂ���\��d��ے�P2ds��B��6Ȳ�����"�u��Ȃ����[R�%�����˞�Bf���:�XvΌ��J��_
�@�m�g��n���>����0H��H�ъ8�r��
Jri��j �5�߆��\vA���#��Z���:+4Z}P��N��p(gz=�)��o��d�(H4j!�p"{�u(���#\���}�
��~(��~ԝ�qj��;��>�A���n�t��p=O������[�kFmSd,�f ����~tb贩��N������tW�u�1T�RH�gL���v��>���Ϻz�f�.h!�����oq\�R��������y�$5v�|ם�����=���C�9:Oa(����cs
i��y@��<"OJ�h�E���|�(VM}_�f���ɱ��-h�}�s��'�qx�3�3şeD��E��:�C�W��@�4Z��)zYI�=4_Io��X���s���hu�E�c��V��K������:�ug����mF:�]�3���ֈ�di�)��j��vx��jmf�UZpY9pXi�]�����]��c��b�r�I����	�⒠Oq_ި�J!Er1
&AY��ˀ��&I�Rs筰���S��R��Hs%L񣪨�Z��lʔ�j���tҝ�li7y�Y�s�
��AO� �r���M
Rś�5�3��gA�_Y��Ag���E�+E
𗌝��(��e2��c/�5�s�N<s)?���nջ!����Ud$����Ě��
��NF��������`��;������?	'B�!�p��1AC&����%��Nl9�|�ܧ��M)���>x,Z1fֹA�Uda�(v���������Np���K�ëx�U:9;ˆe����~����1�U��ҩ5}j'���~l�������](4�u�������SV'.'�B-�����|���d������@������#E.Ʊ���J�KIt>j-�׍�� ��B;���1�#�U
�7XZ�]h3lhКYaD,�-�T��\��&�[̓3瑞��R�I}�0ӭEl�;�	�W�sZ۩|ڒ̶��?䎵�_�Y&�n�6�@��P��2�#�&<�����Eه�S��N�|2�#���W,,ڼ=�HR�n�SW�ܡ�=�myC;�\$ب\f�{�ҽ���@N��%ջ�À���r ������,Z��������3�_�ͻ��[�	��-�&]��|F:O�1[��:un�t�7��oO��'�sJ~&oq �Y�Սv��.<��E�'�����>�n8�냣xt�
ZVU�F�T7�Ebm4���ǅ�����;��X�	�NӴ�M����_�"�k��<�UV1���~�"�q� �,�G��ޕI�Y�.�6��%	�.:R�4�X9W< mz�@��*A�⑓�K3�r�'�b<)��Ȼ	*}�֔SY���A�T!:�˼p��D��U�y���8_m�<��Ɍ�s�gT[�͍�AC`�������܎��ahNiug}����JdU�mf%;M��Q�q����z�xx�g�����@h냖

zЦA�&�e���	 ��{��-p�Ȇ&�t<����i���ae ůW`�M�F$�>xM�� @�n�e�`֤2&C��;<\�p��K�A{�G��fC�X�|�hͷ�<w�it�W��r&�EsO�e`�)�����S���iK8�6�`l���%�,)��.^h� H�<u�;1��wQ��T��a���5�#� ��j��Y��awO�5����]����7_�t����I#�r�ϒ~���U5����pltK������l����1�E~�����p��I���	�u:=F�L��mZ�4@��H�� �ﻦ��;w�L�k��AO��cԎ�x;d�3���-r�0$A��ഉV�6HJcL��X��	`�v9�OcF�M� %��<�ĉq�ż��(r[P6S!2�T\B�{�g �8���N��Qz�����{�{1�p]��А^2�S�,{���[8`��"gdsft�����
����p�J\���/�G��&m$�D�0����7�h�ɑN$�E�ۚڏ�Γ�k�"ɾvM<_T�|�rP�$6{�Q��!�_��܊n�|��P�Sh�AzZ� ;)A���)�z܉����?��߃_�����gN��C�$r��ST�ph�3.�6BN؀��ݪ�9�Y���uv�x���{�㭿��?�?�����뮇�Y�j��5����������6�c��
�W2��1�w���}h:���1E6��ܹ,=j]9}f�>s�闩)g����>[�Q>�����%��!ª4_�勛r���,��O^ߐhJ�ɐ� : q߰s��hL�)B�
�G�Y����/r��&VN c�XR96g5�n9�T99�!_U�n����W����lj#�D�n>�<8�۴c���K��tB�{��c�~��:q`{xr3p�����:8���~�YT�q�8R:\�(���
�%,��d �tj��ҡ�}4�<�M��ō&Wxq���1VЧΒu�i�1p�������C2(����=oȯ&�-α(׺���	�+s�C�')K��fL�j�+�b3�(���8F�q1��L��КRVe!e�X�.i_�GZl�P/Yy��Qb�d��N�]4�S��כS�˿�p��s���|��4ԅt�*���P�\S�h{��ـL��V�X����u'n�f������~�t�<�<'�f�A��7�����A���h�Nm}������ 7��k`�baN-Y��.�w�"��� ��"�㛩y8�=��=��![1�I�J�e�M�A�p_cc�`|U�T+,�.��Q���#��T������b�܈�7Nll�6�%�dy^?�}9t���}��h�s`���V�uu�e2+ah��u�m9?���U�8h�X�*s���'�*5���O�?����̣��S}����7��_���C�sI.c�Js(E;T;Їɨ<z׶�.���K�?L'^!�q�:��c�ֵ�%�������u��!�ެ����Zxߗ���W���_�����.C��$80�u/p:�gPU��ȡ�"ڦ�.���TT=�x�4�W]�����?8{N�հ����"px��5l���1R�B2C�� �<r:wb4�9^�T�O��_�<؇S~��oT�L��������D.��[�tgS������|JW�4By�B����la�`)MEn���|��AC>��������A��Q��4g�z $(%�I6)�â~ԦJ�=�m_�(5Ðs�౜^���Y��}�UʙZ�"Т���$��3��׫��|j����3�#���Ժe4����ey���̍G/�U�FU���:��0J��8\���E��1�"y��z_	��*D Fl;�\�B��ݐ)��#֕4�i�yqNQ"u�K�8sO(n~/��>N��.[��a%Z�S����똧���9bF7Z2��s�Pe��<	Z���FKk4��K9��x�h'�w�0�V�X8�s�PM�2&�u;m$V�ϖ�i����[��켘���a(͕rt���M�I�Ni��5��f�@˂�g�P��¹�NLU�FCFu0����}����{+�g��ë_�8b����*�F �h�KA�3��e
��FL.��Y8>��{�����=�ݽN6�������O��A�¥:���8躸�*n�:��9<z���ᅯ��
&7\��➯�~�D��k>3f(�->K9��Z�,N��V���S/V���j����J�^����_:"D�����ޜ����c�P���g<݉?x�A;��)M���*�RԬ�!���LH��bޢ��]���Qc��kd6M�[�f����Lf�PuD����+�W��<Yyp6���.kmu�8�-�IR&]�K�S�$��+�@GJ�2�"�5\Yph�$xyIA;��X�,b
����
��w��'�i!�%ދ�njnsO���d��_etl��;�V'l�������t����s�����~^�c�����p�S���+� x��b��Q�/���(��z,�Gd�����jZ����~��	vv���tS+�� �;�q�ߔz�c�>���0�Cpו�ɯ��?�|Ӎ'�ܑ�x���s����n�t��4��(P:O�%w���m~y����3cI�1痪%D�,^��j� N,[(B�`���ֳ?H!8]<:	W�דL�;�;�KX���
v�y�}�ǡ�"�T^�,L�:��j*�"Uї�؉��ea�n�.��wYC�	���hqY�גea���-{�.m���ԃb�"U���l��}�]��v�#�I�����c�Xkk�M�ڼ-��`o����Yށ�7�#�?v\��nS�Hy����D�Y��U��=�9���+�9C�b4Q/�M>IX'���5\_���5M�h�2���x1�ak���@o@��*�������'0{��U�,�9�=[&	[�� ���E�A��3T��Pzy�aF�X�΅�̜>������M�+�0_�
���������.s�(���y�{u#�b��҃�E
#�l����>C9�,�cB���d���t�)x&o������]��5����G��}�~N���I��g�"�^��cVLe��:,>���߃}_UY(L�_G�0��Sz2|ϫ��u�;+��\�7d�ӏ}�
�LRD�]�M�v:Z��x;�^�b���=v���C��=_���G^O?u\�I���Tqe�7xYސ�jr�`^2���gt9�xϧ� ��-o�O>�04'�`w��9��J��Һ�e�D��
�:��	Zq�{p�:������}��O������E0�Y����.��?�h����mP=��Fb�YB��Bb7�m���1�Oxlـ�pj�o�RYy.��+�4�SsC͝V�pZ��>��T���@�^_��kĲ�r�Kz��9���֍��2@c%
BD�3����S��/T���*x�tjOr�ġ���*�s3�fE���+U�I;dd�PƂZ��*�Ck�P.��wM#�ҩ3�F�c�^6u�p��Jh�ˋu}�asǻXYV�/Xn�����2�ʧ5�6bh���"Pm�Nr�cHlG�kF�kj���;�Pul_�֚�J�{���@�ˣL;~Z1�+���E���
JN�|��m�< _?����$�1$���ҸAfZ�!X��g#�w!�8L�W��� ���g�fā�fH��+w�3@hcH��rI�J�>l�7�tr�l���A��	��O>߃��?�#�[_{A��s��P�$����W�<��4���I=��m�Af�0vw��'/����w�1<:ۅ�Nu��N�6d�Ǒ3�ظ߲�脭 �Va�;u�<y ��O����30�C���.�D���DL���_�O�}/�8q2�^�䐌s�H��R��L��
��S��eFhI�Da=�&�!�t�c��m���Ha����J���8H��۝JW_Y̮t���O-�G�Q���oaJ^"�ڂ ����-[�4w�3����-�`*�]s�iQ����f��'������:U���E4�(�2�%����O��{l]�Zf٥��Ի�&iqY�D�����uM+��u�2[�$������%ٳf\D�q����""%�̙�9�YEr�io�#6i�z����d�l3 :@�����W���)+��n���Rn��X�"R~���Cq+�%婯 �`���!� ����)8Z��)ߜ�U�W:i7ԾU�Lc��P�x��]Y�O���[8ް��o�qմ06_JFKK�<�qt=�]q�0�3��(3gazQ�Q)�4�9kP�>�Y^���"�0���2�Qף���ј4F���CI1Lez�.l��]�,^,Un��]�!�X�u��j5<�87`���6e,I1�o���-(�I����ٰȏSa��TOU2�ū������~�w�>�����'�����o��oNA��>6Z}���j.�>/��2F��U�
�#K~����S�������>�?q�S'aVw�gUt<��*�:��2|�׌#�U�r?	���K�)���!xǇ??��W�lo'%$��^W0w}�#��u��c�����A��D�e<ɦ��t�&�.|�~��I9�=���g�r��d4gQ�sNo����2��a������˹1?��h�d�	cR�¼�8ta�B�%N-_�M �DV/����Go��l�$��p�S��1��a�4u�f@V���K�:��m��/��喇��� ]ZAsCC��4��W1MU���P;�
�^D���cdY���8I��Cɐ
k��f U,���*=��o�RB������0�4�Z#6;�~'��S� �uSp��L����B�����(z�Ʀ'�=_+�k��ƻ�X�������������Rtc����v���O<w���s/y���~�?{\P��S*1�`�+I��F����W�;9�_t:p�N
v������/}	~�_�|����ε�vzF�N�7<^ψ���]Ž�����R;�>�FP� ������>���y��DT��<��E��w����sǒ�+�!`=E+�2��'*Jd>�%8/�l$gS�06=yK�{�����k�m��g,�;h�LwX7vU�=��V����W�=N�����k�8v��:�R)粙��\~^�"���Q����-�cV)ǉ�F���B�P�|��}�a<��A$��r	;��r�~grH>n��'���\Ӂ�� �����<
�	4�B�*cq���wQ�������q�eۼ��JjI�x��?[��`zX��l�$�́_<�bzܠ哕ήΆ��/�P)ZfiΌ�F��2K%�?����JssG�! �>�L<���K�
L�09�؉�u�=�܍��=�1�����D_ڰI�<��5��'���(�O!��*�w������<��L���|�D(_p^Ո=Dy��+�jHf�6�*	���v������=��|#���~���nzڍ ���`5J�&y��1�h「�x�5��ʠc�Np���¼�?x�����n�ԃ�����y]cU.�I�z�hx3LC�he�������f��f�Bsj~�c�����k��P�8����z�"��#o������\E�U�9�F�ǄG���>��rc���%�w��&����a��2���[G���q��ٜt�$�>q�Ҧ�X5�5���ʢ��YZ跁~kG̒S�T�]�ợmpVU^���/�{��Ӻ�H�9�n����.�9��#�M��"y]=�a���'̑6;��Y����z#n�I 7o�K(b���U kM�>S[��CY��B	V�"#�<(�����f��d��u��J����^�9��Yܩ��.2�S�稌��ؓ��C	U��uԙ��,�%���>q�i��N�����(|䞿�����W}��a�{�J^�R�M���7#:w`�9�8C�r�:]W2�'�K�=o|�[���<ԕ5��zp�22ú��W��F�U�go@}2F	j�*�#����H3�qg�k�>�_����c��������<<����+�?{/|����Ω�4@қ*���azaBPX�؂�T�\�S��ӫ����,Id�lrM:�s�Ξv[.�����sY��.[�S�/�E�!�5Qp��^�z��[�,��sJ�-\I�&=����فyS�7��7kh������ry9p����88�7�I)P�q�璥L|�R<�$oZ�����w)B�h�~�M�y�=��n��N�M+wZ�[A��UOLM9�
-,���E6_Z��VZ.wʦG�B��-m��C�[��t:*�9ڛ��hr��  ��-�������D��Wg7�&b���9k���0+�&Е�@Nk8��튆,�"�I֨df V.Y��;j��XPmtd�HeUd��C�
�vs�a~j�:h�����;���|�/��N�%ce�á��z�T��GC���e^���;qr��>����|���G�I8?��:s�	�-#�5��F:(&W�6�Uc��3{�.nP�T��e���/������p��/���o�g�9��|��_��}��Ỿ
wv����D[���)5�q��P��4�~��C�nyC\�T2�w`G�i���p�)��9ѽq��kd�f�j]
]=�4w2�� �&�6����TѾJ�>mJ���fq43���y�.��K�WS�_�l��n8�Pou��&E�9$Z�Rn�����1�~��WT��x���U�k=�Z�!n.;T�"TE�\�z�+A�����%�W�Jr� R�����TEd}�d }��l�%G-�"v�OU�H��Ju�G�9�n��z+�C�4��4�)9��uO�ņ��B���N�8�t��k���>�$|����3w������y�x�ͪ������,$�z`���a	�j�uw':O<��y��O~���?��<����P�)|xU�C5�ǣ�g�$��0F��L�����t|uR��S���v���W�m�^�
���	g�v����?������4���>�{��Kr� ���Z3P��Vϵ��_���I]Xn�S��_����S������Xl�J�%�,خg[����a�w[c�mY����
t��U`y�
.d�ȅi�I�B˒��F�+�M�JEq*�x�'Lz�`z6�������w|X*�q����y���p��R����5�?{o�-�q݉�Ȭz�tcGc!��N AR�H�"%�̱}<���
� ��g��}|��c��#��#�ƚ�8�(���Hl�@�X[���*3���%"#�2��ޫz�WU��Ǎ�{q�Fj�����c�{R��6��~�d�xv�i\w���i&�Ap�6ꊘ�c�R���kG'tV*�p���o�M����.+����(x���o$
�����B������}7����Mq�6"����E8&����&u�h�֚�@A�Ma\�Y	�ClVpX̡8~�������;���������/�g�(�}�6��r����V������1\��B�6�>��������<��������s�a�Ի��Z��s������9[��+b�-�ʦ]	55���[���R�^������?}�'pn^§W��+�B5�8s�)c��ao��|Ժ�6IZ��πȟT��O}��AN���+�gz*�B(Q��R����F�3�q˛*��
��pހɏ��������ʽd'ü��Ml�7+�j�q��r�c���t���J�u�~���r	��ғ���Hk���Lm��Cz�b<���`�M�8�����w�K��Ь[��c�4�� �"��V�e�v����`)����«7�Fm@�*�1�����XOgѮ%6*���;,�'(.�����c 0�iD`��_��K�g�5T�̯N��O���x�����{���'��n<���¢�|o��]�F�hT��t��q��S��F_���*���{��o�_����W/�
�O5���gah�4�/�%G�����SBo�^e�(�'|�i�����Iߔ��5������������o��S���?�.7խ�=���#�!���\��,9Av����C�(��H����7{t���s���5���o���Lmr�!�V�Y�X(.�)S�L��R�43%�3[
��[;AJ�nZ�ǒ��bE`I�A����j���<���G7tb��;�*	��[^�h�Ҙ��vŚ+
���3�G"<sb\�I˛!y����6���QO}`�<����-�2m�Vu�;5ߎ�׵��&ipm��S�4p.A�����=q9�_]�R��C��1��|���p!j���v�4a
���6��WtE�"��ZA�1�p�B��H}���ɺ������70�8td��
:cHAϴr\͜��]�P
Iઔ��"�ԟ��ࡻZ%@��{�ɒ4��`��57�t�����W5�����=��^��o�
��go�٢�{o8��q+|��������_g�J8e�i('�8P�5T�<;<\�����2���o��5���_»~�VW�JU7y�>w���4�I4��R���1����n�A
�mH�۠Vn�eݟJ+��bS���UPg ~Ӽ�\�b�>}
�zF�,m��ښ$�pB�#X����ʣJ���$���)����8���G/B��j�K���?��#�\�a�V�C鸌���F7�v����h]J�伀h<u������7���P,�I��P�4 y5�60.r��J�X
���a�A*�)�j]�y}z�ii˔i<�y�Mc��;R��KS`#}e�<��0]���Ρr�a
�l	�2$�:xKQr���Y���1:z��*�[>�A3?�LL��T����=���o8���5%�qP�}�<`Q4{�1H#�"J��f�h|�C�GS�(����ZB^Q��U;O����y�2�^���z�2����?��p�=�x����w��}��v����o��oUƃa]WVF3�q�$�ɕ+��Ǘᗿ�^�����o�˿z>]\�O�5��)8��Md��eqSFk���m%��un/�{������xC��c�F*�a�B7�.*����S��F�i�>3��UjN��X���c��
�}#vH���/4��$?���?����]0����T3��(���2�@��f�k��,�"^,1��+ﲌ���c!!%�k�"_�\����w�J
#��L�2e�8��f(�VSR.ϰ8����j���:�o`k�3��*F�l�츪�9ڀC���;%�AP`ڬ')
��]�5fu��@p[s�w
 :��U��1��怏��q��̴9Z�o��'��bH��-��IJm��˟*�J���P��k��C�7��8ѥy%��P�$��i�����!��6T�iˍ� �����	��{���:�[2$[����X��pa�-C� Gd�h�<��N}y���\���E�+��p����>h��.
?~�g�/_�9\�p������o�.4�O@����a�����������[~�T�i��qc�zϜ>��'��rS��׋�Nq^7��1���I��"�GVr�yC���7em=����3[\� P�*r���M��z�OD	��ZF_=���p��O4�{5�7��-�喖F��6�j���m�k�G���RΛ(Ӡ�*F�V]�Y����6S�M�>A�lj��8:�V���1��ݷ*i���aEZ��Y���	�����Իp%�fV`�+/�k�Ǻ��
�߁�����{ڠ�D����H��B�N��k�����Uf&�r����\<cQ;��Ee<6�������94zʯ���x���7o�����[��⭷��w]��}��g�բ�O��;~ ?��{~��e��$zyp�	3kt��x/41Jp�;|]�F��z�Jn��Y������#[����!2��G���5�>P� �����=E�:"���±1�h��p��ATJ�kȴt��f|h1NgI$6�����ع9�
1��.�'D���y:��3eʔ���~���}M�� d'��IS�52��c4��VpL�G�w�w,��=-落�� ���(
���g�q����i��K�u��yf vH�(k*�}l��2����C+�k.z7d�[!�x�����|{U���Fc� �а��� ���4ⶑtAڪWk��H�������yw{���Y���g-D��:�w��*X��ӑ��p|FI��x'���Xo�a?} �7���g��'X�L�����������Ǘ��`qEU[0�4n-T	U�Q�KX�JP��� �L��
{����)<]����mNg��_}͹���^�7������E�$�����lb�>g����1��)��c̗#^_����q�Id�E�.�?��+�**֦7�4�^5�Qy���:�r'[����j�gA�,�R�$l2�D���1;�Y��[���͒��ޓ��#ښg�B�}(k�yq$�}Y���ۣ�l�^�	��]À$ MMn���NEb>%�Z$xa�B�Wz�)f�����9���:�xd�^cY$`���x"c��)��*3�������S�Ie�����z��)gP�+g�`�Vhv��\1j�Wͳ7��5���U-����w�qH�t����у�W�Y��&K��Pۖ@�W,L>�H��@}Ҩ��^�0}u��X�w�k-�8�%�;�o��,��1�M�ZT�o�R�r�4
j��P���8m�l)uyye��Ñ)���!��Ry\��C9�ъsT�'��L�2e���-=$>���T!��~B�mրc	hx����"�k��<��~K�JTD���r^[Y	����:*C����0��0�mCG�I
�ytP����ДL�C~x�<�vI��M��T�c�BW�qY�6ז�-�="���j֚�Q<)�W\��@W+��|�*�&o����E3���Y7,;L��]z�ҋ��:�]��\��ҵ��U���G9'梀�o{����n���R�:���2���B�U���J�FQ�s�¹���j��k�r(��t(fP׮<�m̀�O��v"�1NQU�.8@�jz'Ac,;��#�q#;D�#}m�}xc��B9���͵���8�S�VX^���w�G����74����NN2>��&�2��y�yDq��p�:'��t?����,k��w�<|P?$�Z��y_�*�ƾ�A�}(S�y��J.��U���h�F���aV��U#S���=Tl���]_�Fַà����I/3�"�Q��h8*�6�e2��O������2�
���M�Rā`���Fh#�Ao;��/�V�,eU-dJ�T1_h�u��>��9:�1/ETT���5^��0T��]a�B���a��T��7����W>Z-�]�?�Y�vmZy�vm=v����rބ)���C��7v0�V��oui�RWV�*�E��ҵ�ӯ���"��WB:����R�Ɔ4��*�5�;�gJ,�=hp�� U�|�"_+�N1,)ۀ���Ѡ^��A������|���d�,��J�'Y�$�����Q�]4�Z;b}ikD#J�҉�,S�L�2%iu�Zβ�����4d?�4Ҁû���)�-�h"�C��W�R��c-�A]/�5�Ϊyn}���0�7�}�Nt�(�N���� ��ڃ���t�I�؅|*Lo>Q:��p�~���men �r�X���',Ӡt�L��6��]���q�\���.'���m��F8�I��R�E]sV0��]�B��oXoc]��"�`v5j�Q�)� z0N]Sl�\ƣk�B��TM_�ex3���)���v�,�e��J:�8�EG/QA���$�d,j+�&��q����[����QA�6��*��ℨ����d���R�[K�g�
X�1R��+�{{��p�1x0wJ`=X�/�5��v�!7�r��lx�GIY8��v�e'9����`.��*�!pm{T��%\;C��|�Ȅ۪����x�����[#$�~k@wqT́�r��ZA_�'�ǈ�W��e�֦i��-����+'$1xܺ	�n�^ax�E���d�H��_*ÿ͐=l�_��n���A�_��~�x�Y�$���Q�(���쨡ͳ>^����o;e�D\�>����4^o+gFcS�%�dʴyҰ�ݦH�H��[�8[����%c��^BJH-�J���8mB�=�[8(�N��u�$dڄ�x����pvg�Z�:��� �����q�S݆��6o�qۖ�]�v�Q]��0� !����� �!����C~&ˎr9�<�1^���(�a�K�0*�BR�=K���V�˗h�@��?���?�v�z)w%��Q�G�$�
o��̕'�'K3T��c׭���(M
u�ϔ�[�?�vї��\`���	���qXI�;t�'�}�|���'zcs
�4A}ҪI\.�d0���6ԋ�ʋ0�
�@a�*l��NNS����B��]a�Ϻ�LV����p �x�ڋ������t���6�S��0�!��O�(5�/�t2eʔ�xh�tjy8��������t(��`Z%�!�����e���^��6�#i�zL�"Il%R��4or�$�_��v�R��a���+��7����(������Y&�.�~�8N��ݣ�K�-P� ��)��Q<��x��,�^zʞ 5��L�$�J�R�|��g|�O���2Zq��6 qc��jd8�c��1:k�+$ˮ`\�G����� H�gė���iq����5�E�K 
���U����a�g��z�'��u'I����G���O��h���aޕ��� e�$1�!������*:=��ASm �j��(ld�&Oԉ!���Z$A�;��,�D j���;xS�fw��D�8���$�Nj��^nB�<�˰uD�qꑟqZZ�+��Wa㍽�r��mH�ƭDc6J[)&�N�B�E`z���2ߌݜ\>��t�4��@���Z�'�$B�p^���X��Y0%ͤ�GŤy)^�X�R]�Zg��BB�z�(��\;�/;��x#r� � n�tB��+�H�2C�>��DVZ��Kɶ6��j� t[�QJ2D���2�.;�Q��&�,v۲�Ag��(Q��a�g!���jF���c}�ע�\N	�L%޸�� ѐ�'�j�;|�J ���̵	1W�A��ZC�nwt�>�}̑	���d7H;Vբxc(��˲�J���rR�[M��g~[��4�^M���sA�$�W��2�!�[�m9�7���}W���؍Ȕ�d���'$�e.4�P�R-������5c�d��צ��M���f8�W�#/d�>5(dψZs��=V�U�@:���	Z�xc�ɳ,(dj���2gL�v)$fAU�{��
LB�[�c�|�+a��)4�����un���x"I�B��_0�0^(B��Dw��1�çT ��gOy�HĒ62��x?�;���Ӛ�Ԓ��,�yګ�uwi�\7\��C;(E!�����]xQ	�Ksk��;��w�tdJq�h�>��9����;Q�"tG){�����\B�h�9C��6S�/%�x�uЖ�8kN�Rś��=2��ol�8h�Y<b[ч�+z�*=Z�F�&�	�Ϳ]p�*�<�XF�|mO�
ӯ��ʙK�\Ӳk����J��cC0�T��������(ې����[�'>��t�hV�mI)��ѭУ��A]ٶ�[�b�H��-������o!� ���vƤN�,.4�Р�C��8�Y��	���(�P
�����tq��C{�Y.1������o���P2�E6\��qT�=�)4���}�d�a�0+,�7BA��_��	i&J��=�i����%�"q�u�:��@
�
<'aokn�8?~��h�8s9�5S\�U�̴���	��'5$���^�d��6�͙2eʴ-s�IK�hb��L:��`ڰ��
=n'I�,��a�|�R.�Q��x�>�L�$!�8@K�D"˴c��A�Ċ���1ch$�B�\[q:?����و!��Qk*�r:�6Yg&�[�;�x#�T��$Al(���'+��/�dD�N���ݛ���d��$�Gx$�T$�` ���v %ǧ/���/<�[RҌ"&+��c#(W����8�8J!t+\��L�[0�]>u��
��>��Z �>�:�c�x�[~�4�L��Km�H�����LlԑOr
Q��
P8~������E�Z�NT��9O)?��?c�Oci�����`��xa�rf0ɍ�O9J�L����J��0��/����o��$V�Y��J���б�Ƃ��n��1!�v��<�˄��X�A�����?;D��t�_�����#}Ƹ������<�E��$�aJD	Y��k/ZFF��v�,js��(3�=I�D�QU�C���5�&�(�v���|4�d�"��&0���6�A���T ҝ��B�'}��.�m��C��I}#T�Dp3G��x.:k��@�h�n��g+�b�L3���Ioy�WN�<o#-[���>5j�xʔ�ڦ��������?CC`�	Z�kȚ;�J��P,��Y�X��p}�ҵ�_���Q¬Դ�ϕ@OXM�9:�bmi[dZ���d'��GUid���6�I=e�N���T�����~5���R�vd�;	
S��C����/�{E|8#��A ����6%�OX�n�3�X^���K��  ��IDAT�'�U Q������d�|�w���q»�1�o����Ō)�O^a��� [�"nB��v�;�t ��]s��� ���UKT[ ՘SM^=�
�����֕@+���(k���U��R}9fd��;=%̵[��2N�]��wŜ���6i�����f��<�q���r�ؙ
���V1��n�9l���ʙꨛ;S��4/N0�%˸,]%&H�8Ҩ̽w�f����a�q�Y�5��q�&M�Ή� e8��@��5)�襼��5vo�����Q!�y�ֺK�䛏��@�WA)�bY[�<��2�$S��dt�j�.�'�ՂQ9�f,�{uq�c{a��%�CI�J�IqΡ���e�lTӮyP"��)��ն������ؤ!��Z�I��m(*"%��6�ZR����nŐx�Nd���vo6;a�Y;��wzW�)��N��䆎�)]025�/��*�<2e�4--�)cq��?�6;K�UA#8����6��S�$�i��L:�4feO2����x�e���f�rӈ\&/ ]��{�{���(�K�oۭC3eʴ%dOŴ�G�0��|?���m�|+�SLc��"��vS#���4TU{̓�,�5���6�%�!��w��������+���Q��^H!���:H�����;nwe)����Z:0, ,� ��d�*�WQ(l�8(�|K�OT4��ķ4�p�0OQ!S�;B��h����g�RQ�*Z�+a�[@�s��NF�m�B�_�zNq�\��T�$A��ɟ8�C�0޷o!�7�7�֩��c952�i��(��[j���5��mҺ*R|RY��M8������\J����;��w}=����Zƞ7(�x���v,ˍ��<��+��FJ)�Y_���L�M�Y����ޕV�]�ܰEP��y-̔)S7�Th66k��p9�5d�y��Iv��H��\�*+�1�����ϡ~]k�_4��bsVu5Vz*H��^��(��oJ\K��|���v�kԤW�t,fd\���hp�C�W*X#�8�c}�R�L�D�4Rs�2��*	^�Ӄ\Y�v��7Z�a������Xc�_&�>z̞۝(u��h��#�_#�B��e��逡r�Q��Q��o;$��X���O�\"/�S��ȨIwBX	��9�쀰�P��=!����>1�NSV�^0"�ť��V��S��|����-�N���$SFsy��ub`��O��LR!�kZu���w�0�#��]��~o���U�n���Ҙ*�L�2�B�S,J�*z׍�/ҵY�+/�(�~Y0�G�SJ(�f�cV��9?ٽ��h�n�͸�/	�<D_֥�I�M7Ol1�j�n��-��߈���9q�)S�ݢ�M�X1��a+ ^�pM�11��p^��u�Z:`7��U�PQۜ|
K~�"�ô�p��RM�����{蓬i��"͟�"��2�a G�x���Rd�i�2'`L��(�4�DN:�eH���r�(E�)���� ��fj�����?ۀj$�j��m
�ԏ�0����W���)�H֕˶p�=����9Hɀ$AG��`j^@Y[�e��Y��5�MI��y��%� ��=�o&�.k=�� ��N|��ꈩ��
I�'։�ɭ�;�T^X��Q��Z�)�nP8VA��r���d��nٙ�z糎�W���ޘ^�!vo�XM<��i�$���fπ���7B�'��q ����Q���S�;�о�P_�e��:���}�)
+k�\�2��)�'��2 ��r0*~#A���t$F1�>�F�/PX�'��6��3�z�O�/Ɔ���>��i�ZjG�'��J�,B�Ż����=y��d[�e�6�p���ZC�O��O��'�s����#c�V�J�����"͜�\�#P�h���N�SD4Ti�y��8N���^S�m:��[�3eʴYB�p�� ���\��L[��:�ּBe���eP)�
�*i�5e@���J��=��)S�O}c]*M��MRw�㖺�)Z���������	2)��
A���[�0�2�>=��Z��FȔ�6y\�pf��ahP��O���i�C�&6[��(i��$ۧ'O��M�­bb�hr�{�=���5 �=�P����-k�������,��j?�p�}�J�����	� tZ"*N�w=:�iqCD����c/\J>���ዻ�!s�I����#�F�����x+䳪G*����eʴ���N�׾�`�[��5�`����u�2��
mw�%��m>��(M�0$�PIO���p���-��ۍX��*U4D���|��d����X*�n.���@A �
�L(�w$���M}&E���Qpў���w�*��(2�S�Al6��01�DC��C�;�2(�j���Mt�����(����]i��� ࡁ��<*���**�Es������|2l��$(��'56б�E�	#�B��Բ���݀ul7W�L�2m+��rm�<�>&�E
7���e��	�dR���kR�қ�H���P)�g@I���f�:�x�jW:��ړ�vO�2eC�F%�s���Ǹ��d��i�φ��@]�ݸ�������9-���k��n��_|��m�������l����w��R| |����1�G��EJ�Hb�� m=���>i8�r�!�� a�8\2[%+��]��.i1b��"y���1rS���q^@m�����߬��PÏ!���T`n�s��k��=�{�e'*���cJ�Z��E_1�L�gI�<���K����ޭ�;҉_+� �N��l��|����[�b3���<����iZ鼉7��]P�R}e�ү����W�K[��`��3e�4�wH~f/uR��iß��;|�h̓
@�ھ)�
w�H��=�TZ�Q��>�C��'�Ln��].ej\m�!�i#<�8-�e�Ճ��Z3}��q����1Zr� ��*s�%ʞ�1N@3��K>�6�t@�>��0�>�SSU��ot�>����;���E	��8�6�&l�\��>F�V^��&4,�pT�Š��HR���Ͳ<#-q���W�餗��sʠ���0��^J�OW��Њ���D�L�2e:2�mǔ����X�ц�A��h��BS��t�$]X�PH��Z]�]���Қ^(��x@�IX(b�xD+��u-��X���Pe�u�w��`#��2H�)�ɡ��as-�.Y�]b�&؏p36����_f��5�s��\f6|�ɓV��Qʙ8��]S�5˚����-�A���76a��"_˜!<�HB�mٝ{�'2��n��؈-$l����/���ZDn>(Wy\&���O@>���=�>���{#\�8#����h8m�˚�sq�O�yH��qu3����l�����������1WY���t�wj���ٙ�n�E#-μ��� ��T��"r(57^�'"�8T�S)�y��%�0��U��Ρ�����p��^h~�7g�߬T�0��0S�Ocd����3�f�2��DQx��"�v0@+}]4����DOF��)�
-�K.��H���o�2/�������gʔ�x��:�-b}��t�^'�~��^�P�n�>6�BCJ�E4홹����?e���5�̗���VP�L=)Xx0�,M��kǎv��K&��^��ţ�ŧ�-�q*��jI#����A|����G��c�l���7e�����T���>6t�.�=���b��@\�J ����*��K��:�Q$��W�Ӑ�-\�1-��h7�k߆ZW6�y�և��ڤ׼+M_6:�*j��8h��}W>�t��|�k#�����m��$Tr�:�^Q���� ����]Be�vJJp���nꯠ)�]�5t��.�ԣ������*{����S�Oƅ�����aI��yB����oM��j���2e�~ڍq�V@��; �&���I(��:ƛش��Cv�-��8Xr�y�������;ߠ����R�@��LPXWh�����aJ�(��6���&j�c�e�p��A˷&��w�������/��~,Sq�n9W����k;���So�=��#䡐d�������B�=�zOr�f�U%�W p.�4Fq�x 2�����&7�J��'�
�� �5���@g�� XX����|��[T�'��w��������{S��1X���ZX���D��\]�
���;Ν��>�|��G��sgaV(�|x Ͻ��������� �N[������9���):���Q끐��T��<�T|�u.���4�;��2>�(Ղ�\p�.��D�<, ]���L�x~!����$]��S�@��g\�x�"A�����2�9�M��產񝢮�H��jޤA�R��Ia�]�XV��0� of�!�Z����u���U�3J�F�"�`��w
�I�4�O�]����#ŏ�f�7�S���ȒP�+I��/�c�&���դ2D��B�_�7�6w�3�%Ф�b}<��^ƥ"i�1]6�}Ra0�PV�+IH__�����+�G�!��q*Ѱ`��W(�k�!/��}-��^0��:�:h�}��
�/�n��F�U�hVW5�/Kx�����z���.8wjn��ч�7Ͽ���}���3���*Icܥ��|�4իC
�u�<$�A��?Ѱa�)	��(C"�A#�,�[����{R_ʴ*��I<�5�Tw����
�iF�T�y#��;� {�0������#@�k�3eʔ����O|�LQ����\WC!PyY�z`&{�`�u8��nOK�_���Zo����q�,v�p)^3����?���{dS���x&S�u�AܓP�L�ih?O�� ��_�]��b��΃js�P��A��٫�T��
#��F��1!�	h<H����c;�+`2Q���������SR�����1��E�0�_t�x��ocY�4��[/@ ҀF`Z�).��a�j���΍0{*��ڟ8��CY��GQ�������p]���[�=�����V�+KP�ϰI��>�����������������6� :(ۙ J�hoWiW�oh���Ǝ�*l�."C��M�0�e�rc��x���R��dϡDFՑ���<cH�@G!�?aN�C2��J������=�=��Z%�<NA�K示g�x^��V�h�i*��o(�5�o��>��%��F�7�5]�&�������M(=W~ӕ7�S2��s���j]�7��D�7�w�b/�G�:���-��°�Oi�A<�>���2V6��|7a��-$R�ݭ"\;�́e�����y�^�r��2����
�߄�/ˡl]k��Ή�.-+�U
�����->��f��sw������מ�,�t����^&�����)��/>���+x�������R�~�$�%ZB��	[)�ۂ�����
c�xb�#Em�{Cz�M�&%���M���N�Zz�yKS�"j��L�2�]��x�ԫ� �ԭ��^X�\ۀõ�.���$�^��0��wG����u��]�m��ڐi�i��tJ�~hۜ� ,q�$��&�2-W2��d�M������`­����̴E���"O�i�bWhݵ|�,f�Sz��'�0B��
#z�P���qA����tcى�e�'Wő ����,��F�d�REV�@��w��z��lX`�V�����;���\�R5a��P�&�!ͼ| ��s�����}>���p�m���SgAÇ�9�ү��`��p�w��?�K�|��W��l���L�
�NU'��#,�y�i5�D��y���P�3bxM$OO�X6h�Z��WV�y�8�'����G"Lj�&��8���I��:��b�ȥ��D����ʕ���*��ϩi���ey8�fi(o�X��d�1��+�ʎ�v=m�
�6Ş��֬���q\���|8<tDy�8�t�F���������(�©6BV
y�n�Rɻel����A0=6j�1��Wa��,�O�l\�QFq��.%��N�|�ҋ}��yZ�2�
�Ti ?5
H�w<YO��C�iy{�������{4���ˀ�qX��j�x~���y�!��wí�����T�,5��A��ֵ˸�yN7��7����ß�����]�.}�z0&�#}-l%5U�t	O�2��TN�!�
ì(��X��"v��\w��Q�#�"������{�6�)L�L�0��;RW�C�dʔ)�fֿ�붓d��a]�N��6��A�wԳT�n��2��	iJ�m#��L�[��E�3N;��ɦ�eO��5��/�c�)YWV,3m5��a��?VL�'���h����D|� 8ɬ�� ��&Q�A�()���x�'G����`����&�՗���v�����6���<�&�E�P%��4���=Dz/@�d�l ^�	��Ȓjp;F��O���������n�z�2|S��ax.lK�Qk:�pxc�t�#�qgj�!J�*Wa��%����Sw�����~��3�O3W��Ih��V��Nҷ��D��rX�m{3�o��-x�o�k�+����_
��)��F֒N3J�2���D~#�ao�2ȷ�F�R�ph��롣�C(�l��d�u�˕��t��)Ov�E��_W8�B=%��{7��G̓S���Cf�!�V_:C嚩��]��2m������L�Z[����Fæ&ꎒ�׻��Fb̔Df!e��+�,��'Yfz�嵛��l�c*M�J��2�>'�}��y}��.�e�kQd>�^���|�����َ`��K)c(��)>�Y��P�A��5>�Z�u3-ҵӏW#�a��n�|���� �nt��jՕKp�r�o=�0���~��n���(�]p�5�W��3�vAZ�� *��c��O<���~�^w�����
��N2�lY�:�)���m쒚���:: ��~���ݴ.�&���J�?-=,ӄ�:~��^7��+�
ƱR󑔗��2�֚> L�L�2!��Skako{�Z�7��*��(O�(7��mJ� hs���Z����*��u���p�v�E�����!fH�+��j3=����F!����N +|�t4�[F��Մ ��{��=@+I��T�
H�66��I����6SJ��B�ɣU��k��}ᇼ��?��i�OJ���J�<5��m|�T<o�9+��+�ԁ .RBA�@
�׺�W�6��=X��>���\u�v}�k�4L�r¾O���F�G�q@�$�@2�~jY��~�N������K�$|`Ү���H\N��a9��&���5)��w;kk�Q�Sg��F�=	؋T`q���9���s|�3w�/^�G�n>��c`�X�kQ���s�N��fȕ������z����-T�9���+{�o��Bԍk�<X�TC��^0� �"���ퟢ�]�qV=}�yqH�1����b�{���'c(���u���ϓuݪ(#�]�y*�oï�MU�p�Z��/��
���z�:��`���b���y�&^v�)SӐ:�K�-J<�[��%�B�/!d:.Z��p�>}*�%>1tL-+���Sj�D�$=��T�;�����B�%��5�g�D�	4��bH����i��-4��:'�J^�?�����*��yR��YF� �"�2�']�aa��:$.�wa����z��\�� ���r�+�FO��	�}��7z�����ѫ@��T������G��t<q�A����S����~;�>5s��M8Uլ�H�7���,�7�}���W~�����O>3X��X�<��4
���&j�Oه8��6K�s�i�4ؑ\��UbV��&)�Rg�=���ٰ����FI�����3����tt)��K�r
C
��!w�9�HyB��k�R����ПN,Q,�_�L��m��=�����z����̝MH�����i����/_��X�rH0I*kw���k��xYj]�GI�G�r���t�@����Obj�n$��+�8r��tkVX�x^�q:�N� ���,�d��5���1*Z�w���WX���ŸE=���B�k��<���4��⫒˷��KW��]3�04��}�c>Q��Hԯ��$�{�K&�+��'a9E�����H����k�Grt�G����� �]�(�t�T���h�?���7�;�f�Oх���6.�+(av��F�z➻��O>�|�I���a�,���ٽ��Gܩ�B���k���GML2�9|��G�O�#x�>�u��m%�;�g���B�k�� z�!����|�x�i���-�廡��*k��3�H�?'�t�����Mz�>�H�O��2d�TLj�5Qɶu�Jo�}���N&���L�ˬ2��e�sqsh�H�r-f�</7���j�XG|�>�5�
�2A��s�ZM��":}K��4��2 ������
yF����[� "���$,�c��:�1ѷ��=��ކ^W�����y�X2҉�c[�a;��a� �Ƭx͐��G9�����وh�u��Ӎ
r��g�KO=��ғ����댧�$ht����P�&�Ɲ��wJ�39���7��}~��B]��)l6F���$�*�D�>EE�#"��Sh���)|�cc�ћ���T�,�uS쭩_ ��l�>���d�荔�ޡ��w�x������L�2�"ˮ��x�扏�g��l���
�oC�x�/>��z93�w<��6���U���@*�̔I�d���:īͦ�0�TǓ)�W��D�M��1�Ae֨N�W�;.B"�l9MUV��蒱`	dy�ۨ����*��f& bw1��dӴ�r
�Te&4��cKķ_���_GYi�8��"/c�u��j8���
�T����1���aqx�5/<|����=�<��=pj�:{t� .�c�Mĥ�
�F�X���b~�h�鍊ᖳg��?�rd�Mf��8��m��7p§Q��4+F�O{0�s�D'��n���R8c��MΝ���c�#+K
l�ٝ~J���pcj�ҭ��LK%ҙJv�
ʔ	V_u$/S�)��"4�LFd��8k�����{���g�a��æ�a�j/����k��}����$���*FGk1kc��A���FL�3
9��9�:���R�*�&_,�6j�����:��z�|% ��y�dV�y�����؂I�Ќ	3�TNg���1�0WG \]@Y�-E���n����o|�	�p�F��Nkn���k�2ԤW�����?E��vשP�\YO�sx��;@��)ҋ�PKA}.l6 ���H'NA|�K�A�\�㨠��4��ʼ@S�����m���a�&��SOrx�ou%�}D���ϔ)�5KǴ�)�Z]3s�H�0�Gm9��=p��>Q���3Q�A:� �zխ�OR���)S&����tkcki���1���6P=o�R?ܐdp\��ɍ�~��5��$Cn
X��0�qm��ؔ�mb��A&pjH�<������J�a�]7|+⊟���nALa�N���7�X
p�����k�h2��+ۦM.5�p~6���w~����஛o��O���bϞ:���&��5��w=�RV�G4��.T彡�T���J��L��jҞ�
�>�1m4DF�d$ۻ�[t+�6$�o���h��:�v��g��3�4ċ��[����*�Y1�E7�50\4�%߫��c��ywU�˔i�4d�l�������Z}�c���oU
� ��n��+{�A���E���1�C�<��mK�G�/�X��A��F�O�-Q���%��rp�Jr�3��Қ�J|Ks:n�#O�0��Ad) S�ңD]4�w�׫���y�qb�5ud�mt��l=YX]Ȍ�f���s��W��,|�ɋ��G��n;��O5zHi���rÊި����+����+��ԩ�c�yB12��ɡ�K���2��k��&�u*lC=�Ur�X&ե���8��/�:꘹�cD-�޷v�9)����s����o�ޘ��2eʔi�)�}w�T��H)�Z|����=pЂ�(5��-f�	�dͽ����+
mnw7O����|巰�<������o�x1��\+XX��p*d�!5�@�����.X��rG�L�Sz���
w1�)z����[l�ޟ����Rf�΁�k�plk�]��s�W���Ưgn������B�**����U�ٷy����k���	�:F�ho�p'�%$����it��K ��H���� ϯ�V~�9!\	,�Dd;pw��ڶ=��x�A�~��K�Q��]�q�lNq�6Z�q�(���>��-�����+������{��ם��(㒣2F�֮��4x���O�(�Ʊ�rca��"�m����y>S��������l^��
���[>�\Ʊ�XZ�N�PH���w,��o���\U���~%ͽ3Hq��4ȃ��]�
�7����ʔ�7����FZ�u|�Z_$�NO) �^��4��N)�C?�k:�ٿȟ��?E���3e��i�x9�15t�-0��C��$���}��mȥz��* Y<��+A�<�.�H�5��P�@��/���X1���U�b=�k�E#Ǟ�0H_��3�.@������}� ���0�����k�Ӡ�1'J��?��/*s�ׄr����o�h2ЕT�=�%u~]k>�zW����7
ӿ����1;o�����B���|�����~�q���۠,g_1F��*��e+*��Pa��
J�Eע�dpȆ�f�aa���M>Ͽ�&̋=��HN�7��IMu[B~��B���o���s�b�Lj��a�EX^QTet�w���F6~�@���5]m=�]�j>�@�h��)���^�q^M���Z��*�2e�t�Qjw]��1G!<,%.ƞ�@��e�`�`��4�-�H{C���FS�b�H.��tV�FKʧ�'e��H5
r����m��e$E�!D<43�;��)S�Lm�7�R�ַ�w��%{|������`@ ��y�+E!@1,���d�1���|�6�p���՞�z(-����|�w�^i%�2 ��>q2!�@ (��`�IS���u�18�ͩ?�6F�:��J�N��GFC�_o���.\�	�w�i�2��XطUe�W�k�B����8�wf_z��ç����n9�u1\���PX�̗���Sl5�+AYXk���
F�c���J�`f1��������~�|�PΝ{c�ۜZ�w �*���45$H �ʏy�l��J|��U dwS
7Oe7rp��8#��O�	��.
`xS�%�R:~�sm��,p{˿SS�?��Y�:�xc �[ʑ<��5�L�2�N�l>!!�K���q*}a�e��Kh��J�*���(�F^�j���[A�l�������`i:	�R��W*vUݵK���Xy������@$0���]z�|���u�G�E�B���X�NQ��TB����ce)���V���WE�'��Ӵ�=�g畫p��������=�\�p'���nd�CX,̆�𲡌�ͯ6cX�~�^��h���{�x�e�
��TZw��`����8��ү��<��M`V`ס��x$0>h���b�c�]�}����( 	#C8aT�M%���4�FɴRz7k����K�)'M���4$��]���ޅ�\����z6��֠e�?����y-5顆��$S�C�����x�T�)S��O�uj�wZ�j�)�F���x�x1���L�ɍ&9�iî�����~R�b���Gp(aî���P{��.�ad��|YamW�oWi��,�

ϻ�Ι2e:n�����H?bZ�0�b�, {�W�ځ@ѧq1�q$4eNS�����+A��T�p�'�#w� ߑq�Bw�p/:���j`x��n�^w|��$c�4�����r`�!F�:�*�3@�k+2ZA�S�0
�T�gQW�syZo�&{�s�^��P-��� �,ܹ����=�0<}�n���s�W�n�C0��iE���3�����N� �"L7��<mhr���.��ܔ2+�͏?��'���矇��J�:?��&S�c#s)q���!���G�o������m�s�^S�Z e1����)^C#��!���8=/m0﮹�GjN/N�dʔ)�v�j�F!u�ѣ�\}m� hg ;��k�[����j�֊QE��oNf'�j�k�F�:�K{��r���u�c$�����@���#�MPz�P�Q��i"lUDk]��ֺU��C(��mX�Q�|���^�C�&Ƹ�^K�<��E��>���J��w�_�ʗ�k�=�Ξ:ը�m�����*!ù�X�P��S_o�c�!h�t[E�7Ȁ=��׿~�E�g�ן�ϯ~{g��tJj3�l�A�6�e��5�Gc�t��F���oǰk�+��֬��A�����m��.R�0fy,H�BC`3� ��jZ�3`�)53�a2eʔ)e����Y��w+n�mJ�}8��|��|M��P�a"�d���:*�z���1��fʔ)�qґ�O>������Zk��e���J��8��&@b ^�y�N�3(��~}�aMT����[�~:!"(N:�K�~�ۣ�5R;dK�]"���ш�9�����v���5�FЬ�OcXa�B��� ���z����]��w\��_|��������������T���7�=���nt\�}���bU�q��>�?-��3��`�������;�W߀��>֘� s������U�w�)�ªV�
��  ��C��T P/@�J�LG�v]�01!� ��x���;J,!���׌u(���2e�M��!u�x�#p�S�KҀťL���$/���K��x��{�Z��5�^���]W.C�?�:O�'��V$�P�>,��rzW�����[x��])u�2E��q�{��1^_,�����N��g����#�����;s�ʥ�A{M�O��8�A�F̷�hm��;c�m/�V�#m{�8�2S��i��
Jx�Ï�^x����'x��O�<{�{*�y�����o�T�St�=��h����YÎ;$��F81��ё���[s�U�T�*/>�,^U�Zt�T��qj��!q3e���B�i���J{�:=JׯYx���<�	�I�� ��/�z�ڵ9#^SSC�8�K@�����O�ɔ)S���1�F�O��`�U��BŜ�qm�������}���e��6y �<e �� $�˞�B��m��၎����50B��Mu��MPH}�$��=)�P��/c&:��Z�zd�3�!�^~V�	3�^�V�h�Y��gG�4�։FnV-`�p^��<t7|��G����M箷wA�b�@ɺ����g����Ly����m����L��U*@t�������9�M�O//�G/���w������^����ZڵM�l|T�P�{���.Ǻ<MStP��ݥ>��	Jm�d�E��m�	�߸g��{
��t�vs��,S�L�֧��̾5x�k	�,P(�Ro2����g޵7���p�� �ݦ{,�B �ʫAY�@��"��r�P������nU��ğB��j�w��'�>1i�Ey��3^	�TW�5ưc����҅���D�e�Em.J)�N���MM��o�~������|��N��?p�����N���A�����`���&4`�vF�)�[�����6�7 �۳zϢ��o?����?�?��?��?���>�3{���۔�\h=w=#joM��3���� �B�I$u�@1����zN�?%������#���y�Nh`�u�5h��4b����g�J��z�2fʔ�X(�6��:�P��:S�T館��Ơ+T�$������*�笔$ٓ����N�+�v� +pTP�ͻ#֩�� 
���6�i4�����_�J�+{��kw�:
�b�-�Ys��jj�����fa�L�2]��;hi3��b�vZ��k*��5s�V	W���k��S���]B�VP �0��� �*�A�h]�.*��`����j��HC�f� �ܥj�t��&��Z��Z���w�g���W��9�Ύ�n��������~慆�Z�=gO×.���S���n��n��s3fP]�`f=c4�R]X	Ȧ[�{��1�/3�� D��wv��+�u\�Ǝ�����s6� �]����?�?��s�컿�O�M����LY������M6�����P>��d��u�{�Ձ �Iq,M,����yI
�\���o:'�m�Z�I%u��ۆ�v��ϐ�I���O�B��
�Cta�el�a)��Gh�5��Q/	��|�N\�L�2]{��B|�{yD�z�h�BP��r�����*�i3W�Q$�)�S���Ր���)I��`�Չ�u�������]�TkMUD$]�dS����gt%�b��Q˲�j�N��J�C�)$91NH����|=�JDv�+�K4��9����k�jlkTa�6q:O���0פ�gM��s��Gn:�|��݇/���o8c4��r�|�6��.@x�+�!XB�����L:�(��3��u/���&�(5��\Y���o���w?���+���e�g%�=x?�1�/JA�ͤx�8�p��@L��'��{����Eץ(�_��(�%5	J���9s���
���N;���N�ڕ;�	hR8(:Ҭ����q�Uu�ƺ�'�8�ǻv;.S���`��p�^�t�6�L ���@��Pm�{�	��R���"}�XZ��H}�O+!s��rR��ԇҵ偣vV���.u	]���'jǕg��e�L�2m#���H�)�^0_���˺I��ej3��&�P��x�ԻF�^zJ�B�MF�=b��J8��i)���ro�_�NI��A2̶���j/k!
��������^��g�˺��\�R�YU�-{sx�����~���Cp�����lּ�x�09,��k0[�kW�;u�N���ځ�¿������2@)�(Kг�}n�x�������o_|�����ڻ��w�|WL��9�5���jڤ玠��m���[��B���",\�H�C�"^�0'ɬ1����t�˥�Oߘ�A
��5�-�U[�o5��C��K��ϴ�2e��h�ׅ�\��Q����m��G�6&�ʽL+��� ���лA��k^��B&UR��Ih<-�4-�j�&��!�:O�7������##-�w�;k_����I�0�ua~/����fVs�5/n*��|����ͧ����n<s�����N�R���=�r�X6*�0. �yv��C
�^Bu�����*���a���?�~��7�?��������{������%���aO{��z����L�H{%D����g�S*�&��T�M�Iwx���S�=�x���LӒg	ߺ{�o�>�����T����̔)���T#y��8ᷔ���Fcʡ=`����$���kʀ�͘����\�(�1���P�L�2�G�5��=q9,�3MiL*�	�=6
���c������E�d�Mv�۝�r?�؀ MD
V�P8$� ��B8Nڧ�$��!נ}�/E��Y�ڂxoD��tI#.�%V��
n����M��W�~����;/��l� .��҂�����?g�I��VJ`��_�b��8`Ӟ+�iX��hzP�/�~��������G��>Z �9s�L{%9�!O�L���I
a��̔�n��t%��ӑ�
���L[B�����2eʴ��x�"�#	C����YvZb����-B	�G��*B}H�T��#o0��A�Z��1 �)���Hʈ���� ��c��㾫��l��Ȼ�!gD�y5�
ghaoi�pu_T�x�\����<u�}���?_~����y���Xx(c��AL�E���DՕ����d
_ �������8��&�&]�p�������_����W_��}�	��>�9�3noF�Kl��\��P�����C����p匌7b��?s���FO[k�&�� &���5*�D8b&\wǁL�2e:����ow����y��=��8�F���]Z[�0��Ɂ��S
�S
��2eʔ	A���	�8�7�}������P��}�A$Б��04}���@��\c���Z�^K��Z�Z��1Ņ�젢���*Fડ]n��M]s(`"GaM;�+O��|;���2^6�TU	e��t��'��F5�/?|7��������f�W%� ��];�Ԝ�;!�`Ѽ��T7����W�Y���[��.,6
�1��C]T�W���V
^y�]���?����K��;o���̳g���M��#ম3%�ݺ.��^�� p�G��e������:�[�^ZM�|<��=r��F��8�l	�Up�u<s��n!�����k�2e�4)i/O��t!�v��
#��굗ه�$X-�4�6����<�l-Xȅ�=%�+.�a�tX`/|�o�Y��
������b�J�E�ǵ#��E4�!Q'&u/����w�`�r;��h<nt!���^wR�9�y#�7��իP|r ��t���'�]�'>s7�|�~�ߔ�ء>�����&=������w
k�z�e�7?��,X(��n�sW�Y�0!��ޕ�襟��=���W^��}�\j�{�p�s��V��)�UhEm���+�W��#ֱEӷ�Ј�V��*�c�������Y2uz�����T�-�^N��ǲ0�CZ|	ʷ��͔)�	&��wsrq?b5Y.�i[1��i����?�G�����F�B˩N�E)&�gF��ӑ�,S�L�v��:9w�`"�B'wjX���r-p�V���o����+��m?��]���	��W�V6~F���FkbQF�?��2a�LG䉞�")^�� �NV,��)�;�����Dr0傠$� ��F��Z4�J�����u�@��384߫
��~7sx�[���z�~�����pf��@��!�wl]��3�p�1O�i7�G�ꦘ˕�~���n}]o�a,1�4|�����ބ��<�ͫ������ξC7�ԙ��?_�-}���l�ץ�z�=n��vq,����*�Ϥ����%�A/I�I�:�@�����2��6hF�W=��6 �|0&�U�7d�NEOR;]���0��� h>��`�l�v��Ͷ�"���y|�۽
fʔ)�PB�������P�LcG���D��6��Z����b�3(G-T&5\����ʇT2mļ=t��/m2w-jAY��<��7^��r�"YEJ��y؀]fǺ
�L���}+dߤ�\��Σ�؉Ԑ��x���I�+�#��N�^A�>���@�����R9�r@����۸e�Ϝ�r�������מz��.�p�<�˽&�F�Z�k!�Ր�OV멥W��ƶQ@W1���o[ �Ȃǝ��=z��e	��|��W�~�2|�߆�.}�O�6)�F5�[���Q���W���@�]�kq|'(рq�>*zR��֦z<wɴ;�H�OQBޏ���{->����N�E�P�A���6�HG��-�+��)�'�,ZW�g�5�)����L�2e�(���������t�cZݴ<.�8[�s"hM�h�+TXQح��
Q��R9H��Wa�`xY<�9p��*Ϩ2@��N�2e�t<�ά�*�J�&�Ly�U�y�@u���w���pY�@`�9�E%�����ѻ��	�D]�1�RCo��9U�(���Bh�CM5��w�YL����-p��j{���.�7]*�y㰆�
��s���-�×���ģp�7��3�,�X��E�����`��E���}X��A�(�ٌTi�oޙW5���\�_��x��_¿{�Y��o���8ܛ���9��ҁ�J�]���9�F��X�G��@ �u�����J+������0	���5��EM��-^���NmHMf58*�4�kX��a��$4o�
y�p�讛o�9�v�Y���5.���dʔ�䑦�TyAגA�2y2Z̚�f�o�Uau(#
�h�]�AG���1�|S�7�\���Vp2T�=�6��k������3(�
��`4�J�4B����z���A	���!;��p��׸�	����څ���5,7�;P6z�}f�1�j8��?��t=<y�V��#���n;w����(6i7z��ؾu��^�b�����Q�ژ��kQ���y����h(�&��6�~��%�Ƿޅ��%��O^��~�>|Ҕ��s�)��(vF�S5�ㆆ�>@��wA�}�5��������+�Cf9E}G}�����	wQ�XG�==�~�9H��܎qk�W
9�jl�LY�,`�)ׯ�~�4J�`i�^y�C������R�L�֠�R��k'H{�ye�t�R���JxC]׀�L-�;����ý�.xq�jXOh몷u�o���5����jla'�4)k}�S��iU��u�Z�]�L�2m7M3�+���<+9RYd0�{�<M���A�]��qS��
�@��b3��ӌt{h�ed�+�M
�X|�$a�A�MXE��Xw�Y���Q�E4��A�i��p�ܬ�i4�3� ���­�%<z�-��_�?������o�Yш�W����\�[��g�p�"�0+�4{�Т>* XP/��cxJ�v�<����x�o�_>�����7�� �&�SM�g�O�~ݔS�-餙�5D��mz�>�;�e{����@�GAP2}`p�ƕ��եA�z�Ih�2�z3F�'�\�$�USQQTV
�	h��7�^y%Δ)Ӊ%:�m~�)�8V!E���`�ɵgZW�;�#�.�@^�U*�}�
5�3aL� �R'/\feH!�Ԥm��N0_\̓5�K�i㍰,N�B!<�W��!�q��|\U��a�=�p�7���!���J�P6?�u��}�3ן�g�����zΝ��y�0:���ժ@�����i�1�U�ؓN�%x���
)��)�~�����33X�����������^z>Y�Q�LS��N�i5#���fu��z�SVǑFZ�}������ܿ��7B�ژA=�PN51�cƦ({�s7p��!]��+l��'#�̴
��#��$�ϔ�&}��m"��HgT�n��<P����#=e�JNf�)��n�W��Aw� �X`<v"+o���l���2eʴ��o�9����9E1�*+�5�x��2�R�!�}�[�%AJ�'��E��X�7N�T�wiw�X0-���s���,W5���A��ˆ�J�yèἺ���"�͏��� n�+x��-��'�/���������&��y�0^:�	
�x�P\��>����	''��f˝xZ�ڝJ�l��ӫ��/~��G?��{��>��M���o:�q9��Ÿ6��
;��Ɇt��'{ٰ����Ʉt��uB���X_ĝ��2J�cǼc�I6/�J.1�h�f�d>�,+��z�Mm���Ӧ�%;�� �ez�Wj�9��\�2eʔ)$�]�Pzоir$$��y�8�	�5i�؟'\�c#�m�� e�"bt"��"_�G9��u"E��a�9u4����J��+]QG�n�v�����kt����h��k��ɷRN'j�8��2�����>�|����{�n�ף�	h�`4	0�kWn�K�w��@�G���� ��
�����$m<�&�yW�t�����^������|�9<�O�&֔�,J{]�����+�$zT��X!�+�?�������Jt��h��^y@�ݝ����8��JM�W��ޔi�(y@�p�L�2e�t��7�#q��h-���R�4��Al�1��`+
�)�0v<2eʔi�����,���X�Kӣ]�	���"e�H�ۭu��J� �򄈯�v�����wMXf���"�+S����}�����RFao!��k�p�i]8��ʝ>3��'�U�o��0��#w�������.½������c=qh�s��k�P�ę)��� e�	.�[�7$o�ʻ��j��w��ֵ�;�.���-|���^y~��o�,`1��j�|��R6.����g���7�Z��b��?�×yf�����S��V٢�l-�xS"��;�����*
�!Ob�JqsN��3թڱQW�k@�1�ۈ_�-�GEz�˖)S�LGAJ��'�!lh}��N�8�R��w�d[����q�aBNd���[աӹ��H��b��/!���(��̣���_�".�I*_�"�v�A]p\�̣���8��[k����c�q��Z��&��O��/>v7|�s��#w~n����'�A����R]s�jw��M���:ɴO�E._z4��Ba�ҁ��m%�5)&X��\=��������7���Sx����?�W�M}f%�}8��s�u$h�6�\a��,I��ע(�Ԟ�!2V9�H���$��6>�@gv�Y�E���6X����;h���O�)e�h�zm�a�I �vL�庴�]5���)S�LS��5b�G���K�����;�4ڀÉ�|�rѦ̆W�1�*�L��ѻ���a{��8O�eʔ)Ӊ��&j{��lk��VB�a[O�%�ݯ&6�#���~�@3^b��A�j��̊2�W�v׆�frv�J�)�Պ�y�sF)��Y�N�)�y��AؤVϬ��bq�/��s7�W���7~��N8���v��������C��~�5ԑE���ޯ�=xh�01c�\�l5���FS�����ӟ����x�x��Kp�)��|n�6�x���4��$�P�uX�a�<2ļ`����K0�8��@JŪV�n}�U����{H��7<��u����#ĸ[�����{���18/%���Ewx6H����{2�I��Pz���7@�+oM�՟L�2]k�pÉ�����kf<g�"|�zѰ������$s�i]z0.�ճ����"�L�[��.�j>��vl �u$?��� U��ϭ�؏�_)��{/�0ČE�v���w�eBB��
�i];,������\�R��F�9���O�v5�'n���'���<	n��z�sJ��Һ�h�Y�RX���t6�>�$����~8�t��X���M�Ɠ��s ��Ǘ�?y��� ��Mx�rS����%���]F[��n��Yx���R��A4Ơ�ǱO���?��YwK�����B��'q�4�X&�v��#��P��T��I����5����Z;�39y#}>��:����hm>:Z57->���)S�k��>eLZ
�!�)��_�md���Ĺ@$ԬM:�����JW���^U�O�R���L�2e:nB�K2mI�Ħ:���������ڐ��ơ�_�������"�,�����#�1��6T_��[l�� a����iN����袂��A��8ׄ���=�\����x��ʲ	^Aux؄����CEde�l�wO��T�"�U%晽¤4Hh�-���$�R�lnR܇�4<������c��k�����ro��ga�4��D":����r.��K�'����Ԙ��K�h�A8������d0�92:�~��8�	- 3)'��)���|��R6V���pc��X�L�(��z��M��00𓝍72e�t�����4؎#;�����$A� ��n�$��b���Z�4#M(dŌ=��C���������؎���G���XR+��ԛ����l�@,�F\�X��[���d�̪�����G��{��2�2�*����9M���k]�Q�@��/�L�Ϫ7}/�Z�`Q?p��%�l,�:I62$��:H��Q�t�Q��a�`zM�m�����.7��֟ku�`m�	/L�r���WKdS�e���TƷ�6V�d}V�z͗���qu^�:7�᭷➛o¦+�Ī��:�bw~A{��4�_�z���zې�}a�C�^����t�Li:���)��VS��NY�v����m;��{�U��7����N�y��,�ֶ�kk���u:�7��[d�B�@��*	�wЪ��j�WV��&��p�E�9��<��<�R-�*�p:OX�~P1��qnH)�������P��\���MBBBFO����E�0)�i�b���Ǵ�[�.AԒ�					S����>����8��`Az�H'������5��Dށ`��{�2��)	�5�Ro��	5��>4*0E6Jn�ߊȔz�EQ�8�̣}~�0�ͫ2<��=xd�V�}�f�[�����.X����6t�g5�($#�%���+(TI+�OMf[��;���e%����g>ś{������p��)t�׃�iiC�_���,��1Wx�Ȇ��X~'���Z\��=#��o��Pg�V�d�B��J~N�v#=_:�	���#�Ԗ|c� n�e!i�z/�u����4FC��I^����\2�|��S��p�������\�H)���=p�eǍ9`�3݂�
�υ�]���xm)u��ܓ7a:���*#�M�hPU�n���u�/�~!qMk;���q;�c+�l���2m�x�^si<l��8]�3�(@��^�7u���L���3�=D�G^h��d�T��^�O8���~�OΝ/Ӕy�:�ZVk*��A���`C��p�k`.�em����M�.����
���[1¨I_g�S_���US���q�z����g2(X
����iD�KBBB���˕X� ��	�?&k�15mHʍ]���39A+P����ͭdBBB�Ł�ޫ��%�	u�C�-ˢn�+�[Ux���z�]L����;"�]7"H�sę���Q� ��[�'rV�a��a8��嗅�(������/�7�_��N�x�5�U�䐚Ĵ�Όt�o�`M����-�]���@&�ф�H�;��.�F%23V.��N~~{�}����S{��Щs��U���6�3�f:?-x[{��v�ev�u��c:�ʎ&���ܴ���,��A��u�d�р����L�g�x~�u@����`�`�����@F#i�0���A/;���]d������6�ǳx��!T�,NR�	X���nfa��0���al����S�㷠.�ˬ%������$Bx����VC�2Mrm5�G��"����z4T�
��Ba��*�_?�Ɨn�߾�<p��X{�*_G҆�]k��Eu��
{��U"#�R1��0���/�*�u]r��׻'>�����{v��w��G�]tgg��@��9(c�,�<t��`�C��zP�5ˬ����j:Y۵�5����:q����f]5:�	/0cM��6��8F�j�=���Q�p��$#��ì�]�					#C����D����m���5��/ɤ��F�yC���>��-�&�܂�kX-i��j&$$$\�WRz�[�ӂ�5�w�h�Y���0Ms²�ka?i.�Dwv���
�/����-M#cc�*��w�9JLx"0�����&�ʫ�+��ͯ�ҍ����U�Ǻ��
6%ǆb�x-~��G���[��5��LU�B�BS�:,ݡ3�y�e-�be�ZɌ�b�uކ2�le���A�;D��bF�������G��w������X��s���jV�j�Z�ä���V#�"�*q��go�*,������z���2��dU��������b�rY剉���I����v%^�3r��5I�$���Da�Nl���c�=ʚF��1�;T�"RZ�g�ע�X��OHHHHh�v�r��d�p.l����NZ�$?e0���&���X�>@��#Vnl��8�ɸ�~n&�$8���(�t�?�R�ra�{���LV�%Un����V���u���ΐ8m�s�6�q�%�!;�fJU�Y�;�݅�|��ظ�Z��z�)�k /�����:�j�[���X�i���[�6ZWQV&3!�|��e���$�|c?����x���p.�B��R�)�:/��\i5��3�2ϳ՟t��gӷ��]�\_�T�Y��Q��ˡޯ$M�nD�-Y���%QB���/�S��\v��'7�!Ac�=3����ߚ�.���c��w4�a� ��	+��"J�������0��&��)��z�0���<���p�ZR�x��2�&�Y�0��rֻ;�1S���Ǘt�])���E������FF���4��ٹ�۱/1�<����M\=ԿLp�84/���En�$N�F���iClE!aC#�mjwd�7��ߏ�4����X$(�+'p��^��mv{���9DGb����c���o��k ����Kt��SV���ɵ��,��w�8��RPLfI�fY���;��g�Rz��|t�s�>�.~��n���x���qF�hi��-%zeB߃�W�Z����F�e� ��	=��%)��Nh᛻�Yaf��ՋI�Ş7N�qR�_���Xh(��K��K��X{u�ɺ�P����"�� F&)#5�����q���y��}�n���@hh,ۮ�����:�i$!!!a`���ZO��/�Ik�D�P����d⮗�Wɀ$�b�S0��#�7	�P��1�!��B��oX����>}]�tM�}HV��������`e��*Nw��QIA��m�B%7D1�n�ciхT�̙/p��������vމ�J�<m(�D{�PF�P	V.d�YH��/��6,$���Ud�U�\���Ju��yT�v��]���x~�~�������I|T�]��[k�ȳV�Oh#yfŮ%P��x�5�w*��c����	�����]�����:������N���q.*`䗑�9ç�^�V.��@^��Í���<���6jۘ|�,��uqу�_���D<��������C��Rp v�xCIiB�/��B��ʗ~/X>�-��>&XT]�S�				��5����1�dS~S�j�G)ĥ;sT�Ҡf\z�-j(o���9��K�	x���B�ˇ�<#%[�%��\�=���RX*)����W_��W�*��s�L�s"�5]�_�
>eω<g�`�-UZ�"�M�r��VF]|p�^9��� �>�wO��9u�݆����&"�[�6D��a�A|[YB��
h�hA�s���u���M���#0�a�1NN�4<m����3A����.0��҇p*C��pFL�-vu���x��뢁J�=B})�3<L�qBBBC�<6�E@-S1�)��	/�V��)+�K���^:Om��e���;��V)����VsO��ձY��[(L�]�5G�-s3����-|u��J�ц�e:g�^�CE�7��u
x�{N���U�c�S�g�ȼ�2�_X�������/��Þ����y�϶ [-�s��v�Q�0��-�8�2~��2P��E��Mo�!|�j7�p�(�������@�d�l!X�x0�:�/�����N-�_�sO��WzQ���ՠY��y��餮��1���8��e�0/'e$\o��8V"�/��6!!!!�R�3�`�ȗ��?��&+�Ē�1�x/.<6���%��#��FI�ؕ6�$�"�Ky^�Zv��Г�N]�N��v��Gw܁?��_�Z�;oB���-�ä��:�x��:SˈA2�h	��7�yuu�E+� k	t[m��0�7�_ڋ'��ǁS�ͮ�\����sz���)�Uy�����V��c@3���MjG�ۈ�I	��C�tK+P]��F���A2ƻG9/�~���s�b0�&����"�[&�Y�0���2!!!�b���g�v���8&e���a����(��,��5A�I*��:�	-pV�C���)M���J�z��{���iV4o*X�����N���n3#3���}�Ҏ� :J�Ƅ�t�^���4F�>�$uMʠ\e\n��P��B��wT��v�̩�W�g���N⹷�_x�;����z���9ګW��
{[�yh�aB�o��|��%���3�}b�Ƶ�=(*}�teI��R%X'�Y�Ϛ��ޤ�T2���s��s}#ӓt�`0���/�p?�_v��Q�3JHHH�>���Tx�I���&�(Q];���! ��s}|Ȅ�����Vҭh,���Z4�?��"���飯w�IeWg�?e���	0�~3�1H�GQ��B�b�Q��H������<���2�����5޸`e�E�Ȅ������X#�
"(��2C����x���%��9�W�}O�އ7���c�����ج=��Wj2���<��f�������%-�A�8l#�׷�?��00��}�ߨ0�!�){���{_<�@V��.�7��TF��~Ӆ%5fGQ�@瞂�7OfD9r�L69/0#ӊ�s��cR���������H�D� Y8��o�-0��8	^��7ѹ	n�<yHʿ�޲�Ѕ�SQ�y���>ኀoom|^И�����k�xc�<TH乱ذ���v�����G:���&���6�\��L�;S�V�6�^����N������}������(��֬�ܪm���{�r�Kg̳��w�w�N�p,��]�P�$����7�k�^�}������Ґ��0��~ �W�V��쥮��<u���9�d��1�y��J��瞼D&�~�@�t��"��V.�7�R�q���#��co���p0e��ډm ��bM[�MD�����xv/1ֹ��c��}OHHHHXV�Em�cf��,U*dEfw)�'#�!���dp�Ǟ��U��V)v��)or+�^�����;��aiz�D���<ydɬLsA�f�*l]9d���R�bC]k�Q���SE$��C&ux�3_���!|�ڑ���y|޽ �����9�f�
�w�iw�������}UMr���]OnV�@��<"j�@���d�1Xv��/��\�E���[<
�(�l��<ǟ�;��{զ-d�I��PY�ܧ����Ç0a}�OQ#����%��R��eBBBBBT�8��Wfrl�[�9�-p�2�ಲ�ZL6����ʬ�V��+�PQ��­[��F�+eJ��l8C�Pg�˶��uzi�%J�[�X���s���8lޒ������������ks�y9_�HSzE�X���7`Nwf��A�<6ģ6�(��S�� X������.�X�p�ӳ��W������G��Y�S�Z���fW!W:N�YK����,׸4���C��7�'	ذ*�J�Vo���8�/�
�E��O%_x^��;:H_�O��h/Ԋ��T��s����4T[YUe=���IXn҆Ӣv�M�				������T9����K���d��5�zw9�� ���_�����C[:��P�������@Q���:!!!a项>Ani�>j����+aX4�S0n�;F@P2҇.Ap�7��B�/�V�c�ュ^@U�)�nD�5��!�熎%޲rxv�k���BhGB�"BV@º*{bNgBaN�xu�~���/qdn5d{��Y)�[�,3�83R:��Ħ&Q2�6n��P��ɚ��i_7�b@#ޡ�8�yE�4�>2�0�Q{�s{oĒ�RK��Q���t^>�2������V��J_%LbH:DBBB�ʄ��+\.*cL��]�;���^��n�[�Eb2'�	8�GJ�;���5�hU/
oK߸w�J�M%D�q����M2���tK�)�(��+D�a��u�3�g�=Jk0��?����6#2��_���?��|m/>_{���X�<�1��K��P�Bي�}F�*�u�c�̇$2����Ἡ��f2�Qz`����k���d�:��R<�&=���\�-�NԗR��f��_�I�(��"��r				�:�&'X�!�G&��[c.K���dP��h7�+A�#�Z�����~2�HHHHX^�[a�tSC ���H�g�'�Gynί�K��N0�`¹���]�iW����� ��L����;	31���j�嬶��g�vQ�KcP��E�Ղ�DM��}����
K+d.�gm|y�6���|��K����S��+��ٵe�]��\����J�� ��}(B�H����p$��r��}�[-�2��+-�s�2:�A�-&"%�|�%j��|%��4�K��\�Y�A��@\������p��~�p.�7����/� MA=�t�I�VŸ5�R������&'�k\&�aU�޸A@�ȞMb������e��\�!�<��w������
�B��v�S��g�,�!�P���/�q����/�8���w���dYVw�]��C!�:4�22�c��UAʜD�g�tV�=��,�ϳՍ\�Vi�s������� �Y�i�l7B�g���(����w~agT��K��Yc�J4�:,x(%�I�_��|�$$$$\�^�ΰO,�6=��{��gy�R� ���;a�+��h�x�jF�0��g�������B صC�ƓuH2M#�pzkn�� �~�x�-�G\��󩗌0�8���|������3��48���F*�"�¸�V�O|v�:�͗]U��Meɐ�7��2�j�å;{��W�	F��U������+��]x���������a�''�����GY^-�)��j�5�Ȕ¹�&;Ya���`��\Hg�\�$qԒt̟�T�l��),q��8wQ-+]��Z��Q�V����Źr�>������H�6Q.��N�=&$$$$D0r��OV��#u��fѸp�fuY9��8��Xhj�&���߀p2��z���E�@��\'
d���X�oܜ ^�'cQ)��O��i��"'�6(Djc��6��v����W�&�usmt�yo�P�R��z]��,0��e���߈���9�������x��O���'p��Oq�(s��J����P&�]md�Y]����!Գ�LDtݺ6|���(}��Q@���^� n�Z]��_j�Q1؈���)k�֪��TW�:y̯��}c2T7�ϛ4!�h�wg'$$$\����E�J����s/BE2��� ���XL0B���V�K!'*���-�ę����� ��I�HGd�"K
�0���/�ǔ�4�ے/2J��?}��H����Jnq�H���`\q�gJ�I�z�i�n�۝�p���2"��\)E{��򎏓�3$>;��ۇ��<���2�,�[��g"�i#��ۖ���%���w�޷��. �;�v��ض�J�����e�w�S�x����x��S�t��|լ�������@Ԙ����˲��;��%�0�`�!�yvi���p,�#&���r�50��k��
s�3F�F=�{
V���q�;��!À��#�Q�l�@X��ؐc���7�A4�����j�p�.LHHHH+�kwlE���v�\s�k�����C�l�/,�
��0��MXo����4�\l1;6�r� �мξ����,K��A>�d �:O\-?�[tF���8o��W���Njo��^�$�@Icf �@Bj�Fm����q|���8w��1��
���
m�T�0'��󊡲+��S�C�Gf�v\�6�CWm�÷߈�.>>{��?޽?;xo~��F������ѫ
�㐾C�����l�����*�B��68��ښ�J���cy3~vxۋȘ��&������mXИ�����ꧫ�@���k�T��48e8�·P{&$$$$�>;Nn.[���`C�殀)�����9m`/��rDLŎl�9�̍�>]��d�l�h1`2?	z�����Z�G��>൰��d��{/���ݞ��~�qZ�?��x^`�88�Q9�ɝ	�͕
,5[�,8%�x�x����ӈ��C��u�\�*-���^q=�q�g�[�^Y)�������7_{�t�v��z����Rg|�A����1�$����r,�Ew��Fy�X��<���6��n��>��8p O��O�?�Cg;�����3�Z��T;>�9D���4�e����&�B�i1&��jp��u��G�X�\:���p��P��>��O}��W
���Z����Z�$�qL���<����u��w9�Xc4,���́���}���Eʌ=+����=�[h�v���LHHH�%�5�p;�-���Asi0Y���H�z��U�yex#2����C�O��$����a%2g��S�uL�t˷�X%��^%���7�-#HGmSS���/��gd��J*���Åz�q;+���O�~�������+g�J�a�~�2x񜂤hC��$�y�3�Y�\�Uz�PY~_P�T�lgW��ƭ��kwlÇ�����Ǐ^ه�>��/t�E��u�9ڥ���;(2s?�G��|�qo��=�R�_X=-�1e�y�B��̵�"����i�K-6J]澃}���t:j��O�m��]�����%��gc�y��v�&$$$�z�m��s�ˌ��]��u���ʇ��.6��l��s��d��ٯI�N����������� ���w�df�+�b�7�kMm}W���,;O�dOL"Q������1�>X��n'NZ�|�9ϓrr�q��GLhVn��`eQ�Ӣ�lg9:�-�p����-��_9�Gw݅����:Z��q�v�Ѯ}
$���eA<y+��Y 6�I�#�F�V��u+��f��8|�4^?|��;������Kf�Z(��ޝ6#s�����y#Vrd֨V���� D��7�	�8�B^ӌ��1�o$R�q�nw ��}��.�ϻ�OWGd�����&��Cn��S��3$hz.q�b�;��V������݄�����A�u���
~��~���bs�t��8�)]/9f ��_��7"w��"}%V���ba��ķH�(��k��c������>��Q�aYdV!�ܞ�����ϵ񽷏��W���;���֢� �g>a�j�'��{A�e�4{m�N^n\�cJ'!ofoFn2(
d:���+��z �z�����{�#�X�;�8������r�e7��`}F��Z��}�e3�C@�z�s��N�u�52;�<����ԁd�� �t��<��{-t�(��Yj+�u����8���	���R�b�D���I}����0	��|9`䙕�y�aĶ"��4a��7��bq�G��H�������0��D�]v���J O�*x*�$c  �K^���5Ǽ.�	'N�Jvi��(e`���O��	�۪M>�J���iK?�YcL��U0��&��7�6.�/�g����w���{��=�m7m¬�ݝ�|����6�L�E��&���Tak��n�Os�2��s�X�z����C�`�����޷���wq��i�8���\@Xi�rd�R-c����0Ű�&��4��mgD_W֌to����f�m0���JLI{ۊ&���'2�� ���!H�p`�kE_���R�^��)ue{�>�[�B�<�M�V�|�����0(l0!^�Yc%�S��������F�5���3U�~?2<�Ґ�Ⱥ{��F^�<�Od�0��<m�6��w�5���BYav"v�U����ӷ�b�{��;�?�oܿ�\����W� &d����"/&��B���C�1�A;�񋰕Q��g��j�q�L���ڂ��؂�?=����S{`�����3gp���|��t����H���đ��*�>%���tk��ՠ>���ZQ����*X�ǽJ�v�l�<�,+:����v���c|��,�I�˗�}�;�|�_�����p1`�R��app��!e��U�v�2K+`���2��					����{�t�e{�N�1i>;ؙ*�# 6���>X��\�B�X���u�8�v�IN03vo]]�g��w{*D���5'����NjG��2���D��9p����؇g_ۃ_�w'��.��V�me�:*��1t(
C�e���7)
SaVEHg��Ŧ�ڦ�A,�K
\.f��-���m[q�<w䃓xj�A<�o�|�>���B�e�̅&�9;S(�"��+ld!�D�X��S��0��;a܂�*V�eX��݇1��h�d�n����`�Ԍ�Ų��!�L~�]	u����A��������Qd)�[�� ��@U���$$$$$L1�!qS؎��7^M�v��x��O����Fk�^��r��r����9f�R5nd��"�Y���������=�N�x���O�2F�db�Q�C#'�ؗ�d| �g��D�����-�WΞ����|�E������=;�q��h+]F�0���O�?���Jʼ	���|'�1 ��1��X���Jͪ�[6]v56�5~�q���x����Y��=�m=}gJ��h+}Gt�-��<�u�2� �Ǆ�3�c���A�A���7ʐ���i�QwK�_ͣ�[D��g��pF%\���Q��G?�xz]_���E?WG���$�����������KCp��K�-EXQ��^x
b�6U��q�PJ�7�6^��&!!!!ap8�H�ET�mU0�L/p�G�{�ܤN��AU1�2u�Q�rDJ�{�L�ƫ�'���>oد�{�K��u�y_"���-r�{�B(b�w%�h1�@�gf7�r�[^0W~W�9.�
� ���U��+�pۆ���];������ǚ�L��k�(�An0����~�}�v��I9j4�OcaaΫ��EG�̕Ƕ_{%��p?~��{���xj�<��~�z�#|^� �R�Q�B�s�|a�)��SM�*�L�5���4:D�7�����rQ?�ID�h U�qN5
D�-$�S������a!��b���!.ؽ9FCMD�}UŒq����,a�����@�%B}Hf���ҽ�����6����J��<*4c_��F.V)mjQ �+��X�d�v��4҈�9� �G8��#iW���&Zz����}|�U�T��wW�30��� /xA"�]�CI(��9�"�2Cun�<������׻XS�Q�����Y���O���=����߲	�ݽ�n�׬[�Yu�E�,cA�mu��K�}]aim2\���C�2����*Ji�t���y���۾_�cΜ}{�=�'^ߋ��?���.��2Xo��͕�cBG�V2^:2k`��&P��
XOp�<�Ƣt}h�F��3��x���ߢ�wd��N�^��UT�:hH�6��1�=�8��?4��HX�
,%�~+�N�Ш����ux%�5!!!!aj h��.���x啂E�A8� ���٣XT���*L��߄!ǰ^cR�[�W��yŰ�ufw�hM�p�n�ڦ�K��=}5$pfFz.IDg,;�|�X���7��s�kDO�¬�e�1	DL�JS��#��(O�`��8De�1;��������?�+<����K������m���-����hʹ�Ք�2�0��v՛�H_ϰE��ո����-;h�Ƽ��Z�z�&�z�M��/	G>�/8�����>���*�K��<7u��ؘ�,�9���=��췓�m�["���H|����ɗ�\:�w�5���'���쳮�}V��&*�~DTN㻩_Թ;�ߓ6�*�ʨ�K��+���p�B`T�=0���k5�!�
�6�����M�<��p�a\2�M�=R�HH��R\*2ܨɈO������dt��Z�JM��/� ����F �_�g���,��&$�R��/[�/��.�����ā#�r�Zܿ�F<~�����q�e���}�n�Sj;گ�1S҆��WF��G27w���ua�'am�
�w�.f�sW��_�q�|�v��S�b��K}�^:|�>;����t[mm��U���?��FrC��w�'�d�a��q�}����:�R�<9�X�Au(,R�X0���{z��I�*O�]��'3��S�����0���K��Qٴۢ;�:�B�k�Q_b�TYc�I�7��Y�┐���0~��&����v���wP�c4����˯|��F_D�S��12��P�����(��^��rxW�~֝'���`���	-�J�L��HQ�~O�I����٩i�*l6���,�.Z�dV�(��;�/���C��k��!��w⛏<��[n�ի�0��3�`�IM�6�,`XO��h�:�#�xf�z��*��U�o�F�w�&���;q/�݇|�-���$>��bf����IGir�¸��[ǓV���ILXr7��U:��Qs+Ψ���\�q��Cn�$\,3n�1����T��l�A��9���8o�����Q﷠�������I�PѲw�V�0�c�2�$���Fh42Q�������!�yk�#i�	�qH5��X'�G����^ω߰5�5uo۟sWd��hb�ˊ�/f���b������2�+'>��>���g�����ƣ�v`�5밮=���rҵ�i�p��~�����T��ⴔ�ǅ��������
��ڎO�8��G�œo���o�������|&כK�R�0��c��,��D��c�a�"[�����!����ן�Վ�;X���Y��F?�� �!���W��Z19������?w%$$$$Lz�U�P&.�ah�s/gs��P+"|�nB��_����D�.]��&l$S�y���:�#�`v���q��
�`@X�s�߸	�xV�*��ѕ #8�3����G��L�4"�Rrr��!���Oc�k·�AS>"<*��5}��VX�#א�P!st���@6�C�\��e�?� ��[�m�|�;����΍�j���ht�����xf䜢cHA$�k�(�PW�N��s֨"��P�tk�dۮ�[7\����Wp��1<�� �~�m���$N�e}�/�=3k�F�&�$:�Ȕ&O"x��'}mg���^
��|����C�("Y��R����k��D�D�4��vT�0�i7�Xj�4^h��Ǌ��XLHHHXj��=SH`2>6����N��`�4���ڕ�����K���n�!N�,�� ot�0�?t[p�+ㆡB/�mxaOF��������.��x�Gq�.|75��Z��(y��h����v���/u�Nt�J/�'�S�6�W��K�.^�����~���t=~��{�՝w`�UW��A�naL�3WV�|�U�\��Ofӛ�,���h��u5Q��kfgpͶ����;�oO�������{ṷ�S�p�ԑZy���ͩ�w��T�u�J�.�������
�-J��1���Z��a/u�1/���y5�#֘��a�d���DM��k9H����A���.*�y`�JHHHX�V���}z���8�+?)�ς=%��Ў���yQp��p����F���				ˋq��^�DX�f�u*Ed�{OS��@����w�\�)����@Y�I��A}�4��(�8���<h����N��4n��}F�H2��?T>J�g�w*ǣv� Oʚ�%�,3��v�1����\��c<3�L�j�Z�v{����n�?~�U���b��k���[��=�������b�L$3JP�����#��р20�!�
a�i�s���eywm܌;o݂��k8��'��λx���x��q|8�����\����3<#�S�B�Z#�T�na8ș��>������s����uԭ�f��}��!2{��8<D��U���k��$Hͥ&K�<p�yq��7'�$]��d"!!!a��W��|�|׼Oͮ狟=+��c�#�.*6�-��.RJ%(?��?ڣN5�.��}����@_8�:��N�낊�v	A��<p������iΓ�傲��&�߼�z[\f�
J%�F:��Z���&��T`����������k�#l��O��-��Kw���۶c��� ���Ci�-�U���u���4
�1ذ�2�����6Y�_�R�0�߾�<��n|t�s�;�!^=tPs����)����B�*��Q��~yo�>�xD�g.�� ���P���Ì9����P��n�:�N�W�1����$�����h��o���Uu��ތd�Q�k�E���yHϥIיU����4��������qU5�i�`�c+;N��0��D�؀�U]�@�\�	�{�п+���l=���)6ޢ�����t�����1޷����,z�A!�J	���'M3!�R�m.������s�Oj?��[J���Ɋ��l"��6	q����u;��adDzF��c�]oNܱ70�)�5&¢�������@D�H���*���_iTnZ$,�D#Սq;楽�BX��Ҍǎ"8���6�,,������=G�������[���;p���p�+�9DA��n8b���ҺZk7��ߛ`cK���*b,�NW̴p�M��-�ⷿt�:�~���l��{�,N�_�B��sb�<�ϭ*O��X�(C�B��g��q��PX�YD�jӰ;��A����j��9���M/�8V�� ���Ua�J��k�OI�#/�oNeDmŞ��VOz�Ke����RY!iLO����{�W��e:u�i��Ƃ��м�@��uF���kQ+}����j����"�2��T�%K�of�q�#�}�o^�C���I�>�M�\Q��� 'ul��|�d�\dG�v^:�.�����\>0�<;&�q��)�0V30s�P>s;%EP��<!��Q��ɻ�t�]U��leԎ\{ �V:@�(����t����v�/�ߍ��+��m�������U����!�7�u��;�XS�j��GJ��P��hʸ^b�嫰�-x|������t� �������'����l��_(��L���t�Ύ��-. ��̫����1a]�0�tdzE�'���w�u��q�%5�bԍ�� �*�$�Ύ���7T8{#��D��\�d���j��^����7�T�
4����h�Ŵ�Q				K�Qy:#�ŧ���}9Cּ��S6m���<�	�iL}���"6ߗ���+�*P���˄������Zn�)Ò,���3?���i����("djBs�����1��-����Xl�0g��H0��ƕ#��d�>b9Ae@��5�<�_��� ����(��
�S�-+�0C+��frӆY�FvY����!���{pۚY<v�V<z�=�y�-X��2`~��>ѫ �!� _`l�_����%S%�w�9�O��q��^C
��*1��7݆�7ߌ?��G��O�yO�ދ�?x'�wQ̮*�C�(.���ږ��U�iǔ��Q���65���^@�����5����Կ�rI�����m NkԻ�����hw�ʷ�\��aH]�I`9»,�WSN����-��3					C��=��-	2�4�;~��~�y�8���>���m��2�ui�����M�L$��<Qw!3��R��_0�I�m���?�lo�lҕ����~�9#�oe���3��@.�1�
1")��C)�k#�O�/V;Z3����������Ϟß���������;��=waˍף����-D���)j�~jڐn���ڠ��e�=kXμ�Ȏ1�~͕��{�wx ����#��ī{�Cq��)��9��h�f,�ujYkcx�u/m��tW
Nj�S������"�����#ݧ�M����>�Fɘ���x�&){�ѥ��Hz�,~A_3�H=����0.,�FaeZ#"�]&Ơ���8d)^��|�bEA�H�uBBB�Ō^oz��-�P�:ByƝgD�08��,�c'�(b�!����Z"�?��uu�_Pv�IkP`�Q�R��@%;	���>�ld��&��x�s��L��N~e�e9�H��������5x��<������_x7����܎G�ށ�7a��9d�3���2��%(?����tߕ�<��b{��"eU�Ct�L�af���7\�[�{ ���{�މx歷��x��8[^6����)�U���:�PC��ٙ���Ƕ���3Mۤ@c!��Q��`�*=�جO�����j�bk~џ��A�o�cE�+n�w�]�훐��0up�K�+�h�vl������^�u�����<pD���f\P���`�]���"+��8�a�o��B��d�z��c�\L�aoJ2�SW.�դ4���g��yFr���%��	>5/U�Bo��e�[���w�tJ]�d���;~�?����Ӹ�����]w��;n����vF����O��VÆ�d��Yk�PgIy�v�DT&ݎY�X ֵs|m�|y�F�>��;���O<�#g���*�3��NK����)��2�P.�]��l�9�
�>Ԋ���re�>����]��R�:�}��߳Q=FcaƢ���u��	��ڄp�.a�i��!�r/X㚳F���RP1Ԝ�mp�~T$�$!!�b�R��z.���;�	o"
+0��AS7��;Ble�;}8s�=؜ּ������u�Ll?g�����M<֑=�J5��qOv�8��>�}Ć M� �Y_c��w'I�S�eǼv���~��A�U-f�i�8ӑx��^y�%��_����Y�_ٹo��n��֮6;�4�����L�E���^��R(!�I�<ZZQ��v����������m�m�o�?��8x�c�t�(�?t{>�����I��VK�]�8��dt���LxWφ��"\3���u7�UV�=�Bn:2�|��Ƒ�OL|"��`˾:%B��F�eE|�NHHH�>H�l�1����t0o���b"rB�-U9������v%^.�sO}>�Ki��������*���*r��&c�RE��������Il�!$���>��D�m�v�gë����)/�R�S,�C�R�_3�N��G��?~�����O�M��v`�͛q�5Wc��DW�������I��b��6�-|�
�THbu��͖��^}��~��u'>��$v� �8��ǡS��Ӆ��]Q�<ʚ�Șو��tՍ�Cu�1�<ag\�[�uN����(�K�˚?&��{��wU�{�!�y��><z4��!T¹xd\
V�				h�$��Kp�q�lM��Nܮ`f��/�Dބ������wڸ'��Âu�Z%�(�t�T�9����[����bX��e9��砾�u�ix����{�D�av*��*#H�Ħ��	��&:���n�����1�~G�'8�1g�Ȱ��ru��jp�9BS��d�`*��˟���[���s����E!�8�����z����2�h�$-Sk�|����}�_|��p�����7n���Ư�{/6mX��VX�0%��y� �P��e-纒C�S�~��Tv({�N�|~�X;3��nڌ�n�	��<�ѩSxu����_�Kﾏ>� ��]�F��ȳ�,���m��v��T�l��;:ċ`��E���� ���WGn���}���0�1�hz.�1��yЮ=GC�m��d����8���{��G�!T\�E�}mB����l�}�=�_��hj��%O�0�%$$$�-�xcۑ斌/�B���g3>�x�u����P�|{	��G�/�U�Jl�bQ0��D\_0��I��Y�&��f<�x����7��Ke�AAʳ���N��8dW����a��Ӝ.�D^n�r�K�Ñ���A2,1uU�O.��|�	���A�m
(0����}����7pÚո��[�/=��n���]�\y	,L�*�~Fq(L��4!]��QY;H�{0����57-u(�V�aݕ�x�U��}w�Lg������܃xy7�9�3��\Sޏ4F�*�J��BL��:�L&��Sx�i(���[��$���U�X?�&�,B�����@����LYL7��~�	A�M3�=�s�X�??�${~j�V_'�I���l�&$$$$L���|Z;�-�MnӖc�1ȀC;�+tv����5�[�V<���M�pIHHH&�^�{����^�d#��R�"o*eYv��m����=�iM$���L�Jh�ӓ��\��J��:W|L�����r��A]��� OO"��Ⱦ����d8���T(�d�-¸4��[�T��{��ڡ�.�@�*\q%>�,���������ĳ�~�Uxt�V|�{�嚫17�
�B]LfB���e#V���R����NL�qU\t3CxfR��蚖�-k�i�Zl|�~|��]x���x��a<�� ���Ξ��\��f��S�m�t���--�K�3C�[�?9AY!�m�32�ك
�J��CA�^�u�V]��N��S�:��r�P����				�0F���!$*Z<�h�����i���t�b�u�"b�7$[�n�B�H{�|�0��ׄ�DT�)����t��;�m�2�u!�+���|XY��8A��|g��.��rȋ�ٝ�x�ƻ���<���BXmO��+]퉳��.0�B���.��[��7a�kp�����w߉��؆+/�h)%��#s�D��ڤ�-I��-T�j��+�dNQ�jYS�� ����e�l�wnބ���/a��w���#xj��>�>�t��lsk�@�����U�u�,gz	ӯ��A�s_�냱m�<.~0=GƟ�z�Ş��k�ӎ�:����a@���ݹ��L@��F}z����=Ӣ�%$$$$pε9	��Mb����>��8�ʊ��%HV��$`+�(�2������K+��7�i����Pa\s��w�cr���8i�Bz�0�5�P���� e�*8�n-~�QjU�"�Dd� �M+=�������/�k��]Iv�@�� 6;Մ��1�_2CV~)�1~i�[�Θ��-����)��ĳ�ӟ>�]7^�][o�wl���q�����B�z��q��L�S���킩�^9JD�Ո�-�o}GV�n��:�r���͇��N��ko��o�����Ǳs�!We:�
�һ�`v�e�Cӹ���H��]E��_0i���ģ=�M���(b4u�r��=�=n,u���1����>!!!a
@2_���U�e�d\\��n��dP�wD �jH�?��z�9��s��3�g�,J�};�
#]�R�P���H���} �P��,�!	�y���+�":��0L��5�P�r�V2��U���9�>WZ@y^�P�3��5�ʱn�wŏ��m����[6�������p�Wa�Ղ�:Ԋ��Au(��]}ɟCuPy�h�7����u��O��+�U���mx����ˏ���'�¾�x��!<�� �Δz�	����һ�Sha�G��c�(^G�U��zx�R�xh��R�#��w.-�6��A�걄%�5�`�c�觟R?&$$$�`8.],�n3=\ߊ2�p�X0�MRJ&��z�+~ɺ3!!!�R��Z#2$�8a���I�,i�ju��#۸�p�ؾ㮘N��`2]O|~nG��o��D���>�X
�ދ�U��%�&�O���d��JJPf�W�H^R����5"�jwZn]����0aW
t4	ڝ��{�G���>�����|#�{��Vl�������-dѱυ���s2�oz��%�0�1��K�9Q�|�faU�UH���y`����5���}�Η���>�_=�3|�ͽ8|�,��נk�	��H�%�m߲��sH��û,}?�=;���Du��)���٥��72�'�K��xi��eS�za��Tx����������A�X_s� ��fV0��z�H�I�O��L`� Hư��L���2^^k6�9FI$3����<w����z��t���D=�1Bp�7�򪑓ٕqU�J�Z]\��;$cI���`[׵ ���c��m��W���u�ҫ��_݋����՝��;���M�q�U���ZV����{2�h�J�����~���5h�aZ�g����<ǽ7_�{o���G��=��?{�=�33�U�lJ�jg&�lfu�L�R~��4FP5YsmS�#s��V�������t�.�t��ˆ{��0�5!�si"%$$\���<.d�a�m4�Ji)&�ka}Vl���b0!!!!a�h?�.����g�?�Pxr��9'V�F�����Wvp�|w�c�;3�:�;��p��$~���0�2�Ĥ��	ǻ��h�[�Py�*�{�,������.��6�6��p]�����W�porX���2�W�\�O�cE���V��[ֻ�6�cff-:��m���)<���`�?� �n����.ܷc;6�xfm�&F�	�b�U֦J�,�1G�
���dl��E��p���NY�[�ڈ?�������'?���s����,��v|d�m�.<�Wr�ڨ D/7�!�"������Lv�4�t�c�6gD+�P����d������{�:,v~���rƓ�8r	�"�[�M^���s�O���<o%ke���і�$�O�Q�`Ļ��1��������uYz��Ly��� aQ=(-�o�a�F>_�78Γ�ʓ�`4"�w��%��H���ϊ���C�)�+>�h�o����y�^��%]��c��RgX�.�
�c���w�A��ko��Y����ؽwc�m�b��#�tu�ڧGaY�9�d����cІ0���'�IR2ȯ#�~�V��7v>���u^� ����^��t�Ρ[�oYV��*���x�Ū���,��"�c�Oc�ޓe0�B�'�}���L���ЬY����\���ؑN�#O3�u9�^Z�翎=�)���؁����ޘ����MG�9?ِ��ݏN"��z�Cؕ'�W�1��~rȦSB��Q��;A@U�v1ޭ��eM�i�NHHH��E�3g��L���[:��.��oo5؅k�زmE@l�&& ��6��#6�=>c����*�a���QF0F��"�9G�D��'�-5Y���y�9���ULm�ާ`'�eDn<�j���!�@�f"��3^E�+��*h�¹Y�o)�Oy���o��ڠC�?t�m|R����������3���k��w����b�5����P������3P���8��6��!<���p	���"Ǎ������������)�ΟAgnU�g[������ x�s��G�u�C��}Q��7��u�y��Zb���L	��p��5-Q�gv�M#�~�8�;^�{1㌺E~��C4�����|p�iD�Wߍ��$�c					�*ϭ-7��$|�g�F�J�I0�LsON>��Q �G�C vNI�iYF��s4�8q�CW��}Y�tԖS����F�~�t��Q��I�E�P�qE7�x(q2-�ׁ����̚��Z�T��0�
��g����������:�k�[oĐ����L{�(�?�л-paf�v:��/�������_�/�r��s;��&�_���ҎJ�NvC���ƛ�Wn�~�oǷ�s�A��nW_8W���;����� ����?�֬BGΘ�E��e��r�}MLD0��n�ћ���;.j��_6�Bo�	�-�S���(�~�f��������9EQ�rӽ �t�Ľd�.���褤�f�&�b�Y�署�i��܄��"Sc��q������S2%+��(�Q%�1���cO���$[�	�<D� �d�a�<�_,�7*�(-!/���u���2R�b�yQK�4�"!!!aA�b����������k�@��$�n,%��?8-#X�I2���=��C/�z/	�ƕ��9aV$�e8�I|�5��N|�c�3/�1��}��� #��2F��_I��-W�w�t�%���\�(ʿ�2MG��X��9��x���x��1\��x`�u���;�k�M����07;�LyQQLhg��@���3 r�4J�q@���)"�#1WJ��nێ3���/�]�J��&%~U���N��5WvW7J�K����>U�h4e�ɐȦ���b��R������k\�=9�����:b��<�!�/t$$$$$,<7�ỽ^�`�w�󍺄;k��ƵF�Z����﷗6́�V��^2����e�Eg(��H�d��H��y^��:
�j��ɽ����a,k.�����Vp��ɒ땂�Gh��{W-�k�����]����q�,�|���k{p����[o�/߳[6\��׭Ì2��v�|�Yk	����4^;����6����t���wf؅����k����8��|��=XX�����r^b�M�\��z�&}"�,z��t!�s]�v�}F����G�K��\~qNskI�IHHH��G�O�ǯ��L����6ٻR��P����t0��&��������;�����aq.!!!aEC�.�bO�)K��dm��v�T���^W&(��Z�3�v�Ik��=\����ϙ��k�\oR7�����fU1Y��א|�$``oA�+��'-���s��L@h�琈H<tD��hֆi��l���/�6B�P+D�e��!'ZK��t{�<�Y���>�3&\Jy���=�.���븮���ߎo=�%<�}+6�Y��5��¼�"T*�sN����5�q��������&�sE��/t�+>�g��񽯠�U��\%M���<n� ��+*�(H�����n��S�o�����35M2�\��������愄����V�,��6�U���⩟�F4�y��l\���0��`;��o��T�;p���K;'�^�uo�n�I�r��^8O�,Cd5�����P^q:La���U��^��Lx:J��2��}|u"�'��_�`H�/�/Q�o�	ϔE:'�P��*u�\�'J�Q�,dy����r:d��f���/���_¿�����k�{��w~ [�����U�XP�wa|X�ے��$3t��C�p�;Y⊹�����>�/�:\�T:��d����͎���ߡ ?��!X�M��j,���/�Q��#�_?>ƃaޫa%3Ą�����Ȍ,V֛�V���1X�+���	��)G㋛S�ϊm�����|ss�4��1�7���sK�y࠲�s֬
��*�##BJ0�H�Þe^#��C�8�D7����9FRC���f��hO���KF�q١�;S��9�Y�թBr��Հ^@�,˟Q��7S�q=+��\���Fƥ�9�tU�t wyN ����8v�(~p�]ܰv5vm���؆���^�N���}-5��A�M�uk"�kv�)�Ө�Ct3��9�~����7�4e���Uw�.u=!�'����<�E�Z7�v�BNh��
�~��`�J?�w<2
a����}�KHHHH;FW���B�r����#��,A��6qB�ʜ� I߁�6k�-��T��۫��0�)RT��`R:�rg���R}z���0T����Յ�X��l��Hv,l)���>��j��C&��[����兹�:s�����A8L0Hi\}��p ]�n(�V�o���+���3/�Ϟ{[7�Ǘ�n���܉]�܌��)2��
v��4�����tcõ7���^��$n��z<�s'��!�mߤ�Z��X5>w�����"���jm�����Ƞ�>9@6���A��cQÛ>���^�Y��z���C����[BBB�$1���i�g�-�/zf��AB�J��da��$��D���CBBBB�
�W���!B-��4�Ḧ́�{E&P 2���r�Rt�����>�������D��`��g�oF�h;g_�v��&B=&Ǜ�2$��Ί1*�ȸE�E�UV�~��1�s�Q^���{�c�j����F��$7F��\`U+GwnF� {������ŏ�܋[��_�y3��.��z+6\�����Rt��������g�� �Dp2V���#�cӵذ�J���ڳ�ٍ�g��+��q$�)TF���Ͱ=9�^ߡ�}��h��8/���7`l��B6�;i�dk/�u;jc#�A������@���؅z�����A�ŸGSBBB¥Z�T�ޅ���Z�36���#U�a���{%����ʦ��y�H������LU�V�jx�Ή��\!+��*y��&j�Uu��0��P=��'$ӑ�E���%P`��;�u����W�}��t!|��'�<��/�ه�T��e�8�U�<��j,t�/u�7N���_����p��W��m���]wⶍ�cm�kO�2�+�MF��
S�P�!Ŗ�+{v׶����[�ׯ���
咛�{�G�1e��G�ϋ7-�MM�ڽ�L���u�����C��Ŭ�"�1�Ӊ}��z4�cV
^���C��C��a�MHHH�|7�E�ޙ":>)�Fh�Dm�]�X��1��\%'��d�)�I���vZ+B>3A�%���C� ���					=�^��Kfy�w�ڍ�������YֹT��p�,s9C�p�#����pʷ�	Z����)^L&pq�-�I����ì4��Ԓϊߟd,q�G<g��� &�^"��D�3/�[�Y��A����e�l�l�,, 3�g'떢Yݼ|f�`��^}i��ŷ�i�*|m�v<z��ش�^vf��}��ؖ&Xǁ�edY�w�C���r�Z��#+�2'T��O&i<Iv\"p��h�Kjvj�ň�:�7�F@��S�������Q�V�����u��� D��_�HL	 �+n����l�{D�8�VO��7�Hv�	etb�,� ��G�1O���ӌ^��N����ޡ�B�	"�W��6�1�7Pw��;K��ѽ[�}�|:�e� u�(�+����C�:/<W~����@e��>n�PM�S�:�99��I��<����qO�ͯ��?�-��o�Y�<Y��V�v[����G�ƕO�w]w�u��6l��\1��|~[�]��5���Ŷ���b��Jd�?u8�.��|m�G͠��B�j�h�2u_�ސ�-�����5��^~�Ҿ����_���I���w]��qm�g^#x�A�k���B��Kd��-�WR=���u�
��}���1���e���C�q�t�a�+��{���)�5�
�>)Y@ʋ�{�`X������Ke��1��P�w%Z;m$$$$$L�b��]M�����F�B8���� ���*E$$}���;��*���a��sΕ�/���1�鮃�-p#\��ʒ{D^�ܛ�1�����8�3��DvF�����-	��V�!29���<�9�u�%3��U�aWv�n��]1��R�:\�T��܏�u ��]|��-�Ʈ�p�m�aݺuP�Y��u�M�v����v]a�4/�o�Av��_-� eVD�KwWaV�HDE�5?'5)������I1�9��{?L+��O\)]lW��ޯ[A�d!����DL&$$,?�ʥ?2��4'1(Ҕ{� oXM���@�CnG�Tk����S�!.z�2Й�:��DuuYz�B8�����]�B�;n�r]�_Oc4^���<^�i:�OH�KOV U}���P�#\\�����|kV�N{	ko[��|_����N�Tx���:����Yt��.H<w�^��ϱ��gp��9|k�N<�s�l܄U3m�[=��{��V��Yn�Q��O�L���vV�ͺ8�t|��Z�<�n�ꁾ�$]���
ߎ����f3X��R�8�V.�<�:��|��� �H			�F̝����˧K3���;q8���+Q���LU�T��'��f2��t%$$$$��E���3�[��
PТ�R,܍
ɸ�i��ڮ�jK�l�������C"^���b��b�N�ZV�{���5%�3�)g�Q3f%�ˈ��+4��:��]C`�#� �|�ݟҵ##٬ǌL�&���L�!2�ke��E������ً�q����u�M���m��曰�+�:�u�h��Ϙ�j:܊�71��*#S�s�=�>���!<����{�ns��:d�'97YӝqOU���4��,Fy��bG+L�{c�K��Q��/=��~�TH�~F>?��KBB��{1`��G[ �s��;��|C�qH��I�1,P_B�)7.�zM��Ixzݿ�a��w?�A�{E�\�7_)�hͮ� �?^��[��|T*�x��g�V����u�!K\���������	��O[���d��1T�ܨm�P�߿U&��3�B��~X&~���x�~��?|;6o�C�n��۷b��aݪ5��B�+K�HdRRbKV���׆��B7��^{:�屙�a�.c�6g.��Û����v�YwD�|�"�˦�o�n��� �D�u�1e[�<���9[Ng��1g�$��9�pԷ��̙N����n3���$2%@�O��f'4�"��W26��k���J}�̗���0a�u�|NԼ�GA��P�͗�C{C�O��^k��'e�/BeiɌ:B��6mmii2��W�/D8I7��K}I�x���	ϻz<�_�{V�<>�n�"�(ί�x��0�"'1`l��*��h�XD�N�c�7��4��S�2ψ��0uQOM77���:~�+��ⵗ��_��:���޲	ߺ��i3�\�-e̡\��QeXW~�pe!��8q���?�'�2�\[�T%�V;�0&(�^�̋-u���~��C�����}7�p���k�ol�t�R,~B�R�k�0����[�]8�_uW��X�y��^�3�U�=�V0��G>A�8?�S�����Lѣ.-Fy:9V����_��R��=p����=��D������V��/��`#�mw/5;��h4�^W]��(ԥ�e8��)O���t��ezw.��]I&�c�Ǩ�z,�}��I�C\6>*>W�uX�u������'3a?�s�=vX"����[�13��ay��c�����`���`�u��������w����f�*���v���Ima�8���{m/���!gf���Sy�B��p�f���{�W��.=�j�sN�o��4M�ZQ����˼��oA4��	�FiBL��I4����ݴ������V��c<cԨ�5�k�����^k����Uc<5�*I;�����bQ�^���8T]O�W��>k�q$�i�q��+�ڎ�?��)CI��~Fpbbb�}�����|�rvGG�h���4��8!|�pt��o�8l�ᩓ�"yk��&�i�Gvʵ"�u�R��R��A�S�B������V�����`���LQ�D����ϳ�tA�V������~�b�˄�d����RP"�iM+J�<_�!�ggk�~F$b�a^x�H������z�>_�HV�ˠ�^�O��K7��F��K<K����^����\[ro��v��jH�?��?�Ӑ~��	~�~~��F�O��_����ܟ�3������v2ǟ����v����뿔O���5��%����A����?����[�q���.�Ϲ=
�.�@s��[�[60j>�T�r�ԐI)��ㄭ���(>����Z����'qG�v&x[�Xr�`Ҏ�D�ث�1�~bbb�8h����W�gQ���)��pyj$��?��76���(�'����+ޒ;YT���l�Ë�r%�VW�MBj�F�L����+R��&kW}ߊb������rmp�W��N��.���ڭ�&��/[4�R��I}|ಮ7me�YEoH���z���j=p�Y�K�}��������w?����������ʯ�������_�������v�������_���wKљ���� ��ȗ���5�����z���~7�����n�|����cD��o�C$�[�MQ�Q�t���ӫ�KrwK��RތX��;�����׃�^t�Ж��Qbl�;�l#'MEz������?�-711�QA��
�k��K�Yg��ms�"�s�!��/A�"��L��׻�7R��Y���(<�;�D�S��nq�]��48�TDڦm�[��1�9�OLLL�����]�?��䪮�=\�ce�g����9���^ex!�r�yvK��>i�^���g�	���U�`�~�������]�R��`�=�ģK��:����t#����J�[MH��L+�����]I͘	�oq���[����w����]��ׇ�����������9���_���χ�O�r����4|[w������_�_�=�o��÷��\&r�h���ldA��:)E�N���9L�m��Kt���1�g@oܱbW��O�o�JOLLLL<�l�S��S�R
w�C�!��`��|�E>=���7s�I�b�I�e�Wq�`�����@�;*��Y�>=��Y��@|��Atb�R�&��2R�6z�g�2����h	>�%��E����U�)u�.�d���|����Qni�R��W�g}���O��������~���_�_���m�7��_�ο��ÿ��t�S���C���Q�Ϳ�����_�o�����:��'߇�|�N��ƜHyյC�!���/��U�.�<���U�����e�g��C#�TN�t�����qFZ'A������J���$� �����
ԉl��w�	���e�f�}a��#��'���'&&&&� b���	+����.N��ĺ���ȩ@�Ò7\p7�9��`Y)7{��	��f�X��F�w�C��l��W�h�v<i�y2_K���U��Y5���Ae�3Aӯ���[�-K����z���}/��n?����~�����~�/��?���c��_�'¯��/����8������������~��}�	�K9�%�;T�ㄽ�W;�jO�֢��o����"w�xET_�[�M��Sw)^i��:�+u����p�.�:6���Rz?F1R�aa]���xڔ@���ldR�b�A�����j�{�ڜ=��L�:}ݍ��R�Ŷ奴/��ĺ3v3r훷W�g[hYk����}��K���s��|�k�������~�!�s��/���������7���}�1�?�C�nՓ�©�Suٍ�w1B��)��8�bJ��$O<����̗�K��9�MLL|U\q�_'�o4��s�RNf�a�G���u����7�8"��@8}䬍G�@�O��c��211񕱑e�=	D~��G�����
Y���Z��I�Ս+�E�_EJYNO�fo������q[�u*��J�G+e�ŉ���0��1*-r}[<��.�p�����Nơ�(OL���������I�����S��f�m�����o�������'�~����-��'?��?�mA^�-e��*Pc��%1����3ްש����K�:D��Ѳ��X� 2rܹw�=��O䙘����LH��E�9�ȵ]Gq)���L�X�ig�Ȃpv��P��9F��#���+4r�/�3�(�eP jS1�PF�%�3q�})q(���m .��b���>B��!)��u,+K��%a���>(�[}��z�k�+���s��s�e������\^����7]�Uz���k�_��^B��oK��������K���/?|^^^?_��j�/e� ��!�� �Ac	WH�mu?1�}M���s�ң=��[j����GG���M� ����Z#�[f�cqf���x[�Dw�����i�j%�����G\����[8��7���Y���G�u�l�"(�?!�G��;����O:�Ήbb����x0$`�L�>�*�G�9L
���]ݏ2����F�:��d�ӗ��� �¿	Z�d�K\"p�a�Po�W�s�"}�FK�Gc�@��^�R��Ek��/�����	��:�"	Q�F�"���7y7\.����'	���m���_�o�������/?�S6b>ec��,�ؿ�3n�z,�GNsN�%rުݮ��-�����+�(�� ���.\O>��;���	�q�;Br4Mܡ�c�����9�}E|^����gA��|�/3xȼ�sPWnN(I�E�����:3����O�|U��r��a�4��QG������ڴ,�Ӣ��ʛ��Z&IZu�O�'ph���������U�Ĭ��h���ZB('~���~4��jfu����@ۈ���1d0)|��	����]��1�(k)G�g����6��'��Z�l׳lgx��Մcӝr߉�� g�x�qIųQ��
��5�t���ї,�_k�v���W���.�KCj`H�R~d�!���Y�i'K�<f�OLL<o|(�}���2�ܲ�:���v@���G ׌Y�&�����d��a�[R�,�\���x�>�Z=111q��8�BD��V��I�2��5@b�iR������sEB�k����8�iI�#a�ء�mp��9~��a�B���~��d�Qچ�W;�L��O[1��ރ.���ޏ�~I���P�r�N��谑�1/��J��v���>[6�12Ju�'>�
,df'�����=r�<��u�Q�2��8o�y=�	�V�X��k��-Ќ��Q�E�������e������7���NLL<5h'�ʝZ��@3^��4�-_�q;D(
���/7�	ї?�r'p�� 3�H<��zUP�I�����$i�	b�����zu�����Xv�~u��I8�O�8����|zFx��u%��N���d|��y+�51f����u��_O$\^r�[B1� �7Xk�������T�Eo垈c�#��JV��{ơt���@��>�g���pq��"�8K2\�:N75�n;� �� x+��NQiqO��W_�sbbbb#F���24�v)�C�'U߆�'�'�u�.3K>pG�a`�}�R�D�c-5/a/�ʀ#���z.e�]���Ņ{P���&&&&&>�N��Rz4�p��glP�9#�]�j	�D���D^�=�U�D�D�7/bgG�6����D7�*KL�Er~kҒMR��,�4E_�G��a`��@I���KB54ɱf��z@a;'��H+� ���v�I�Q,'�-�����WJa{T�O�H�@�XO؝��`�f=�0�P�S���Q;�G�]��FJ/�e���Y`cy??�#�0��g�MLL�%.�7���u���͏`��zȓ�u^M�6w����c0��A��C��'�E/
ʏʈ2��B�M
���5ҫ��,G��ѣݽz�R��A��\����O�|G����;�� ���׳G�K����/��f��c�Ƅ����g۲P�$��Hy�t�v�tg�PQ�[s�x�R��a8'�@�279i����0�b��>
��������]�����Ɛ�S/�*�s7�-Ze�'������8�@��79�!��;I�$!��m11111q/<©��L�m_,(9���hs�\�	���݄'ϛb�`�7H��̧/�E� 귵2�6��9b�O���B��Q�G6���~ğȓ�v��R��J)��-�-˹��^o�ꛐsT5T�Z����m9�0��e��"�#m%�YP/�[�.J�z��7`���c1���_�$�$��D�Z��x#��ZӾ���<	��V�ۣ-���z�^���;1111�8tǁ�=oH����(�kWǹ�]����Af��Q>����{ �u{
n4@���Ė���A��Ȓ&���K��ڮk�MPuֺ��Ӱn��SO����8��F�q)h12����Y��^�T�N�.u��n�aA���)�\μ+��̞i�q�j.�;:���m�=��5�xW����L��gy�Zʉ����~��N�y�깉����311�pt�$,�Z�l|����i��o����x�� 9�������ϭJO^!��T�Nó�����_��'�eebbb��Ox��j�BU]:+a��C�zW�N��Z�ҞA�w
�ݻ���׋���B5�@��H�O�mUH[�/����z���������6I�m,���1�f��k�b?-~�N���FF�oUjPZ�g��?�#�'��3��O��j��"�������m�4	��,�����O�~<һ�:��9�ү/^�8ߕ�#���
��*�5A���5��:N���������%�9l��9��e�Ҧ����?:b� ?_�T)�xţUX��w��	%��;���~GH��eW�e��A�Z$u�4?��Y���1Cɔ+[�E���^>D�"��.0*����Q�ߢ�C�Dǳ�D��ms�;���;Jx�4���JDPQ���Ŀ��<c>Ч�.]��	#�|��W�ӯ�<-~9u5�W���t]�{�/y������=����y��C�Mmow��v����M�XD�Il|�~�>��c"cfR�Vv���&/؈U�c��jqk=���~��<�?@����DY�bx�R��&����(�\���������
�}s��_^$w�ߊod����<O;^��M��	�B����Żl��&�e�jぜK��2�s0�G����Ts�2h��"5-i��pE�b���bY7���!���ĥ�'0�0�I�!���1�A_�"e��Bh�^]1c�Ws�l*��ָ���F�+�/�?��t��Т�G���v���;к����87�q[���Ao[/ǁs�?7��Nmۼ�1��V[4߄�\Bo�;Y��#�+TXd�%r���A��a;��Qܔ~@�͢G*�o v�����vy���=0�lO�#�x�U����:��v�u��~��ݎ�g���5"��G����ˉ�=g�n��R/Z�gɐ��^9U��.��9�*:�������x�6�Mt��%c�,s/4v%ۂ�������K�m\��n���jޛ�xۚ"�����(������τ{Ɓ<��Y�NQ~�1���T85�[�z=�2_恻5��-X!�o� C�l���8�2�#�J�KK�d�K�&��|�}�ʇ�d���^V�rz�	9����������#ߗ�(��c�3�E�tP����D���(�SJ0�F����>$�����4 ����JDk��7zT�ƍ�8��#21�qǏ�:ϰ4*����i�U� ����$����?yJ)�C�z��� �zBc˪Rj��Q�A����}bp-�l��hm�\�ee��!v~MLLLL|�W�E�Ѹ$��c5�{��G��?�84��:��Ax���� b�����Q�L���0���z���c�FW�:���cq�%o�rk)��4^XV��!>�qm���١��8��G�/�+,Q��Hq�F���]�isNy�XG	-D������V���f��A���Q����E^���'�$0T�;��;kdu^�������1111qd��2�f*��R���䝦}0uH�Ɠ�Xz\�@s�'��1#��t4B��
�9�{��11111���*������l88w|^�A����vn��
%G����J�x�����9C��XӉp��&����%4�܄�woh�A_*�U��2a���|�����HS@�
$�3͓���ԐƁ�V�:F�6�}�������a�(W���4�Ԍ� ���ʀ;�&&&&&&&>7b����C6ޒ�Ӳh�h;G���H�)Ѳg�C-z����Hf��9�Pg��mT�fٻd�Ix[+���c�X�sr����i��AUG�q۰�Z:(~xR	�tQ-0���JW�>��{2�����Kc��?�2���п�M�O��c����nm�!�?��ˡ��]$��,k-!��p4��j���2w����xhΪ�7Y����&<&�-�v ǽeo�&����!�|�q�	�*D��~QR�U͜�'&&&���Н����P��`�V;m��q5�Q+�D�!a�B��>�i��Y/�CV)�����}��[&�K �-�[��rU��?�ړ��XT;�@�qF(QMH6�8��h�|$S(�y���cU�R0/~�>�fߚ`�w��"��"��>>�&[���c��5&�&:���?qs�KD_��;V:;�M�`��Q��gX@]�G��M�7@>{e\-��A�[�)�Dk�A��j��3�����+��,7:�]�o�<��v���N��J�Ϝd��σ'C����>��'jV����^Q��b���bD,R'����s$�Q���p�d��W�N��&3��=�pO1�:ʕ��/��D�d�x�b�T�I�o�>��=h$lRig�y~�|2{���ׄ�u/�/e5���x���qM�u��v�Jzq�{�x�}@_�I��}|�p	M���J�{�b�6���'&&&<�����TB�D�����#�8���/�f��Ѯ3&/Q�����]�)��.�X"��Ey)��܁?o�Eb"����g�Њ��M�V�s��0.{��o�^��0Όr�W��R�{A�Sa�!�����*#ړ��`��%�K�F-��)#�b��œT7`�{[�5�s ���\0�*e�}��8�c+˯��)0��/��o7$�ղϗ�����w�h�,���7#�%{s\��u���H�NC��'��{���?$ݽ(��C�,�F9M�� w)1�DdЋ��<K:��]��g��Z��n��|Ib%���J	��S���f�"zj�k����8_��s���մD�#�S��CzL�F��*F9��-U��x��A�)�)�7����Ɠ��u�\���px�'h��6��w�^�,��7�Ƚ)1��;,J���
Z�nq�������,G�={����F<�<�*�b���c陹߻J�Z����y&�_m�d���"��Q��=�^���G�� ���DQfd��������ϷW_'&&&>��N���&K�ܓ��x ���,}�E����ju�>�t�;��v�L�2�YB8��n�*��b��BП��u��o"�ܾ'm�3|j����"�vߍ�$�#�ZELB�I��y`�Eg�ˋ])ҳ(��GL�E�Deȡw�H���c�3ρ�w~{y+�������lw-|ݣH�ۣ��ڿwD�o]>4��R����ym7����3111�� �������n��va�n/av�Ie13߅����s	5��v����i�O�Enl�I��9u��eN0�Pr���I�ULqɷ���J�J��Xj6�8n���5�̦Qk VnWژ<q]�c:�y԰�����Ʉ��B}*�|���m�NCJ����F��
P�L�Ӿ�#y���Q�.kF��]C�I%A����BgU�Ϣ�/�ҞX��/z�:N%�"'P���ٽ���`oQ:X\�C�>K��?hnE^/�]�ώ�Ż|qbbb�,�Ɂ�c�$�T�EM�{<�=��Fp\oIa:�XD=��z3l�O���ȼ��5l��� d����/uG�R��	gx��ؓ21'艉�	��
zb�WX�8@dL���`�vt�*<<����w���gBh	S�&��Kz;oHҖ��T�F�t^p����t8Ek�_ӥuj�a[[�v�����o⿭xc�!��G�+B��x:�C�p�]fB-qW�����צEX!9�|�'�{����#�L�OLLLL| ����bh�9-��O.k�m�lA#��}���x��G��	�����9��Aތ!:��p"}(`���s���:�P!v�R㹃�(�5��CQ�a�s4�fN<-��;��|Nm]W�3)`I�,3��(\��E���#��-�dL���:;��bO�Pm?W��U�ߣ ��U���P��b��җ�vct�Ջ�-�8��y>�������,s]��p��^�W[�N�i�{Z�M;n��j�UeL��s�w>&|�W���̂�cO�������ą8�K)b&�B���x>x�39m� NS�Q>Ч�=�wY1"��{��4m~���*�Vhf�@x<XD}���^��Tџ�]��ci ��g+�VY\�r/��Y���`	�t[���I+I:���$?MGm��F��v��P\s��������g�*Xh�I-6�7�4�[84q�]�!���v��m�s^~7$--"9^�?�Z��f�P#,zE*�]�|}���5�w�t�v^o���<x
��`��і�E�-ݧ�@��O���PS�C��#����Rq���1�h#n;`�j$]�E��0VO~��mѮi�m��8 �������(Ӎg$����Bo��zH'��#Vc<�Q�YR���;LLL|e�&�0�uo�����0�����r��ד�[;��$�>�6��NL�{+\wp<�p�[��(���>�C��Ԕ=bbbb���0^-��y�v�Y<�_c4�n���2ޡi�1�U�["j�'�X��ɰ}�IM&�JS"�;�ns�T!u�LmD�%H��i��T�;M�gR�N�kK�Gtz��:*�t�Ub(��o��HfuȔv�����k�ז�KUA�WI��t�!{&�w]��{�>��g�'&&&��]�YYL��4� �Q�>_��G��1�Lk�
2
rU�Fn>��zP��bn'��ڃvM_�&U?�0���d��9/³Kp���QQ68�%���ǥ���j��\܄�y(ŨS�Ng0ѴBm[���ӏ�Y]�ϣɓ��<���P���'��R?���X�蓥=��'[S�����\�$�M��+O�x�S�>"��P{��#χ8OR+�$��������dO7�$4��*�j����+�X�μ�Ʉ�ԋ'&>/|�fl[ݖ�$�$��V���:�c��kI&{~G�
���oJ ���%���yr١�\(���2p��9���J�̷�P'��p�r��6��7�Y9��'�
�S|������
�2rd�p�A"A��<��9��PĐ�y)~��}O�����o��j�K	h@<���\��9�CC�O�&^~DN�z�pًO��߭�ٵX�7�Ǆ}�Gf�Ƨ��xߝlW��7�8�g�m��y�,�����L��!� Y[��O�s)��!U4h{U�D�=����q�O�F����9m%�K����$��0�������G���S[7��^J�Ev r�^,��g�3m˪�`���Bn�;�]iۣ����2��(�ϲ�5�-��^�&Po%���������)?M	�X��"L,�섔.-�����{��l>���1�y�����ӼZ������oT��2������:/��� k����=�<��l�<�ڒ��=�N����~n��HQ�)Ct�/b��ɸ��ȼH�ً'Ϗ�ܷW��'FGE�,MT�pf��F��%�J_�+c]d^@�<4l/��O}��n�����%,�gK{g�g�7'&&4ԛ��KMtn�p�ԓN���1�F9ݖО�)o�ׂ�IMj>��'�6��nk���]�^��bڀ��-��8m��G�\�6���<}�8����s����(\���_Cp�����(X��u�u�����Q	@�H�P�M�%ZHF�m�]*Q`p��-N~�E���Z ��|w!�E4�*aя�J���&%K:�g��l�(�[����o��l�iq����5��R�A��wAc��&����}ؐ�J�G��s�v1?����O�4��(_1\����34zܜ���X9����H���8�&rjS�:\uN��T
��mATI�Ɗ��&����;7>�#1�A�<�/jbF{�}�*�>LY�d=u[��s���*��<�q8Y�֊���_Պc��tOP�ԩ��vi��]��<�]��T��ZS����=kC�u����D����1{ȎB�+2��&�9�Q��O�p�~K���H��:��dP�����6���� �`��y�-N�����HA�G�~��p�.s��<�q�e��5$}F�X�)����t���H��'#�F��?m����غ��Rz���&7;q&�;MLLLL�'V��t�S<��uΑ�)��Qf3�⹾ӹ,����Vd7H,�!mZ��Y��,	Ȃ�a��N�Z��Exn}�۔��G������#'��U��	������2iyd	��Äs.p4 Οo�>V�r	el��ɩ�=Y39�ύAX�[�l?Hgc~NL�jbbbb⣃�0���F�mBײU�g"�=M&���q����b����S�_���tXY����YbIN˚$��}�'�V��|&+}����~c��6��-�K�������/�WHAI��Y�A�k��C+On��T=C]�7L�T�'{P�Q��%���s�������1��;�S�e����hbpv4���K<���M���mx�N`���d���7hqqbb�s�A��G�8�⎴�U�3��I���#�^���.�I���};�"�ܐ��ė2�X'��������cZ��jT�nߦ49111�ިɖ$B��%�[aU'p�S�
P;��n4�(��(1.��l���-��&$T��9�ެo)?�������x׻�B@��ec�^��ݒ�-"�g�a����p�X��9״-@�[��b���/���7�ԢɩG��ڬS��Ŀ��Lb��>e�����9������g���=�{���q�(����Fz޶�����"W�E��'�:���%؉�M$!9ey6�XK2OyºH ]'�,Xҳ�:���nWP'%"S�9��㲺��*ٶ���s8�ʈ=-�BU{��5A��Yj��x��Uջy�q%p�n]@�Q-a���N��*3����>���ꮼ���+��e��q����'�}
��F�򇬠�X#�q���.a�T��/ԏ��{Q��G�6X�t������}�H����8�;6�ް���{��Pv�e�cÞ��*Y�n8u�s�7[����#�#�g�I>bHj� _YBmd�J�sL>�O�2�������8l���+��!����&�[85��T�ʖ��D������ ��6!DD�6;��\/��pg��y-> �GO]?f�W�(�Ju����~8�I�v�8�O��5��4��aLv	�>k�Q|����]k� :=B�#'���yi�����]!�-�œ:�y�1g$U^|�^;����([���XzHN�Ɵ��,Zq>�j�-�U���Hj@�;1?l��Z����ģ��$�#�&�9v�`���0���ax�A	5�$ޞuf�GO���m9��wTۓ�	��m�ɾ��d�����]���џ�C��K��7=��*���߈��u7u��x�l�J��^K��ӭT�%��Q#;�nUc%�Qg���LG���pI*H�5u�p*z���������_1�	�K���r�X��0:��W�@��&_��AIyx��Bc9�K���t^̗ʣ�M�r.�|��ii��|��A���w���t&&����{�rx}x�O��=X�7�Q2�6yQ��m�Q�5ylIF�ak����ȷ��1y]�_?�����/"�z�ו����<�h��/�jճ�=��n2�تm;�B��R�b�}�l�ʔ����}\�vbbb�9�N�+��MH�<���B�R���O���\(�%F�����G|`��8Ǖ���7ftb���*�7B(4�(�+�k	wc�G�ߙ��¿�,�=�HK&W�Ϛbx��I��H#*�ԓ��	�ƫ��µJ��nQ��E���tK���ں~1G���;�h�iѸN� �2��2���$�_�r�joW�Q輰ޑ��������orGc�BU����}#��|7I�s��V['&&&&�n?�7�͙=�Ԃs�3�m{�@�[�����8��=���ߋ�VI���^�d���4�"?��i���C�p�����F)g������+K�3O����M�Ae��,�����ǽlņ����d'�n��s�xZ�N ��N�B(8�@�%O���{Z\?�B��M4�_��z��f{��;+����$}\D��x;�ɾ׽8�ֈ�-iq+�I�N\h��L��;�U_�����>C�qӉ#�d��=%�=��jx;�=Ô�	�=��pW�9�d>�m�7��PƗ�q���~h�Z����(gu�����"{=�oJM��~H;���n*_�
R1Ov�9qMLLL�#�T7��sQ��[<�<ἐ��;+��p�d�E�a���E�-�	e�>��V�Ex�if!+������7 v&9,��d�S�o���(�H��sv6�4S�9Ɯ���{%���%H1//U�p�{�r�q�~A;�<*�+�ͭ�L��`�sn�]�)o���*�{
�#w=#Z�0L��G牉���1x���!O��� ���C��4��Z%Ӓ���%#7��:y���h�s�q1�a9��� ��U���:�3V&O��ݫ�Pj�}��Pn��3/g{D+�=}%9n�<4T7�)jk'κ:�F���P:�n�����4�����I�2����ា�w�{��<�Ũ���UP"K+�Ӓ�y�u���~�Xtnǵ���0T)��Z����}<��Co��V���O6g#�%��b��8�`�P�hW>�a�5��J���]_ȀCl�c|���O��ԡ&&&&>3��[���s��*RS�Yd6�,����}�=QS^��+�¿xk�A*���&���	c��`*?�cH憎39�EHR4%hQ|���-�Y��u�#�Kj|Z��q#w����0|�&w��/���_xd��@�R]_���M��/>J���.}~��$�T,����G��2111��=�)����c�=��w+WU�=�#�w�o�B��,i������U�Yj'(Y�������x��Δ��y*��yЅr���M?�9�Gx�'Orx�Z4��1z8�������G��p-�I=O~-�JaJn_�HO#%�h;�����B���*��1�	�t�	ċ�.�����6�b���ꓳq'&&��X�޲������0P5���L�����|_!ۻW�P�<��N9�C�GHWxxg�W	`��=,T�^����n^��;_�֞���xnl$�z�e�G/���s��Rf� �E����i��L�yX)&�V��N���L@D3.�*s-��,;G�kR���;�S�c�d �Xڈ��٭Ф���[�YA�06�w A\�#��3��ns�=�v�E�݆�4w�L�xQF�mg^F����{G���c|�G#�#����r�ǏAz'������)�Պ�{�h)o;��c�t�'«��\:�7&&&>"���͈�,���=��^A����K�_���X�BD��q�XhѶ+O�ZD.>���yK�*9J7OE�Y��Q�2Z�����ȍ�sҢ{�"�)���:O-��:����	��'�ȁ'��@���RE1
P�����ian��U�9n��1�-�Zܰ]�ڨ�a��z�\�0���z�uVeՄ=3V�S�`�w���oQ���E)�K�@�Ǿuw2���M�s�X{����1����ѽ��h^w���Mkb�A�*��yfϐ�^��Ǯ����(�=���xC�{�N�b#��Ѧ�l�"�hB��vq��gK�t�LV,�H~�9�-��p`�� �ٯIJ�vA�_e�;��y#�q?��}�8_D��ؘ�c�u���c��
JF!9���?
@g�LZ�@C�^+�
��i��3(3m�4ىHLxJDBl7�R�G[
���>zX�hJd#�"�����"��fH�R��<�͐�6�V��VNu�1lp>S���&!BSB$��9H(.��W��-K��n�A%1<�����)��؈ϋG꿧�U���.���i4����|Ģˑ+a�w摺޺�z5@|ɳI��ޱ*��.��;��O�Xn�R���c�z�G�#�1�F��A}������٘��W�BY����F�`�c���eo}]�[�#�%�N�H !<�r5��o>Q_C��wB	O�o`����1�"_�<��Z�J��߈p��ۺOU[������t�C�Z�Y+HO�Q���4V�3YQ���BEVLР���P7��L�u�\~�S�t�Ԉk �TI�AE}�QW�C��s�wM���y�x�Θ|6�~�*��=�7�C�lБ��G�|K��e^+�YU���:ŵo�&�[
8��}��,w�ݕ�'��X�#��Uz��ǋw����G~�zv��1�l�Q�[2"X�7��"��Bک��;�d�=,��)�6/(�o�����o)ܾ_S��5r,`��'�����C��R=�Q�0J�:b�2���9��u�-��v��W��+����*4�GIXdPB�9�#���3�//NLLL܏u2_��W����;�Q?��|�E� ܱ1���6(O��Z�;���WB��d�d�T�H� ��Aq$ݤ��	�4��o�ԋ���-��(>�?�¸Y���d4�*Z�|�(�� iX�y�v�Q��R�7�~U�%���7�I��+I7�U��,X2�'l��d��a�o�U�8X���8u��݉zy�GC���3ekbbb�<.��\�d��H�Vҳ�ɡ�p�������_���!,��,�G�Y��`���w4B��	����c�v9ݲ8����U�ݸ\j��%��D��'�D��L���ֳ�y6�B�`hӍ6F�j�gu/���wO���H֯�6@ǘ�*"EB"��G����c�Uert�^���{\�ꅸ���x����ٸ���e[�:x�����4[̲~�8���ꔒ���K;��k�MS���ƍ�n:1/���M���qҭ����1�?��{�ݼoR����[��	�3(P�a���쥅�&d�@�V�K�3��0q~{��O�3���ϋ�zV��I�q�dI:�<��jJ&7h,a�/��G�}��$Y�m�o��8�+�5Y�{`��h���8��3�|Ns��,�دO"���s�4@�k�lG�(١">YvI��H%C$Ṕ��x�SZ$�X�I���\'^�����{=�E�a�H�p��G�9��u�1!�&�s��7ē�Z�f~i����]=���~[u��lE�:�W�P�v��ү��>?�:qսr���[����щ�UB�a�,=w��2�;=�[)�MK.�5����b�\2� �d��hF�ע���ƅ��c*�r�tD�,�V'p�ɧ͎HH-���g�.X��=ݧ�BO�Ba�ɂ�s��A  ��IDATn�Pk`6'=}��Ӫ�,a�x`0�Ս�\�ܷJ����Ѫ���6&�g.|G��v���kc��dx����/磪`��6�!��C�T��2�E����Eu�;[`n��������n�9��4
ۗ=?��g$�+��wL�Y�UP���ƗczGl|�G//� B�!��)MKt�-{<����ͮhS�quʀ#6�!˗��@ɚ}�{J�A�p�5��X׫F+^OAtbb⣡?Ɏ��yN����<��u�s��/�<|���[-Yr���e�*6$$~�Xv�g��Ӏٍ�X�DJ��I�7��%&��3�����	�P�П�ӎ��j��1q���*spO∍�R��~�Y�/��L���W��c��Kq�#���mݖg�6]#z�+�X%��]|u�\|�`�����h����P�R�� ��N��y�������������Hy0m�}�y��T_�^^^ʼ���qt�"�}�{�������O4�l��ў/�,®�[�LD��I�!��=���VQ�eO6JP��r����tk�c'�U\�Ɖ��*���}<��>F�[`3+d6�"ѡnP-���ij�Hu�V:c`q[�(�'��>�W���<��8�hpy*P��I=��H�A~�A���%m#K$�Ǵ���<�;w��d�p�{o�箞9u��_d�Q���R�9)bs��]ם<��ז�sπB�(,c�)����A�Z��h��G[
�7��7�0�j�µ[��S�2�"($�b-�ɣ��xqV�������o�����Q�����%�v'�x�mĬ��s��W����^g�#���TK��1�f���B���LJ�_ͳ��I�<��Y��<�u~��۱t���줞%�U�=�-8��s�$i�r��c?l�f0���́G��H>�kHWD���Z�h��yj������8��Q�Wu{`H���؏���[�*��(h��6���Jh�q~��}P�䁭txy�$�7着vbbb�#�e�󃚷�l�t�?Gc�{��5���<unIS��7Vc�9�{l1M�V|O�~��G�k]"?l'!���J>��,
F���m��	G~��<*? OZ�����G��Z���iCvy�&F�l�)�����<�X�ɹ��������t [Z�V�,4�U'q@ƽ��Ey���õ�@}�u��p����}���ҤG?�R�>�3��y���%5���$���cֺx���'B�l�v�a{'�h��[)�G�0��w[֯�s&&&�"�1pE6~��faN�x/��U�������v��l_��p�1����E���H��i���)Yh�☾q��Y����4p̀#}o>��t�����Tsæ�P��N�j{"'�%unʃ|��{Om������'P���RQ�$㺔n��6 �?*2i�$�.��G@��G`k!�p�s�v�f�QMa�BIy���Di���0<ZÒpe�z^4�.jc��ΒGʅ���������Ǽ�P{N�\2.���: /I$0Mr��$/5� XƉ�3֎^`���VB���E�����lSZ`��ncuKf�)�z'oȵDwT�5�T���&v��t��h�)����%���(�{�-�N���y��������:�ş��Z�~�����G�d�1�T�	 E�o�)��o8y} ���E��|$י,����v��繱~��%S��|R���5b	B�wts-0��x�Ή�����h�.Q�b3����N��C��d��䔢��i-�SJu�$~���ړ��t����D��OO�W��t���fs�g5�vQʁ�(;e�����zE��Wv��6'���vc
ד0;���~Ku��a3��b�W2�HK.w1����Qq���_\��ꓻ�Z����v��%Q�R�Srԟ=����2����A��!�x�
�x�������>�����r���75����0�n�,��[��+������^�l��K����H����h�#�w5'�qQ�YT^�~+�����
�׶.���t��c�`�1
� ^.y�.��VM��Oሠ8���(�a
�̣��:���"|$��ₑ1ᷔ�� ��̛\���(;_�@2'�,��Ю� ��JH`ub9 U�J�ʍ�/ܦ�8����"��d�"�E�+ߣʷu��G��i��I�%2��ܺa��5�PV��HX���B��6�[w�\ޕ���{�,�W���,�I�� �O]#�8r��}v��[���/��5蝵c�����G¶6$��Z���~ވ\�z	-ɮ���_c����!ёφ�X��5ۜY�MA�N{�3G�y�-�c�M�7,�Hbk�'�������S"=#�������� A�d�j��£�c�Vt4���k_����sVxnӱ�;��`�3�8J2�'b\	©7ۨj����f���ad*�d��p�NC�]*'�'����vђ��E��Xø�ҷ�ZȔS����=NT/��]�;�}\c�R"�F���4�:OT��vm썬{��+��1�A�2��~9S	�+37I���-���A���:^��,��%�e�����P�
EوD&���$A�}>ubbb�ˢ��,Єr�R
��+����������EvvAS	q�P�L�"7� H<�"�prRK��P�E�7%4V_"�!Y����3j��7��E�T�dRD�g�����VV��-��%�$�M�d]/w�C$�SЎ�d��U������[����-R� <��H�$����Ѹ�r�,V���pOZog�����{|��ۯ����111�A2%�Ǽ�|�Qs���N��rA>q��������ϾW�g�+U�������#�?��u�����H�m�XPgbop�����LI�E��:�7����'*���0�&8*(��4v���x�[��F�������$����!�Us�aHn�&�f3�D�ȿ.��v�)���l���@G�ϖ����0g�z�v�����q���@=�k@`wh',�V�������6��N�hF���\9C�\e�1
4ЯO�m˴-|(��+h�
}w4��#�)|LLL|�����KGT���˲l�ፏd�o���5�r�����`7���$���5(���Bg�8���g��m�JR�9YB�?!]"�Ʌ �ʖJ�:�@g��DJQ��&Y�@$%��j��c��lϭExZRo'i'����PS�`�$��!ɧM>�32��j�{e�k�s�W��K&F�G��,s�Π��R>:��Ɓ�<�b�U�%�xXއ�M��Ӈ����%��&&&&>R�c���nP�<���7^�����Y E�d����S����a�?�}
�X�ݝ�G��EZ{I�Hj�y��S�#��^�n9.������������u�5�M�)iFK���WO�M�E����sT/j�,��n$�:Q��B�7��|_ieF=�^�=��=O��~���c��D(��c�x�R�o���v�<o��<�8M�p��vVpKU�~�Q�8N��"�_���G�r�L�.vFׯ�^��4������5l�����}�Np;@�񒝗��Dm ��w*���K����q��x�˴�� � �n���/r��L{���d������ջie�p$�����%������=Q�4��� �׹j�+�2������b,i�	,�$-����B��&�"QN��.Y@J(d�����&���p��;���,�n�!���W�Z�J}�l�U��Tx� ��e�[�=�LЎ8�����A�9R i@jB���d��R�+L9q^��@m�Cr�qL��$����Xӣ�zu;��"=`1�s�ջ�Qyn��n��t����к�s}��~����f�t0�{���n���n�<tj�.�v's*c�(���﷗�g?�j[&��h��6�)�۰כ�4�ۖ'~/�=o������ &�%���eo�2G!�ne�]�^,z��6�$�1Ӟhwd)����|���ܲ���Б�A�)�"3է����8����e��:n��?I���x+q�P����s����:��DV�j�eyʨn%��>��G��z�B���:a@^*�'��a����ˋ:��>����"��5���y�/����*�V]����>��b룕�A�wK�4����	��$�Uh���S���l9�4�n��j's����Ԝ�H=ʵL��dJ��2�%�9V��N	�n^�P��*���{Z}/��g׉���+����/3W�a0Kd������H������ʣ�46UZ^�=�\�:��6��S'p(e����}�V����˒ڳ�?0�^Y�q�����ėj@�x�gT�0��������	\T��Q!\�U/���E�!��-�2 d�
�D&��1J�I	&r�5FCτ�IHL�ɻ!Ak$�&:�3K��g�Z���F�TJ����#���N���/�������-A���ޫR�~�
�}�z��n��ۭx��o�C��M�G����^������穉���.:����bE�@R�}#����ՙ9���Y&nK�WÓ)�.�mp�,�z��#SBcm�<l��N��n�o��<�� n��~�?:R+�$ѝ"<�r	���D��|�"9.���2xZ��lO���e,�a{q'��y��cTqSI�ȀtM��c�c���b�mY��H�Z�>��r��C93A�Q�3rgk��W?����)=:�F���2���2�Q�:܄ɐ!e}һn,Iڤ�$�3��7�;p>R��)�5o{6��Hsbbb�~����U��d���������V R�C���Q�6�^�^�Ҧ��y�*尖7�$v΀#R�����)Pv�2��ǥLLLLLL��(��h��� ��9]"����* =� d~+��%o?ܪI~���]���MR�کV<nqq!oI�BQ�e*",���	��������b�C�z�X�^��,�����k�ۨ�$p�l��{�+0���ٻ[����>/�^F�u�=�����-�;�x��u3�]1�|��:9fbbbb�M�,q;9dCZw���˃e1~�vN�J@�dy(_]}%jO�E��ǝ�(Kl�K��K��t8��FQ����`�*3���#����3�ɖ�VLm���p�~��N+�>\C�H��lZ9���y���=�p?�j'�6U�Γ�s�q�L\���e�gk�E�&��������A1�n�5�w�8��yt�o�����Sq�S��c�w"��!sd��{�x�9MKp鴍���i�gpʀ�U�%�"!�Ȃ-O���dbs��|�➔��&&&>�m�cn?��$�Vo��c�H�~C�{teRyH�|F�%IJ!�Na��%E�Ù7����h�.���b�HKɌ ���)aǒ� �)�D��c� ǀ��6���dL���[iWTsx����B���w�������ى	m7��yCuM��룈�g��ҝJR+-��x���]�4^����5+�mOn���0$؝	�!7{���䚀��-�"�I���1��4�Q����1��Ǡ�۩#��_�Pig8��~�����kG�$�02�`��5b�H� >Χ>U��W�g��p���Ρ� �h��süւ3���L��<��7�N�O�b�n�~��bb��t�����hU���C��1|�͢	�}��z�M�&�.���g���I}���ٷi�������Ó��L�VYXo�\n	D�$�|5��Jg�����UeY�Ӧ�};�)�剎�ʵ�PjdM��pN�ꇈʃ�wR�;}zے�W��6��.�LLLLd<b�რN�&�c���(�)��PL��5�����#?G��ǎX���.(�<W�z�].�k,@}���L`.��H��R�2���:�����eQW��x�=ԏ���~K.J�J䠸loLn�O�?�/c��~?�G��5l�8�h�����:nW�W�-�5J+��(a^Zg��º`�����o��{�V������F���������A�9ʀ��jэW����������	nGG43m���ad�i�PC�H�
���)�d#ݮ��B�����Rxs�y�&����@V=9�,����^����֪�I�.�8)#6��|QO):���^��H�92��C��3m�fv
��I�s�_�}D��t��Mŭ��Oԋj�9V�JU	���}��{��K�y��KO�9?��&�d��P�'���,�l!�E�a8��p;V�TU4�85�������U*$x#��[��_�gMLL|H��PZ�\{L���b6�ȧ���Y�dU�j���n�k������
�rI갉Up[u�n§8L���c�
ˑ��L�� Ѻ���ͤInm�%�a�8\S��'S����o5�Ȅx�I�$@����&�b�:���v;�u���w��E�x0Cg�#B�b�߭.�5�A�X�	e�cv��f���|�=�D~�㞙;��Jx�T�$'�"��',i3Qű$??""A��3�ʮrHϼ�p�E�L>�I=�&Ҡֈ�s�ٕH�n,A���{/��t�>+f{ J/�6|��w5�F�Tk�^eԜ�5��p}#n�v���^���0����ą����y+ls�M���1.����㿿�U[nh�;�?��8111�B��t`!�!'lr}�����]#f��lV�9j% �9@���'p���Ө\I�!h9��[�ǌu��[!����r+����X.�Lȋ��]s�(lqF�I���㐌>U��t���R���>J�!#YS/V�Pn���"��}���y�ZDt����|�z���~_�k��������1�䯥�x�A/Q�t��C�I��:���N�z\���W_��`ǥ����u�k�r.��YԺ�8�����뼷�G/K?��K2�i/��W�gX�a�PX*Ř��_Ͽ7�<~������M�/��>��d�c�E7��te	��%��71�w[��u���6��e;�Cr) �V�Ma����)�����K���0ۓ��7���8g�af�u����B���>��o�1/�|�:�����-=�����>�u�]�I�t7�����2�!�dI�h���N�� ԋ�.Ir�<�	U4XR����H,�N2N�/!<V�#	��_t��	REj��*�`I��S����[MAZ�E^63~�?Ͽ%?�-r���� z�mݼj�^�m�s�Ha��>���e���w� ���(V6�V�<��w�8��x��m5xG*O��6s�����[b���Ɵ��Y�f|P�s��e[�*L���6FWk�)���FN]Ê�L/��nPV���D�T�HB%Z�(����QM�*~���w�.ʍ�t&/�!�\'����qH�7L>����~i��e��a��W�V}��G�<J[��~��:�2{~��z�Q�)����M풋3&�=Et/����rD����/���gH���x�/�G���:?oG�<��n�Sݚ��xT�����)t���K�/��{����O�1���$�ft�R���pȀ�Wb8C��J��`�����t�y'p��`21111a!
Z>Uil�j��E��Tfя�^k���\?�o!@R����/�:jB��N��g�#����Ji^<�2�S|ꤗ]�]���^�q%2�C�x�re4p�Z��]���ٷIL�2q6�y�]�%TT����\������J�Z�U2s��<rJO�wϠ�H����nN:/Fl�h�E���T����������s�#�xr�Ȅ�Ȩ� ���FG������1�E1�����϶?}{���Ph-Q�����9�`�
�c"�t.�t�J��(�$�����T۔�N���}le%S?�p�޻*5Q�������-n��3�E��ӓ#[�Oo0��*ݧ���P^����`���t�t�������2����a�P��6����wA�-����?ǰD8n#Y99��6���p�)ǽɴ�b����>��5��E���\�\<B�rꁖl��§"�r��+@��|����=11��S�wB�w���-]{?gl	#8 \��`��1��@ �H��D)�M?Nj��!E�D� ��X)�ɀ�+����2����nSQ>P;��	L��ʭfA5������A���&M���K[�=�E2Zb�E�ڼ%����y��y��D�}��aQ6�9���ǵ��'���/^$	�q�GǗca�>;H�zQ�����*������~>&<�~bbbb�|1���/�1� R���䯑���V��bCm?6*�\Y�9N����j�!	�ϩ���6�GW� ��'���u��a�g��I2ViMGgR�@<ȏ&�o�.�����^T�t��BrfȠY�>���\���0f��!s]���0�<�8�tO�ы<칵���}l����r�C��<}��;}�x����_��x�F���A2@(_���xyl�!���c����8��h�=�]����Y���r<��['��dy�(�,;e�Iiյ�E�I]��N��ڊ�R&�q.o�8�q��RA���*�d���uvI`�D��B�^�	"	����N�X�$:�p�u#^�7^�W���'&&&�Dk�s�BC�k/�%����2f��XȞ�����; ����GC�F��R&}rrG	�3�us�Yc!Y݃,����,j��@���Ɛ��F���:���M��E�I�N��8�.'?$k����m�]�dP&�ó�_�<ji@�ɚU�V׷D�/ԘSj��'��~{Db�̓WQ=��,9�.��?�>�}Dj����c��=�G�����}nǦ����B���il�KG�M��/o��_i<�'�w���ty�S�_����{�9�����]z7��C��-yLLLL�`w���"��)�E��$��d컁� �.){yU6~�柸����ЂWɏw<���M����\����E�<s�p���z�0���ڻ�q/N4��(��K�7Ө��%�N'�99��@�Tr���rSBE�:��O����J�j�3Wӫa�ԩ�����RQ��(����TiKR��VG1� �����F��H��yv4ݫ����[��v#�Qm=� ��g���S�h��*H�8It[�y����v�*�l����x>!=�y���h�l^qM�6@<-��{u�z�q����U�V�#i��+���ݟ� �Egˁ}u/�������*���T���a}Y��pR��$�H���h��������Iy���'p�rj*C�=�	]�d���,�E��/����V�A�{'��7�w��5��$/�$<'&&��q��Z�i��G�D�1���X�⌨�T�x���������<}��3ǒ���]4d�T�ROA"9�c~�XDR6F�!|R��z�g�3l2�9<�t�#�ի%=L�����%v&.���n�<I}���g��*�n� 0��t�5~�-��Kv�$E4�_o��l�q�{o��6���EK��#R�x�c�/�'�'� �a~˥����~@y�t(}�uXs����5�����us����WEkNڤ"K˳ò�?W���b�s��(-e�ĥZ�o�o/��7�٣x�3:�ڵ�������_���
m�%/�刂�~��h���J�8�G 3=��:S��-�7����dd~���*��\��F�a=�ԥ�����ĉ��-�/_����)&f��؈�+�f�mO/
�g�	��K��᨝���,��/kq&�������gо�\�6gdu��7�l.٢"����c��`ޖ�'��vQ�V�ֻ�6���t��v�S�r6��Mˤ�o����po����h�W�5�x�>|�f�Ѳ�I�~�T�.�[S���f@�'���l)�a��<�Q�ֳ7���)-�|P�%�C�z����9:Ǒ~~؀C��_��
�;���tꄒdk*��O��b�[������ոTA~K�Z[JD0�A��uy�^��l�M�:�X��|V�趒Ҵ0��I;���%��N�V!j#�[�f*c��v$Lp��)���D�O���.p�û��IK�B����a�9ƒ?��|�͟P������W���,b���p��T=���I&���+�ͳ����;���k����p��vl\C�}I����$R�GH���?��*c�������؝�G����|Xc� ���=�Đ�@��:?��|�e��G[��0jԺ�g�8�+k(�./D���w�ΓO�(߃�5)��BzA��n��I�\�E�N ��YQ�,�*������⑕�U�yz�����A
@uL�|� 'xȕ�6=���>G��Q��^�g��^���5Ty���Ӷow��\����y�H_�xxLL������1����H|
M���� ��4�9���}���]o��2�_���&>*>J����y�5M���S��\��%��U���@1��Ԯ�4�w���;8��:L��2@�co(�ls�;�����2�.�aT�Fa�|�}bb��c�q����by+����hk������B�gasdGKo�<N�"3��IōHc�	���|,'�����9�����~��I^B�#���Rц�ɀ94*�L8̇�0��!��|zqA�^:�����X�MS���<xn���zh�KNѩ)�ѫ��:���4�U"�\��Y����vLA�3t�Ǒ���X��uKѻ����{\�n���u�l �p�}Є�GZ6w/^�Y'&&&�8�\s���\�R��G���p�c����k�6tu�G'��tyѐ�P��2�D]$rP+�	ُ��9;�3�.��:������I�h�Ł�l�uOϡ̰nBm�.�W��M�IO����s��!��>�ߌ
l����8{q�n`�䶥'	�r¶��v���m�P�Y=pw1k/2v�z<�+�!�[r��)�bJGSG����@����qF=}��䥅�1~<<ۻ� *�yx�������<�uz=�q��"y�w���Vy���Ƽΰ>���>NpP"7��}0�|��:\�����Wg�#��G�����#Q,��6�p�Z#�����7G9�%Sψ�=���ͽ��A&����R;}���8�}�!�t:A���_c0�}�����pcerH��ɪ��3���qUݣ~��@Z$�SC�-[������l����)���r��΂�K�����H�ˑ�bw��u7�p��
@��E*0Ĳ���T�y���y�pڲ��{e����z�:��8LO�x�&<��8X��1����=oY��S�H���n\aK�o�%��AQ(m���v���iI�e �ӣ�'���y��n�\��*�z������|NLLL���n��p��+>+�6��>N/�VYBh�`t�|��s��К��2�㍑�Z���x������~��m�����O�����73Q>Ppt��,����2�Q~�N *S�C�Gu%�p*6��L��̈́���ptrG�2J8r��l^��w���zDFE�-�H���F� �~ѡ4�co8kU��9���ɩ��'�Ղ���,Ih�R2 �n_R�F"�J��o/2?o7w>�y��[/o#�7�p;�G_��H2T��7x�'.�h�H;��pt�<���G�{4��x������pc�ĳc�r}��m�^e _�~:kY�86c���
J�}g쑯,�s[��N���"��-1w�VB@�8�Vw�Xh�l�����P'&&&��6�"�����n�<.��:C�"������:�-�QŒ������Q����ݏ-�
-��Ca����"pq�.`�C_��N���;��nVJ	G�/R�����l,&m$
*�4>uDv���nr��z�D7�pqs2(爑0Nqj��^�k�Gjz~[a�܎��Ge7�&�?��eKu�|zf}� ����1�A�	wn!'��&����l\������{y��h\Y�o�}5YhLllA�U��:���4u�������͝29�)ިKs���v��e'���\�2<H693_����u&]��Kϝ �,(���J:c�f�#��voUqb9VN�6�E�$��	iז��\Y9�'։�o�7TG��}8PXm�!n���@W<�
��r;��ēᎸ��mB]0�n��1C��.����'@��[������m�yc^t	�E~�n�����,ە`ߖ|�����:5hPOH�-N�Sm�܈�+iӢZTq�,��7��yi�	a���r$/?GgO��r����q����>'�-�k4�H<��N��K;�G�L�����8sҶw�H����o�T\=�����Ո��<�l_2w��oٔ�����5���9"ڬ�q�i>���mq'�Y�wv2�X'�[���{<
a��sS2�(V�E�2T�G��A�e�$.'&&>
Zc�u���T�]�-yA�Ӥ@]�9�GxOk�~�G���.��#ɉjW]�H0�2�f�F!C f0(F��=�"�y����Y �s�YP	�tȱ���$�q�����rSuQ�3����bHU�QF}������m���V�k�9��w�������N�&QG�m'�.���)��Ss�؝�ۙpGvԞ�Õ�p�`K?fc����_æ�f�?�r\����{�c�Șz����Q���c�J�����Z�X'z�����o��{ǽ�?:Rog���W����οد�E:��n���ːnQ�M��"��-�m�`BgIt�d�yqY7��Ò�~�t���<E	���4X��Wr��]��6�D^�u��[=�_vK��iȖGw��j/�3�)����q�-ǯ��>�D�WD��S��N���U�����VN�7���3��3m�x�	�����g��=��ѴF�˽x�N<G�kO�~4�3�Y
F�軩��2�B%&}�{�L�Q���wV4p	�ՕZj(�,Y�fwV�b"�I��8a��'%��R�'&&�
/L���Z(����u��z��Cu?
F����{�o�ʝ�4�+(	�&�X���D:&��JE�%-<rx"41kfj�]hMe�i��R2G#\�q�� ?�p�K	=c	Ǻ%�e�/,Ay����n���?�rĎ[��^\6�u���4���x;��1J�h9b�H;���	�v�����Μ��$<{&�h���D����!��w�f��=�U��N£c������C�d4J����w��:�J7�]k�7����;��?���YN�:ͷ gr� ?b�6�%
K��/R�e�.NGdue3�z.�{Ԧ]���o<7��V\6��a��:-�P��j� �t�u
��{V�E O�:Ө�c�����N8�=+1��C�u������#�.��q��������z���۶���n�9��a����w��ٿ�I�m��xd??*���uU~���v��ǜ��5�Q䴯��[�s՜W>7�u&P���S)������M��FʯJ�;g�MJ�#���{�������x��`[V��P���x#>��dD�7����^Upe�X�Y�*w�U�e�2�;L`�֧#u�\��@N�[��!Hߋ���g׶C>��'�I߫��j�M�'�"PVC4*�h�%��y�˃�Ύ[-5�T,�\^�T�n����y��G���S��R5��2.�s�?�B��w�ޡ�*��5N�c�U'bX�8�|mn��2���w��H�
l����=�*CUH}�I�5�w�N-���ա�t_�I��`��A�o����ĵ�Ƽ�G#װ��H]�1��
e�zs��<��F�3�}&�!�.,�[_���?��bБ��!�.RZZ���$��H*{$�*9��:S���j���nT-�P֌���[h7]���9\�h�B(2��+��q�Ϭ�`kI�z�\��$z�qL��n:�}�ݸk�����0�c�Y�����%tb��?����;��l��0"�c�-z��e �ܙ���'j�G�l��F��Zxd���ѰW�����(���yL�[�����pP�`B;|�I|��u���M�n�Md�+TB�#�"Pm�Ы�F|1kFn*$Gfy5m��v�O$!O2��N$��oF˟�$P�q7u<H4sM*W�Y��^%V�kE����s��>)���n5�3��-d�����Gv�g�5��z�Ֆ�-�w������S��0e�4i��If��[�\�#i��#�h�y�8o���L�{�̣)�Bg�?�iDe�uo���R`B��hbf��	l@�d����	d�D��|M��?{�	���<���w�Y$��@�&�RS����B7�h�X�ֈ��r�q���e0n�N\o�Z|ƺ�[mX� �3�aB��uz��"��w�9{Faގ���3
�ƒхo<��Ik˻��)p�K9�Xƶ%�� (H>B{��w�����T��5����k� Ba�s���[FP�}�ӎ�2ǭ�˂�}�F�U]�[�j��1������ĕ�Ƽ�\���xX�ݴ6Ԓ�πd�>��g�?�d�uNX(O(�� K����s[�
%݈��
���`�Μ�r�7�[������Loηn�m��meO�q��L��'���lP�`[�t4*ຑGJ���Q�H����g<�Bx^�t����7\'ٍլ����>#�ͨ�E4��	���3��)�hd~�s���N���ae8�S�>�
��o��T���|�+��@����Xu�}z���mp���#��댹�^3b�aǆ�aǞQ��sc�+C�`{��8<���j4&x�a^�l߯YL�dbb����^�g��������%\�$����w�dR���աիpt��;�E���ܸEx��W�Z���Q+g,��X�Zf����\�~h���pSx����M3o1�L�WL�����iSo�F��6&?jr6j&2r���%$[�R׸]\�3.9���`�J������&'��K�01j�'pH�0o�v��\a�.�?��uG�h�5S�t:�d���θ��tzUQ�O�@�U�΃����O����#��q���n�V\��CӍ�"j7���n����J�4� ���w�5Т��c����~=�7�����b�=X�ZMʕ1��x�<s�uA�1�'�瞤>�K`4;E�3��	kڼ�����`8��J�{�uS���x.T������BjN?�	J8��H�	��52�w����X��-�z�K�7�2r/y�z�Sc�5�g��"�W��rx���-��L9;7�Lr�W�<��+hrreQ���x:	����>�"�ɜ��Y9ݸq=�m�w:��	czQO���R6�v^�"��vr*����}ｙԇ܆�i���{��{:�51�(�lE�C�䷄�-cQ�'n|�N���C��z\����m���J{o�����3`d��qtZ2�M��N}�ֺ����k�ʏ����B�0�S�ϼ�7����v�����cLC���b��E(�]k�dYa����qDH9#�xa�`4�B�o�����Ꞵ&�q�Ɔ'U���{�L�J���5�L�4�p�����є5�EhB� �#��P��_NVO.��h�ZHˊ��`�U$;�C�u�]7�s#B2IY�C��.��w�v��:t���or���V�T+Vy�#��[�����l��n :�j� �Q?��TxdHNbU��*eXkW���Y��i!Em+�^�l��8���>J8�i���������Iy�I}i�*��5O���9Za���G���n�"~b.N̴��rvIɸ��v�S:o�f{�Ekq��<Xy��~6{�g��hٚ����Åb,�K�hҋ�<���s�z�r�Q�(q�=��������C�C~��D��8=��Md�M,c<G��^d�3[�ݖb�m@/�wX��C�������l���a'��pC{�B����c>���^��a���r'Z��EzQ�/LLL<FO�j�5�����v�Űmc楃�G�"�4�s���8�@�v.�+N����Z�=-t�Ś||���P���\#ɩ�7��{�tm��w��{��U�����זgں��Ϥ�R@���p�{�
��}�.��!�m�b��{��1�|���#�P�jh~�H����oQp\յD�{��?w�̔KB`p�T���wW������*�b�ɮ�ɖ�8��ӄ�֝��H�U٠�48�EMS6Ee��4^XS�щ�X���tX��b��\#0 �HE��&��\���0�o5+f�.g4 ��pjK,a�8}I���jQ�D<o��ڞg�x� _��4�b�d�8u�����*�V��v��'p����&���Mr �C�&SBJ�����6X�`�w�0b�~��m�~k��'ͤ��F��{C��n���8��F���������jA�$):���q��1l�0����c����WE�@n�������:U��S��7=�z'TYy��2�|*?���[yﲾ\������'��L���sϪ|�rHz�[D}m�ٲg�깹�q��eJ��a�������|��¼���O*y� ��:��Eu�G<�Ġ^�&��.��F���am�Z���5T����ǖ�W��8���q%�3��;�����5x6�3G�I.+m��X]jPb�)���z�|�T[N)lcg�v��G" �oa
�������de?N2�YQ+YM��rrݙ��%�	Y�����B�I��W���gȶ�G?���U��m���c����#�όf΄'�1������`Z(�*�94������-]Ο����Bq�}_���H׈q=7���g��lP�A���Qv�A��zq�,�Ըӌ����n4�9S��j�T�:�О��d��VX�g�R���c}͖�bd!L��I�1��t�R�=%�=Z81_St��� �l�u���<�.�EWݶ���#����Z�g�׳Wl�^�1��Y|�}mʫ�<�a�|����S�����}�E���lr���?�XQ�B16��{��T^��(K5n� f�yi��0"�,-~&�Oj��k��>����E�(ƺ��id���m3��IYI��C����y�#���4DL�^8�����Z��xN�����}���k~vt/��z/un��!���+z~�B���j�'���
��UwÍx�I%�a������'��c�ip���t��� r�t*��Zyr�w��#���7��r؈A���C"j��ҡ�K�%B-^�{ߨ��A�F�;�Μ6�� 5�߿8�ߏܺ�3?7{��٧� �ƽN�M�4r�6��/ly<���}4afG�M���t�>Ώ/�qf&�(�����}�T�2����c' �ޛS����v��(9��#뿰K7+��,��$�K��*̈��W׫U�����ϣu_�`ߘg^9#���QY{��Ż���m���?�1�c:��8.q�]�E�C�%/>M ���(�8�����c�Wr��yRt�^կ���0~�����
��o��l��ԯޚE��2^��\6��8��� ��s��iE�O6@��T�yT���ͥ�LS���Gh�C�60�������JG%��U���*L��%�ۃ���"_�*��(�J�)���1�{�H�{Ӷ����w29���g��?2�N��8��u^��O�7Zq<������mhL_����S蕥9$��9��/��o�ȡ�ĎÉHv`��4��>��?Q?�N����[ps�C�[y��X\ս�ʞ�����n��#x�߾����Mb���U����۔x��N����D��������:�pM윑��-�Sd!�a5J^xo�.3ϝ�)�����o�TT߹���2��m�Z��ʭ�<ne�/����w0A�(�b�r�[�Ic�oJ2&>�+/4c�J��2]�[��jΣ��n迮��M@��Sg9���;��kV��8���;��K�-���%7�˄ൃ�K��%�X _
Ҏ�U�$jf���4�V�i��Q�Ϟ���e���1?�E0z�1���z|��W�T��no�H2�=�����������[�����v�����G�����fmo�%X�E�{�&_�Y��S����)���9�>>#�ӯP��-�5�*f�����A-�g�MTWVɢ����R�)�AE!�I�@��n�4�|^���m�ǻ�-�7RP������~)�s�j� �Y#���xO��ˆ���I?� e�j~7�M��x�0�P��U^O)l~~#�v�ɣ��Vz�R��:����c�����
��1CVɼ�:�P�Q��Z3,�^��aX^���<�����
3ӈ�I6��JsC���e�kFS2X��$L�Ì|��:�h|e�&W+@۶e���K�=��՗��z6g6F�Z����:��3�r�tu_�J�wۇ"�V��W���W�Pzm�I�ÓLv����n�g떏�\gK��%�����w�3F���8��3uG߿�݌�O�w����ü��P�m���ʺc��R�g�6�l�7���l��������_}����S��J�ge��dS^q����
Aq��\x�k9OUP�[��������ײ2��Ow�*�Xڲ*��>�{T	Xh_}�Y���p$% p3�������.j�������k�'��»A�+�q��q�L��§��f[���%����hc����+C���WF☸�����oëO����ӷg����I�1����2�]�O�8ʢ�f�-6����0�Z��M���xo�� qv�;��
��)$B>�-�s��붰�/��F����C9j�N��E��y��!���q ����{�LCuR���Xu��a10�IAٹ*$]N`H���["Bz1�Hp���ڳ�G.�KT]������]�Ey3�4�O�^3���֘Z��ʡ�0��47��0�ec�x����F�bLk��x��nF��:Su{��d]�Z�}gȘ��
�r�c���Ni��)�1�?@���/\�t�H�٨ 㗷��N�&"�������vO�Qx���ю}���py�4S�y���1�>UBeV8
��y����C"�A�_�-8=�x��������YΤ로�X��~��^��t��p;�'u�+��)��a�[��NA��԰yF�m�e"\�O?>(oXN�m!�S�h���\����#f�@�~���� ����|���XXXX�]��D�X�%��ޏ���i���x���@q��V/�,�,���n[�y<�����o�1�p�H��`��ՋlX:	����Y�~��.\���Io�{dX�"_Y׻!�W-3����XV�ޙ�OF�]B�"Ǿo1�3ovl���ʀ�xL���X
����J�������1�Wљ���G4��5�M�	����G���7��E�*����JL0VbU�f('��:���BXO���s�-ǩO1VBAR^���P+'ڤ���e�Z�G�q!��@NXl[���;�&a-���?���N�Nj��	gH���ԵQ��)�P����s�R���읷�G�(�zy�W�B�t���Kn�0�&u5�Q�̳�����q_�o���y��:�¿���>M�A�e��؎�������7�������cv��k#���q����|2)��&g�L��	$|#������'%%�Le���|��I�L�.e�%[N�C��m��T�I���>F�r�%Ww�('�0��r�QޡtM[�aC�y�H��堓��� 'u&�'�� ]d	�{i�tV��h�~x Z��� ���o�ki"�v�u����¿��~v��H����O�|���!��������Q�&�)���˿�!�������ёl����$z�B%��s�W�y��� �/��@Q�A���O
l���q�j��"f��E�K�U�Վ�o��j�H��w�U���|[ӑ&�e��~^��AtEJsO��xl|�b�b�˲ �z�祖�� hń��r�wGG6v�2�N#jCbkG_t�f�=�mn��[P�d%�8�Ó��!�ʢ�ش�����ᱩ�C�>Q��ͬ�+:�k��`Z���N.A3qf�|&a�U�jä�T����	c!݊b����Q��#�v7�<
��J�9IgQ57Tˎ{�`ļ������v�|���q���=�?�u�����~nXy��#�� ���H����Y��}q�ˢ�;b���(�K��r�1��n\<��/Cy���M���c�	F9K4��Dk\XxV?�|��.^t:��Zh�a��L̺̱е���6���V�����nS۾���E;
���Ϟ��-�~��lr�BP�P�8s��ng<TP9T���R��T�Q�1dcOlp�E��S���k�fo�R+�EQr= ^or��EV�oq��"O�qWX'�6.;�*RB%�%*���QYW��B9}��>��\`�U�s�c�U�m۠ / Z�"vø��.���S�x�<�P�z�/�m�����Vg>�i#�7Zv��~NAOиը�?xT�B�P��mKI���8���QԖݹ�봱�O�`����(�Hh0�p��^U�.hQf������[:N[�ڡ"�2�T�j����|��6���oU)����:�h��P�ס���׷L��;0��f#I�07�D��16.�᫙9[8�A���f牏=RX�����Ee���?$È7�6<y��̹�n�_��}C�A�R���h���"�>������j9nU'n�JF&�f�q��rz2�<}���,y����[lkUVd�>Ȃ��[ɬqZʳ��b�&���Mg��l�&�Z(�ܿw�Y��9T���a�S��:�I���z�*�E6
��^����^�K��r>���3V1������F\����=^��,,���=�1~N��1�%��,r�-����۹n�@#O���v�p�nq���y��ML\���Lm��Q��5��I��|Ŏ�_�!��OT!�u�uw�gb�.\���0&��>V�G���E,�P�x��S.F�L�<����$/�>؀���E:�av���r~R�����P>l?��z�T<yoɪL��P %��<��W]P���;m��o��V�w,,,܅z�{� �j�π<��A���<ؓ�Bv�x�9g���t6��
�`�b�݈����#�en�!?� �|��[��'P�՝�5gi���Q�F��I5>Q������U}i��Ű�F�J	A��0h��>���Qg!4�䛍�-Hov
"����7��4s�I�A'Zjɜ��@��V�����W� ���Ԑ�k~g�o�4ה�єu�㉳Sy�rl�jshO���4ךa\N�^Zr���N�°J�0}-:�[��ZaŸ��?k�>�@U}�wj�}(,��˹�N'��Uq ܶ!>��H�S��w�<ek�Uh����W�T���<nERk�Y�Ë�4ӯ��~V��\�^_X������S���x���4�G�c�}��B��=�g6𕑇\�ɝ�?��Kw����&q�=ŉ\�JB�+���Px��g�K�p�`��k�QQz�16�� ]��č�=�=����`���L#�Nˇ܂I�SHE �JrQq��Uܧ���>'���7Ot�E�oNI>��ex7�b�uY8�lhO�gK��6'�l��$r~�9px�q�L�R���tɗa��G�R�6��6'B�H4$v*_ϭvv��=?��D.,,,0���;��X��0���h@8�#X�ÈX7~^1j�^�b��3�.8�}p���e�w)ՙ�`��/4i�3����T>y�=fEj�E�ژ��F&�����*G�c�!']3���rl�T�I'?Z�;��0�mu�i:��Fdo�9J���'խ }�y�@(�yk�>��6�|rL�'��d}5����ʅ"����>�7}۠��bNt���@�oRd���p^ws�e�_XXx���c�[�"89�v�?�u��+�9Z��lγ'p���(�����à�&�B�D��W�f�2%�&�z�}MZ��
?�����٬�49�ų,u�t�`�a�rzs���6�}D�N�y��y�a^��m8���	;d�{hŞѧ���Mh�o�������0��M/����_2e.,,,L�=�[�}f��ι�3ZO;pl������V[���K�Q��9ʸ�F]W��=�x��&�
5
�Yt���N�N�A9��h����v�k���σ�g��v�~�)cj��!�i/�;߶�IJR�u�v�b{��9�B]��|xG�}���\Q�`B�$��d��YG�q��OWŸE���l��0��(��W��6��r��a�Vza0�0/1J���X����r|Y���|#��A��ѱ�u,�R<�%�cQ4aJ>��5�H��~��D5PC��]���7�o�6:>\}���;�[卄?s���hq�	E3�(���q��/%�(; �\2D5�B>3��q>��|ۉf�G�����������{��i�6��[r1��0^JV��]PL��&��8q�7�7�׬\W��N>T9o�/����:��&ȯ"	�y(�t���z8�!m���[�N~�	�>�Y����0/*��9:?����Gu~�dJ76z�|9~�;��kg����y�}F�J/]
j����!�לX�yt�9\ ��H�?����_>����C����߳'C-,,,0<�W�-ld��]��B��"���WY��1���q٨{x��c���������DA^��a��4�u
GO<�+���y��R�Q����G�i]#6�b�[Ĩ����_�93�.,,�������,R�V��.�Cg��8���%[���JDN������X�z���1DF�}�Q�*Y��P��G�"S3�ㆽ>�k�NXY�y2�E�8a*�`�GG~�"qP ���M3���H*\�����-N�+�F�X���*�{��5r���P�+���4�	^��Tm��#�H�B�^�InXɭ���p���*��Ql�h�4�Dܩ(��o/���hhl�_�ݧLC��ipS���B�\m�~O}%ķ�N.�{�{-�{}v��p1g�-C�ށZ�B�[�k��R(�b�������fɜ达��~w��~�r��9}�w�X�y��t�	���Yei���9{�����ٰgt�^Y�����Z<c7Si���s�#�d���)�k�㞁*����$I(��w�j�^��m����������ʈ���HO�b��嫢O�
���	�q�W���Hz�Y	MI���E�NAx*�5'�p�uw�}��l������8_)W���a'��V���+�p���{�1$�������L���Σ��I��Ok�2H�{�>�޳6>����ot���!<��/�������i,���<��ϳ�ǒ^�^��a����SN�+��:?;���G񴞳����[����AaL�����F�hց��w|������'�TƊ꿙XC0Z_�(���� M^_XX�^M�7 �ņ�;�ZN5�Ȑ
���c���(/��v%�]���|c�ܓE�I��E�B��%P��>��6T�(,eh�k,� ���_�i�;�X�@e����0�t�����ͳ���Z�x�̄yyj��56�봟���v솝�ސ�etj���K� �8�����:�xil�-r�9u���d�y����B�z�X�\���'�R̆��q.��F'�oB�۫�����SqR�K��u�yC���C�މO}e'�p�ɴ�1�����WZ��:��͵�{�hp�(k�S�/�V���W�-1�U ��8BQ:��2Gg�4��+�"p�a<�k�Em�L뚫�s9FO��X/��t��r�����*�N�hp�ǁf�^�;����"�@�&�SX�Q-�8ۍlm%g�g��l Z�Җ��Q����WC�W��k4���h�8sL�uM �uYW�жY�=�~|֨=G�Ju�9�S�.�����l�yQG.��*�{z��T�2{}Q�G�>���bf���1�o�C@P���~�Iޒn��n��@�$Q�~r��͞����t!՚�<#d'Ha-F`���Q��_��wbH6�*֯V�tXl��&�M�&��g4u����9�;�TX����Xw��u�6����uv��5�A4�r?�UVS�g��z�[��f��g��1z�3�$gF�;<nA�e�1'�t���
�A���h1�������5kė͍��&K�K(���/��v?����[ �=����j���śz�N]�C1j ȋ �"�3�N-�{"0=/U[�5���^<G��K��Us���;���iGM����6��N�K=K�����-�	�u������d�����r�����E����(�����? ��N���WaҘq!�^�r��qaa��:%�WI|�8�J�?2_r�����a�Nb���Y��U�|/ݩ~Vr؛��8O�G�y�w	;\�m�_XXX���1#qҸaA��x�hc7%���X�׎�_9���Z�2%C$�"煵�.�i�
�X�y�va��=����;���V����,6�N����(���7��Mc�,"�4v������E2qj����s��Y�vg�dn�fD�Q4��`אړ�lX,��S�:mG�VƦ�^:��=�gS���+a�!�'F�Z�?��8�UW~-�390�V>��gr��,X�_G���|b��g�ORI'E�WA�!����h��]\�"�}�j��.��Zgaa�Ӏ���	W�0N�e�����1F�s��#���y�&/�'�=r�s�ɴ��Z�i���9C�t�X�x/�%]�":M���%���Hs&�\T��QLU�������$�_R�-e+�#u����)=���}z�(8�������r��m�J����m�Ζ�Xu��Y�����(R���h�	�s4oa�_��ˏ`BQOcH�os�f�|�a��"WYXX��7"�J?0�Y�����rځ#�/B�)�;5�'��qw��'f� 
�a��X��?�P�\�T}���"2QMD��V9�#�l�lG$	����ۭ�V���taa���).�%y�}�. f햽�V����ر�v�o!%o+�A���70�sZcrORt�`ۈ�������I�g��wb�2����s��מ��FǬ�Ü�)vH�zbT�̻u��t�P�j�J��9�	�FO�pU-/O�5ҝ�7Pr6�F�����E*촜ٰ�z��|�14���'"�'�3��N����X����w��I �X�:y�'��cc3z<��DyA��.L��d#�q
�vVq�E9J�V*�[��O�#$]�{DٲN�d~�L���>"�zn��l�-ϲ�����
F�Z������,�t�h���q���~Pټ���3޲|���=�V�ۑ)������\�;��l~o�=א�@��U�5v���,��G�_(/�G'��sQ�JM^A?���C���@��r���U��N��x�>ʔ�s�ο�7��?�d�0�~Ԗ�G"&�WO>���}���p\˃܌�@�r���[���mŻ�s��E����d֑�䯹��<�8��n,�x.M"{r�)�������BzBm�� �����������ɾ�Ӌ
�������3�p�#�*��O)���ݞ��2t�-�	z�wzo���\S7�����t��]1j"���JF�B���Ĕ��K�_N�h�d��񅅅�c��X#�����<u���ע{����{"<�LNy���<W}��p<�n%w���#�eFVF�l��*�F�mS�CBYL�`�p'6�Gv�4(�1;����W*w6BZu��h�5<�m�b��_�o�� �P��v����8��*�k��p<��8鬯K4�B����eק9���s`�@�D��oHvVY�m=�A��+�i��#��O�C'������7C��G��|����Q�6\��I�.�����s,�乂x�قڵKy�0�w�ɑ;�>�|�ؖ2�/?�L�v��WI>ԡX�q��@б�č�|��w���*��5�t�����ϏZ���^�JQ/�F�<�f�
aV�1rj�)��뻔�P<lZ{^_��1���r4q�F]/{�s�@�At���	�:�9�����]"6:C�5B�<jv�veUe����J�|��p�+�#�Gn%���ե>���$�AnA&nu:�!���Dv�?���0��p�=^4˙0�#�q#y<�۱jS�������x�|�f�ˋ��k��0N'~t�G.p C]�w�2�WL��U� �e��`���Y��0F��t�\,��+T�M�m�lcM���h�c���􏕯��� ���fKmG���1��R�1�B;,,,,��ʨ^�q49ۍ/`�\��R�	!C4��x��s�H骬(y'�)M[�w�gP$*�*x��W���2��_��xg>�{*�� ;��� �q ��p�)ذI��J��)O4\��V.k�R���H)�k�0̋���r�d襳��@XO� ��3�Ѥ|�rύ����x��Y%�`�l=�S;G���[~6n��u�8iW�Y`�3��.�7��G���Z���q��<~=J��ʽ��$��Ms6�@�O�8[�������0
�V��P��+�k�s�������/;6���b��2w�<��y�k</�e���cf�������W���������� si��1w��2K1��f��	�tXJ��r
��e��[q��Q�!UJU5�}.��脩;�"��l9�p����3��`��	�Fª��PO����H��G�
a�,g.������e�h][�e�vx�+
s���ُ��v[XXX�m�{g��,�d���@^;�ŴE��TՑe�O�ƨ8������4@�:�X�mR!�O�(�e&�����F����d-,,�S�Ǫ�����S��cj1,h�C����mǎm��C�kf�6�!���r?N���xMWw��k������|uW�ݰ��K�Z�=�W�y7Y%��+�QF����Xd�{���Ʋ��|�� ����h&�[}M]�݅���iu�ʓ LeT�y����0ucH��BO�ؐ/8�
�WO>�~�I�k#��9
UE�4M�"Ll�C]��<�֐��lqx��7�ݍ���i���9�כ�H*p?��ǝ�o���7�F�`�������C��B����g��=�rhj��q���aaaa�8��zғ������p�(:z��7i�j�����A��\�e8OI�zꐦ��R;s�Q�c��]��h�/��h���1ZN�kYz��^�r�tO�ׇ�������p��AQq�#5s���LO��B(��J�ܳP9 ���wjI(SCw''L�0����Y����n����!^Ԫg=�;0�|�aN�Yٛ���|=��q�㴇}Ub۫�M��������8�q�?ٕ��,$��]f�Qq	!w���lV������50��T>�>�L(n[-��+1_i���߯a�x��F�.M������9��6*�ؑ��9�8Q~�Z�Ī�����"
�d�9bcj6�V�{ G^ �8�W�<0�X�W�`C���y�`#�ف�
�⼑2���?��c���h��C<W����ur���/٬z�\�qrW�bͧ#R1��ѶT�J��Ĥe��!:yz2�`���6T��7�za;�#�U�#*3�G�R�tN�]@4�VT��Yb3�Wo����촺;9���Wg����v����Ƚ��8^w�G��c|�i�ӷt�X�J�hI���YA�;e�T�v��H�2���]G;���Ҏ��
�a�ys¬�Z��H����:}'#K�,�Ǥ.�8��F"U�lZ"*�/	Mcu9����z�E�Or@�."�J�׺y')�9�n��u��ޟ��g��xO*�g�;�m)��P�s
�>�=#������fN�-1s+�[�A�_��02��������ܢ�׷d8�O�+�k����7r�J��H&����^?��@B.��:u��������tT������y��N9p�o<���#Ѿ�#Q��(\��X�z?�
-�;|�d��<$ϣ���o��2���;�Z�dp}<����C��9v4g�+�#���H|�Ez�5*ߖ/�z�m<��-o�~p01awr�= ���?'��?g�����ga���B�����#`�Kǻ��(�eeQ�O�/���*��ܴ�s[H&ʇ|�k���l1���#�V�A�x��T���r��>�?¾m�����i�;걿:fKFPzl�!� a�Q��l�ٻ�9o<�T�j�l�2���,�+kR[V1�����F�ϊ������(�XA�!�e[�R č�_�	� �vsk���[��{`P�0Hg�J#��d�����0�S�����2���Z���|�m�v�֚Gdw��h�����W�p	L)F�`��Y�W���3�Ǭ�Xf�p����t|;g��:�ɏ��y|��H�;䝹1��#��d�
���h����f���OS��_�q)����F�oN��N���I���1X��v��ăB�w��ş�h���UrJ���iF�7猪]�\�ȣ��mᱪ�$���D.Ϣ�k~xN\XXx?Zsh95��X�L�|�ò��8*�.q��Y=���߿o��XMv��s���{\�_Gz���IJ����!��#:�)�.��Y��mK��&��Y��±�����:�����I�������w�t������NAX=O�@��K3���U��eAfj�+%!|�}���X.���MPA���/�w�d݂���U:G9f�\�-grtw�=�>t�zz}K��ȧy��W��wZ�'L�5�[�7ċ&9S�Gu3��l�}�I��z�D����m�ֻÆ�a#��ͺ9����3�qr$Z��Ǽ�C����.���I^7�����p�V/��h��Y��yR�r�E[����&I�3�e���g��	̓��u�h���n�Hd.Q��9�+��cG=��F^=��(� H5i�v'��}a��U-���Z�vaa�3�F�j�0�^;�'<1�U���ɶb���{���R8�
�(��7�s�1��V<�9f�yrZ7�G��}��o<�,���a{�2B$9+rAN�����:��Y��6�9�h�:��s��Fn��"�ܠ�J��@��^��kF���@j��(��#a�'��
�d9� h�U	�X��	��۝�$G��mQ�F�b�M��d�	�>a�V�ϵƳ"�J�iy����P���r��f�z�he<0��:�q:U`�jښ=<��N���+I������r\i�����~�.�,����[$&�V�g���u��/�'{�����Z��L��`v����֩n��vx�*E*&�B�!���x&�����sQ�Dr��s>�=�&l�O|�گ�O�{k��Y���U�)��*\��+�h�= bd=^G��Q�q��PN)�j���弪)�$R�0�;��q�U���t�g�tw�w�8�ˋX�a��uyQ�[X I��Ы�(�;�:�6l��LH���Q��՟�bZ��ͱ[��qgk�|ё�~�y��÷��Ǝ�9����V���X��m�Oڜ���#�'<�W�9�	����E�����ƒ��2�'��u�cB�y��1;��9p`ޑ���&�wM~XN��y��S{săY]���_+#��6G���й�C��Hw�q�oDy��ca��0r��=S�q�\c����X��Y(�Oʰ����C�s���d5���?l��N��;�;�����]�l�۟�X	��=�;��Xy���,��E�J���"�{`�]�2@)�J��SRC�*O��e` m��Z�D�r�B��Α�Ԫγ�(b�{a4��7Sm�k��%��ʴ{O	k�MGv������+�^רi3~5��zM �%�횝m2M{�g�@e�ZY���G��K��x.I��r���[�7��G�F�z�K	<��)>��x�p���~��Ki]�l��Oɱ%�y.�P=����˧�������Ĉc��ϔG-���kS��1.��,�
���6�7�@�kibH<b?��Ǟ����1�~1�0:���	T�=��dt��B��Z}=t�U?�F�0��mc��%�վ�������9�	ON7$y)��2�2bXu6������Xwg�ɴ�̏�O�<{:��p-��\Ω?r�`�WD��V��v7+�m+���=�rsQ��Pݧ^cރ�X"�Zx�;�%�͉���ƭ���������_�|$�z���:pT��l)ϲ݉��=x8�|��_�*+-�/P�c}�Q-��ѡ�^i�H�4��kˠ��q8^���N�#�~
�O�v�ܵ�1�L�<�΋&rأ9<���jP�϶7�~�0k �*V	:�ip��J��
]R)���M_f.Ac����LA���v{M`t�|�pR���^D�U���k���m�{<7<����h��r��p��_xQ�;r౤�\C�ȎƳȯ�k��xj�k�3�ޞ���	�<ǆ��ِ�
3�pؕ=Y�Q[���`���N��_��]c��Oe���n9���נ�+@��cO����=�����Q�7{��(W)�FL43H��838G���:�{�1��x�ǥ�t�E5���D"�i哉x��:}���.��Fq�rL�K*���y8Ƶim\����V������a�y.�����&��9�:S=�S��5"a^0ߜ��n��b�P.B;�a�K�ZFw�&~���#����9�a߰��;2�&nU�"�ݙ�!�|�\�񼾂?�I�8i
��+�Q!��ق��*�{̯;.�0��.�K�Kz-I>[�f4��CFȔ#:�!+�E�r'K93������n���Fmn�����=��M��/��r�s����a��\v��Yն�-;�Y�:�.a���=({ �\����^��W뙶÷�M�>A�+z�߉���{�m�=O�`�p�Ͽ��Y��T�G;����Թ��$*�1�ˋ,4+#i!h߁ ��nC�Mк�Q�h-Bx��`�3�VB�ז��?[��N�d���g��4�k��ÞQ���d�;��W��8���RޝV
L7����Ԕ)���Jw��*Y�$
����5`��y���V&�f�6�$=�8�`��V���]n1V�i�xy��tz��S�R6�>&����������� ]w�Qnn�?l��>�-b�늆�X��]kE.���A���"�1��A��V��Gk�c�-�i]�D���y��dWa�����;	�[�k?�Φ���:�<�2;��*t4���at,��޽p�jٽ�� }�:l�����5�z�-N�������d��ў�5��m�Ϋd>�	U�I|u;�?M��Y����&��[��.q\���?A�x��DD�m�.<���w�O$G=K�	�gr�%����9��S��@Z��V���Z�!Ǳ��t���3��*�qx�����>/j���#ţ����㤉A��v���Q{�R
HI�M�tio��r�N���ے�'���y\��s1P��)%�{���]����-�5.s �a�y9�8"OWf�����2��U)�5�6�6u,q���VS�,���<�g��y(������7|G*�����~Se�����\N	�j69F����N�R���~����5%�	��aWyGSvh�Y����4��ΞI��S���5՞w�Q�ɛ~�Ux���t���j��&XȢ�3l��&I�;�7[QY��"�&XXX�K��ň���#�x�lw[�
��B�s��L6�1�q�b��p	�ʎ6S��M7���O�(�ڞ�N�ʔ0)�Q�wW	�w6�fgK��C���@/,,�MH�=��C��%��sDs����qJ���G�R��ص��	8���}}����x1��H��L�5(���bӓKM����cQ�U�q5_m�<rJ}nb�� ������2t�����a||���K���#�ض�=���2�~�B�+���$�5d����
3ys�2��5��5����7�[k,rddW�
N�c�32�O����S/��i��rT[��g�i6+zs�9{��Z|]c�H��j�m�xv�n﷽�}>^t#*+G��qx�P�c��_��ݽ�ޠ�瓽����Ưt\>Dܶ/H�:����i�#;h`+S:�Md��mX�tg=^�@��,��*q*��'��o���s����?��g��Y��_l��ܝ��W�}[��>꟥ �\;b���1�h^1�׻���Y���,��� ��y����fW����GtW!'�e�yK�7#:��8YW���	!ٷ�?wDQ�R}�a��9ۿZ�BJ�&;�[�f0�C7j\�֩>)/�Z�#G�c��)65+��au��I/��a��������Xn��6O,����*����Mn�a=NWq&�����GE� �s�Q/U.�m�\���ɀ��7��#�-*=�eR*ohˍC��B�p�${|����\W�7k���9�����g��O`�YYXXX�xX΃�#�d�7������I��_k�����0���"`���`�i�(1���3%��{ƙ��֓�v�Jy�]L�R?�hx�quaa�Fq�Hs�a��q+�s�2d�������s���]���z��.��r��}��#-��F�m�ݴ��D��pѩ�H�zR��2�J�rU�kh�φT{U9V_D	�؂9$/�)�%��ő�,���B&�)EU�Q������U l���:���c�~AEE�%_ی�l��se0�*��thxkďq<�U/)#B٣�+����+Ea��"�%��쳸K�?��g�m�����vp{�O�O��)�����xw�6O�O!��Δ�#��%K=��p�8��۾�9>Q0B�����ܫ��f�Q����36��X=j�\#n���(�?�72v�q�v����!F>{���a=p�9�N�<�3�sƺ졑��?U��U�e���R�j��e8����gvA�H�!Y��t/���"��%GG��9G�8��4>�W��)�MNߩ�H��G��M� ���O�L�Ώ��%3�HI.������ߎ^�p�-L9�}�Ա�Ɯ2ę��#�����{~IOs���+�z�������MԖ|��1^4i�A��}�����M��cW�v�wj�C��X��ƛ��c�����¿q2��n���ޏk'p8�����@�s�aZY*��$֐��:(c�9��UZGd�BZ,�����=� Wkg�O`9o,,�h�T�c\��h�I��v*_8�<�a��0�el~�v�_s��� Q%uI��+�"�e��`E�,tt�v4Z�{��Yz��ڠSfE�b{3�=�5)B�S�ݤf�"�l|
�ｔS�^HD�n�]����&_���t�:G9yr^�9J���ڰ����?c�� _%É���T|,ۦ�k��S壘N�?-; ��Z�����;P���ʄ㦆�Kۅ�޸�aw�o�X�"�1.xm�w3B�m�j�����D��D6ƼEyh����[
C�%�5o<�� V��˓�������yr��9b�2��mbcsC:Aύ;ɂ`ޘF�yI���kIR��6�$�޼\���Z�|k������.~�y$�ԭ��sK,MQ��
˃���=R:�쒿�1������Ci#/�R���m�,��E���m��l��=vd���w�v
:�f����N�0��F�U𸣁��"ı}�?n�<����3����z����8}���v*L��,��FI�	(�k����$��/9���0��!�^����6�o����T�ЮXm�y�v�/����jK-j��2������j�Q���9�J�����]��]�?#eF�[��%/�T|�׮@�&�F��Lє�-=�A&�ǫ�r���"�9Y��)������_�-�h-y{5�wJ����4`�w}��i�w��挓��|�y���S��Ds��t�8=���L�{+���a�MU�W}6���AFU�@'aXNK��|����J�+���|6,N����}O�a_�y����j����8`(}��t�3T����x�l�"��܇�y-��s���((�L��1�]��V�g.;n<e����N$N�T�&P��v���Q���7]ǖLgz�UrE?[X�p���7�\ȧ/���:�����)X�58ʵ��f�����y^`'ܡ.��<��F!�ԋ��=R��_��.6�5����tt�3�8�r�ʟ�)}�����1
���
+"��ϓ>s�:ʈe$�þ�J��^����-�\��M���us '�q�*,\sxQ���������хy\A��	�h�e�ȹ7=���U����ʮ��F�i��g�g��܋ﵱ�̜��;Oc�OA�~��;s��{�r�XXXX��x�Hy8m���o�� 
/ƥW��mK�����2W��y�X���zlH�G�]�QV�Jz&/I��.PތB>�8�>�$��.���o"�d�
��Q�i-�Uʙ,\����Yw�� *D��<������N��I��=Y�|Zy/,��
0�UG z�=��T�Eo�tQ�N-�}?jR���Q��A�>���JC�S=/��;���P��������������2F��C��������k�__�����~���!������ll9��8X�N��ӏ�X�N�bmj&� �ZD��{���F3[��(6^B���L�fc�C����L�^y����a�G��2�!ZF9�����a��i������H��{ً;a��on�_���O�� ���1��3�݌s+}���\*�vl��=$�/3�-�����7�)�#��GF�4R��B~6�(�����U-ߥ�?���������SYP���w\�՘���Z�	�ݧ�Byu�c'��t�*t����_���С�A���	;�,��a��w;#-,\��s��G9͕g�G1��ؖse55YQ��gS������|�f�~Ε��Q�Լ��vx�1����LpJ,��I �Ü0��uŬ���u�-���h1�L@�A�	m��b_�0�A���1��̺��Z(�t��8�^7��s@W�����������G(��W�;ǱE�'�ڃ�(:N�Ã9�0��r��(��ϩ�!�.v�q�quȏhyǙ���bZ���+���0���28mԒ����rl�j�Y>edn�����>!çaf�q��ҳMb|�,[l{{�/���K�n<l5g�<��������?�`�k��u���)�?�Z���Y��å�<��+T�� �%�' ��D[�8���KeA09m��FibOM�#TZEى��A�G�3S#���mB�LN���m]��g�,,�g}���=3w��3%��`�R�	��b6��ƹ�İ�-X���A��e�?��_���N:�����SF�<?3���]ׅ���-g�S�qttu,����PM�hqJa�1Α�@�ʎ0�㔝|иv8 ��65�|6:U�����\N18`���SFs�s5�z+��#_�O�!P]�nq��3�g�2Q#O���+���r�z��ҙH��*�i?��Ϊ���۱+{���j�V�z7�'Ac�g�t<�{���D�	��o���C}�|
�{��!��$��(<�3	9�u�i�J�α��7~_{�ϛ s��bg:T�O��������|>�<�z��klT��T<�3�n|�-��y���eh0�TF,���Έ8Z��-3�m{�̆�.4��s�_�|�=�o��fY�ωOP� �;�O�iBx��\2��W��P8��+�� �Lx'SN�\g9��g��*��gcSX���މx/j�c[�è�3��z�;$m��QɄ5��<�f����q/����(9C]�w<�>5�j�"`� lkiq��y�:ya�������W?F���X�6�Bo��H����f�K�o��Cm��2w`�x���%y��X�)Ol���ዷ!��䄯ϓj�Wc0�fYx]���c)?����}ǳ�*D�]⅂pZS�j/��o�^g��|N��u$���cml�h{���f���9�ye�'ko������ I��v����6�v�5� %_����^6~�����`$��_�|b��SyQ(�lҩ�'WLLFQ���8Oy��t&,�S���B���tR�L^nX�^��c�^���F��y=�G�I
��]��N����4n�4�s`kwZ3�dho�w8D$����QƴC�!��b�A�p����'�w�ҋ:@u�r��	U����������v���ﴇ���ֿy����˟p��s=v`�$w��r�S�/��9�:ͅ4w�v�{������@���w �4�0�|��rR��x��8|%�	��2�S�SRv���a֖�p�}��w�g��@0aC���������Gt�Q^d���o�Քᄯ`9�>�v�P���s�{�r��>?g㑍��5Ɯ9b�旳��p��s�<Ny�&����Qǃ��켰��� ���7}
��&�O��!f��8f'��_`Nt3���fy�|��T.�x�`gJE���V�����t/���/U/��v2>�fE.��h��2u$Ɣ'9�[��L��v��R�`��%��=�����Г�v�Ў���Bg����z��@�1V���x���R�C�0W�྇���Zh��}�W�NK���E&���NF���0l�~4��� �gUA]�V�gҹ��I�0�yOz�2��� *��MgꅷWdqZja�-p������Dk�h�3���u�Q�o�iO(bS���j�Ȝ������L����I����Q���)���%�`�)8r�9�}&�1dCU�kǶ5T��П�z%����u�8�����\}���:,
8�Yn�o<]��:g�������q�3���#}U�F��BƖ��G&PF�u�dQ����$ G�5���Sw�����vʋ �3�����$���@�x��*�'C��y��m?��ε^}<z��WLkx��PE�l<�qw�i7�s�K�f�;���m��u�}f[
=�]�x]�#��;^�2���V���.!�![eo٠�'+V��Ɇ=*;ki+�l2����Q��u+�ʙ����A�G	�0$)43k V�� �_&Ȗ�\�F�3G��D(��ܯ�-���4I< y�3�c�&BRζ�K_�c,��a'4OdF�>I�u\֦r��XY�+������))�cb��4Jc�>���|��c���Ce�:�#ڏ��ژ_5���U&�������i~�p^�O�������m��,��y�_�k6//��C�>dv����Ft��Y,3���
������R�Z,S!�������gSŧ:ِa-Bݩ�>�;�b+���Q�	#���0O�P�G��иnۚ�*�#�C���{ﶻ��Cw<5ʛ���p��1��Z�@�Ɔ|���Z�4�i��徜��S�������¯.)�_߼!��G9B1u�G�)�Cƿ��r�����͟�=������9�^��6��N5:��ۍ�6�h�*C�b�Tud
i�%ZXX�w� ���{�i��AM�������4&���;�R�}�����h��c�YY!?k��A�ڲ�T�«d.��E��_G�������8�{�:r���*�źə�#�"G�3�b]L�q��ȳ�� {��nR�#��[`K�H�ЛA�>_���$8�<e��p&���e��O'�o'�a4(�o�0�~�>�0�{�rgjdUec�ʨ�S����>�����v\�c�(��ý�>|�$�[yDoG���߉��^?����N\:�]ey�G�[7��������N�JĔUCjW$kZ�
g�hO�EE8i�J�����:�Mw09j����@�4c��j�ۉ5���Nc���B���`!������,��F1%����*�:�a��ծ�o���4�L	�����*����ûW<�#2b/�X����9Z��Gv���ƙ�3(�#m���M��{`	�F�V��d07Ɯ�2dJi�ت{:F7�}%3��pF%//L
�9���4���6l�^��3�B���ԑ}���zy24�sл%� (1~�2����l:_0{U^�0�M��(c;�G3��,��"�#�UR�䓘^�v�5�]� �8�ɽ��y�?�ݿ���`aa��"����=2:�+w{c�s������T~�w��l[1�	4�^j�ɡ�5=22�+��M�-��+���l����)	Y��YK�ʚT���m\��GL�A�X �	�j�z��{VwrTpx��>���p�f92���O#Li�P�S'�)_�A&z_�'���9��ߡ�����1zB�+�8K���:�l��sV�4i�����G������Y<�GyB�s�De�(B����B�I���yPH��a�=�+���T>���W�(I��HϸE�d.HIB���m�gI�Y���J��v:���Q���d:�ե,,��|�
9����E��lY�a����� ��.Mb�����AoMY=6�?�	��	9�:|�Q��]m�C�ѿB~W4d�8�[(��0�:ER29=IX��ds�a��5��`��UM<��W������*�h�i�s���U]�	��"O#�ueo�Y������qd�d��o���E1���~�Iw�YX��	ail�sU��t��t��rd����x�	�l�J�����f��c�twcq����jţ
�s�Kuf�Ѹ�G9w?�菍|�vp�JAne>����9��M�G�m����Ene{6C����J�b�W��Χ�?GGR
~ʓO�D�S�v�/9���-�"9/O�0)�I�����)C/��}0�/����t#���v�x�)�q��� �h�Wm��8�t��XS�ODoS�l�j9��'�y|���	��3���&o�7{�N����������¿�kc���8D���W�a��̬���%U������sh����>:o�\�����}@���^XX���9o�>��<k5`9���:���w��!��J*^k쳸r�G��{'G�,_���b+'��H�(�>��GHUf�;���E�XG�h>UX��f�Ɣ*O���^��|��^�:��:��F��O���0�A�pF�Z�m]٧e)���d�d\�)y�^�ì�_>��$s��>i�%�Q;�[�WMN^X�#h9y��;pΟ����c����7�?���Ů�Ü��,���������G���h����?�wL��zi==c��)x?��]6)8��X?����(7�R������bȋJJ�
��vl����*yXo�x�g�r�ٰ���u�y�[ݨ
� _8��:C_�T�[���~��<�y��}�n��;2�������3���pϬu݁�����I���2��IS��T\��o���$qd�׿I؃H5���UĊ�
~뽢U����2�x�~�YƲ\���n��#ݠ�k�f�'L�R�4}G�Y絇c���ax��n��2\>��<㈃��,}�Y1������5쯷�?�r���6*�{�S�W������m��5�yu�z���T������z�ĸ؏�/� >��hNX0y�gT"+K��|W�໅U���A֖��*�py�ض�b$2�r�'_�����-�?�ܨ�֊C4$k���	Q�[�9��E�/ϱ�mY��q�@$���hP��*�^���ӻ����]�6��>B�|-,,,���;:Fo��56��Nv1�,��z�Y�W坥��'�$��c�o_K0�;=e���9�xe��^�����i��LP�c] O?�k�|%rY8��]�B��F��Ix�G��t\�I�Z�}<���.��ꓜt,_���0�^�k*l�� :j}��z�ڡ���������G��G�UR������i��_Ǝ�r&��z�~4����eGag�+�f$߅���O�;Ǧ�ꔤ�������8��Q~�G�.c?�[��N�_��k��LQ���E��#S�����b6_�4!�4����K�a|�{l�E�q��h�drTr�1ת�&�������s���|F�Xb��=By�N)�9�2���'_�}���x�!�xx����L�����#�S�(���9⾵��C���Ze����W�::Z���3���^��*\�2ӳ����;J��S�T�ذ��!%ˮ�ܔ߉�a%}���J��Ѱ���^��hw��k�|F�Α�ʳ#��Δ�LwrOԵN����0��!������q~X����C�-���'�yc�g�<3p;(���1�K;'G�G�ǂP���Ũ}�����@1/y��� ��!~=d�����|a�&j�}포���4�|�ǫ��;vS*Ջ����{��~���Nw��,,,,X\/p��v��Avƅ�цd���'�Zo�?�Hš94F{�g?5J��ݎ���o;����3��:ƴP��B����~�[O�h��ݞ����s��'p��Χ�_ɟ8.��֑3��M��6���SI��%��S±�=�Dכ{��V�q�-�j�g���a�	�~w��D�3Yl�/�y<���y5�u���sl&��J䟠<W�u�3g5k����{��wy����V������jL�@�u���Gq�˜���p������p�K���Q�j{�s{���x���͕�r���^i=L9p��#�E�N�G�U�(7Q�~\�驌N�	y�/�&��ӛ�:���sX
�������թ�a���G��ٛ��b�9J����I��GG$�e����F�^�p�CRu��MI�/י#@1p���g6����ǡ[Q���8n4,b��Gue�� �a��݅&��t\�c(���5J�F�Pק֨ʮ�QI~֛�Q��Q��B�^�}�d��h��2�D%>T�ݻ�ܓwH7��Dͺu+=:x�o�eT���C:>ҷ��S�w
_���ՠ�x`�����H�C���{��S�sۧ��5;�.����p^5�<3or�q�T�2/�9�ٍ9v�R�&!�Jc����w_`|8F��S9��u���$��an�Ϸ�s���X���3t�x�FP�9��ȥHW�u�E�y�0L�/�pEI�-�)�hP�G���^�-z��r�88��0�}��n�h¤���35d�Cn��76]��T���Y~�a��'�&���{��C�1����g��0r��������G�� �(�:���0ܭK,�����Qȶ��28Pi��T�q�N�`Y^���/�B�z��� 3�_��L`#,�\� )Ӑ66"9[zOQ�t��%��>�z:G�i-����q����M�sdc�y��>� jg��ʵӝf���P3"����8r�e�#��X�CN#F۠��ka��*� ;�J9� ��q�����5�g�Z��l2l�V9l�nȇa�>�%s�>�qב�:a�rzaAߧ��^{��3�)�>�z�4�/��D��a�V��*%˘kV*ڴ���'B���zw~����8cȃ���y1m�KO�)�_�b���WS.��'v+|�<�=5��t��X�������ɣ�;�.@�a��<�s�;�gxK�A�5�nyv�3��E~��,���q��3��K"�ELV�.3�"�LJ�r�!r��r]�u���ҍE]���I�0,����g20G�x�H�-���Q�敃����g��-�a��m[L������C�(���;���N�{%j'j|�{����gA�	�o9.aaa�s@��~"�5/�u:�,.9pT;y�� ʮ�'���B�<%%3��T�y	���9����3��d��������n�V�^XX��0i�{�H{&_4��Gsn����ċ��o�6�c3��+`u���G6�A�\�k��6XPI���af�X�O��&�L�`C�6�φN�VF(ۍ� 酕:�Ô#,�W,G*�{;SN�ȧ�C]��-���E���j�I_;�ڡ�aPvuOL����ڤ[��x���*������P鵋�q>���/ڔl�V��F�Y�yΠKN9؁�ϲ:]�ݥ�C��8�Ef$��_��ɝ?��뉹�Ң�'�]��ߘ�~3F��w�T<����)O1�Jғ ���]8^w���U��f����	^����N 9�r4�C��x1i _}���
/�e��c��d�N-�'���*w�-��[bgn����N�Ml���c'̕}���������
�!�tG��}�zI9F�^��ȧ�	~^����>[莛�ә�Ua*�]��>��Ӏ�r�����*?�O�����[N4_XXX�M��M9=z����#����M�O���a��X;~�ǤL��Z[�:��7�xL4�;z��#x�Gf
���ك�jԔ�s�iӦ��Ǖ�~�c���O�����ى?ϧR�%��dl.��dq�0�����LC9�����-�D��K�;W��T}+r�e�T�R�F����b͠�'�x��=��Z�2E���	JI�D���TT_<����J�yW�V^�v����'gG���a-ٛ��Gu��y�d��h$%'o���y&�+Tp2��O<���R�˻�a�B����y�$(6ϻ���^���JAZ� �1�r��A*L`��q�zɶ��-|�?߿��Q`��,�:��x�3��TL��ģ�2��'�����B�|��7�{��g�Iuǉ���������#Mۮ��eŞ4c(9�1�fź�Lƞ����	[��e���޵�{B�ڥ�N&�8p�e^��W�y��W45��$ g�^Ò/�AxN(��_�S8O�5�����voa����5ֱ�xG��O�f���da2��}l��6m���*���S|Ż��:�m�������[��F��U�;�.�Q��n|��{GL|�MHp��4�ۨ�K�1������/aJ�}9b�Z[�C'}<�׃ބW8o�v��1�m�K�X]H���ͮ�{.��DX(�٭����(S�e�lbn�}A��&���:-d��������h,�0��L�<�Uw+	��W������k�W������VG�|h���ȉ�r���eJ6�_��D��S{Dp�*=
����Q?h�@4�%�
�Q_�NXİ��:3���L��z��u�r��ؐ�,�+ߤ��^����L����p�9��h$+�@~(��)��x6�dG3�G�8.b[FHNզ4�s��&%���6�/>������,Km��)��~��3� f�[XXX����	���N�j����(s��ّ��E�b�rr��.��;m�wA���H���Q��했*��i������}_	ȋ0䅜��`%�T�<��8��Q��Ϟ�aN^�0�L��
�t=N��3v~w�OO�N��h�煝֫�G����1�qO��= ���x�bX���~P'O�X�t�+z;�p;�P��g��͍@ن�ȿ�q��|�a���
����4t�ܺ����B����'p�h�{�G<����x����n7w2�V���?��A����:�H=��&�0���4�}�z�d��T;�"K2wO+Ư}H������� ���r`����2������q(����Y����@�I7��c(���_-���t<71R:�5��r�*�l�$N=e��n��dPj���:yp��L��N.��;�۸P���3#}���o��]��ceU��M����P�MFҹy9]�H���ya�z92��ܰ0ض��k��{&���jI9	���1���CZ��8�m����]��ht���UU\�t-c�ױ��ā��:7���_�=�����;zC/��m~~g�5�9%�y�n�JJ��p��+>�n�3GN�硹X��OÙ؋�X���m��+yP��2�aCqvl�W����\'}K�i	C���)����rD��:!��������n��Η꼺|�ǋ��%��-Fd��i�y������5�-Zy��\U�5ҡ��*'�,J�3b$��c�]�]��y�4^�-�<7_�	���u�gn�7f�N�faa���n�O����'j�U�7�V�|^�åW��(MM�JF�̼����r�'���f߅���[�]r����+C�O�.�����5{�p�B�D4z���ŞB�v����g� ��G4:++%a�t1*��Z�t�~R粓C�7�?[�U�V ��p%~���qǺ
���]��o�R�`:�C(#j��0Dk� Nw��dw�=�kk��F���ސϓ��ν�!��`�%���XTN��u���q��V����3�����1J���ŪxLD����]7сA�xE��8E��7�|�4�?�~�91vC>�����W��[���gn�<�RH��hO���$����_1'p6R��)�V�Sq&���'p`]��˫�;N�|V��!_�kr�f�Z\���l|V�5�0,�a|��(�j���m������+�̑��ÌC��oF��`�1^��0����Z�~�4���D�f �k�s࠲�Q���y&K&:�7LM���K�`�}c��J�Q,�U򾰰�~�.8ޏkT���~�6�	�$[��{ğ��U��"��kD����q���8N(&h�NzE�� 	�bX���2T]8*7�ʛ��*��n\��ڝ\�'�h�c�"'O�h.�։t��w6�?(4�n�#'�˖3<~X�Q.+�i�^���5�ݽ'�ֹ��&>��i��!�'��;��Zg۶殁����<�/���V]��f�N��>s����~�/��a���.,,,�a��9��1w�+Alļ8V�r�9���"|����cku)�@'I�p�o;�����9�y1(%5+���s2s/��a��(�0�N�9�כЍެ���]��t\����Ɏ���n����| ��F�Of��,wl���Qy5�兹m�2{�g`�t�?k�����q�{u�O����z�q����,,,,,\FCa��o���/��Q�ϛK�MHoR{bV�`��|K?u�6㭛�x
����*[����4Z�6Ǽ�Qv�����~"|�8x�Xcs�{/�<9z��$&�9�Y��E,@<��"> �J��$���Dk��Ǒ���G�@���[1ڑ���s^#;�G��]ha7�ߔ����%ꁖ�Xr$��+�LF�x�Z�rx�]�����(FǑ�a��f�g��k�4�	#����l��גO�SNK,���Mgd��:S�a�v?i�fX�ql��z߭h��G#�Xr'pl5Rr�Ŏwo�﫜�;�W���!U�ƥ�(����>��!��1%֞��dC_��r�{���=�7y�iaaa�`���TzdCu SY�k�J0�yJ秼d��s/�?�d���gQs��(!�|�eh�%O�����rZ� �BR�<���H�m2�����< ����5~��ԛ��	 �o��ҙO� -��/*gd�cK���Hj�����=����=�a�O�#x����"����{�(��z��r��I;�T�Q'��$���n��U'˕x�q�5�I�g��8�s���yyi�7��Ej	0�	�1-��rq?ZXXXX���9�	gfJs�Ƭqe������w��g8�3W�O�T��P��{�|����t��Id�h��4&I�fA|�&u4؋h��D_^XXX�P�Qͳ�������6�ܫ�&��rh�j�Ȣ=.����S0�B�ze�	f��UFZ'p�wx���:��@��4s��4��m�%e�[	���T�Q*�i�g��b8	UBe��OrM�q����9��FP�>��$�S�5�Z��^:��.r:�U���uҶ�����K�"<��i��2p�d��\ fv��h�<����窱��F^s)�+��W������"��";�s\�i��԰����¿�d�6s���Z�����4`V�B���������B��qC9�N�G���x>�y���fDd�+�~D&9��t1�+ U��e�hh������C��U�J��������ϸOW�?�S�WX�P�����Yy2�|�=�,��pX60o��,g"�����hq�f���kQ�pϡ�,�]c".:}���K%������uXel��)%i}�C t�6\;�C	p��yPT�ޝ�6MU�b9�X��q4y}aaa���|i��iF�!�d����8C����n�0&|�ᣅW.�V���,�%Rv%�!�mP6���(�5��<�2��6�<|C	���C�;�]GWf�v�:3�՞n��L�������/7��@X%��\���p3u�OO���5�({�[��|
B(�QOPQo0zU�4�B��=i�e���#�=��c��qGD��l�@p��w�w�q�q>k/,,,�N�:���:R2��V��zE
��g��lѓ13�h��Q{>m(�R=��T�
�G%�(��+���q��6	�l��,1�΃����z4�ku���ī��������{��0�4�TC���g�Ty�����W�<���LC�$@�Ҵ��h^]����qŖ3���*���B.,,,,��|��a>�0C^r��4��.�|G�d~�vw��h�>��~?�x��x�x��u;żW��
ޮ�+NC�J\����%W�#X�0}N�:r��]g|Z
H����q���j��v}#rmI�|�w�P���v��ly�����|�\��Ӷy:̫�����Զ6̑����L絭�Wm�!���(��P�l�q�{�@������y����ّ\Ƣ�L��&V+��������B�g<'�*w�k����Oܙv��S��{�g��cF^�6"�\#��k�1��E�=5_I�/
��|`�^��A⬁��r�@�<��D�r���Ԓ�/�:�4�t[�2����c�Y�/s���?{m;��V@�my��w�R���;t�W�V��,q��|�U2i��gaaaaa������R>g�u��IԚ~���7��<nD*<l<e���G7y��ޡ�n�6����q���_�w-,,�Cx�XEǔ4�Nj�����U������t
4B�B�0tq3�����^ڂ��=ϯ�y��Q�giI��%%|���A&~�P��9��M��ӌ�>��c�l'���!zT.$�r�w-r�!�?F��uy"��Q�;�C�i<�T��)'�y�������S�̶�sd!#Fr�:�j21�IX?{��'[1�v�^�^>�L�����g���z�����^>��6�ۜ�BWJ��!�p�x�z�����@k�Iy��5_���=�>Ws��C�&Q�픽�ϓ�����F���,����j�	�ֆݽ@��Q�#r��Jۙz�Æ�e��B��I�Y8���_
g⤏r͔#�t&<}ņzZ�yD??�E�d��<ݽf���E=��_��al[M��`�zmt�s�Z�U�q�6�(���ב1y���xUƱ~|Ns�錟q
M簒g|�S	��@��*��؀����������8�ݮ�������8�M�����ZD�O.?݃}R߶��J�����-��P{��B�HmC�hl�� [��'�5g��KEYXX�tx�ee��i4E��;{���_wBn��0�1p� ψ�1dxi1�����1�۩��C��H���Q1��*oȁ+m�_�X%=؂BՏ5�bX�<9������
`$S��(��Ͱ���ʽ�Γ}P>��v�������L��N�ȏ���6�a�|&�[�����s�y��o�h-�ر�u�FkAcd�j����|gea���1�Ѽwf�Tn�;VRL�%{v�XXXX�=�<���S�g�j~3��iB�n���kUdQTX٠�i��/�����rq2�&����h�<���8q���[N�^}6̣"��e��bm�' ��(�"��\HJ�9����}/��¡jK��y�S�rza&�fX��x�yCv�`Ww�>.'�5�ť:?�����wQ�U��v����_�~�?��!D�S���9zU��$!@�}��ߪ��Jd��ׂ#j>���Cs彻ⷯ�Sx����C:��,���z����wϓ-d�
�ó�o�vq�(�����&jz�A  ��:Lk�Γ�Զ�Kcc~�������).ϫ��_��z��;�����o��MǬ:=3+Z^e��8*�\-�OJF�F8l�;  ~>־R]&�3b��5M��(c��b�o�A�Wٓ��8��9}?X�'J:-s,����N"�L��j�C��U�������3��V��٭�˵4���x�U҄�,+O��U\'���\>~]M>~]�U�iVy&�1Q�2�כ�϶�S���,M�O��l��e�T��{T+ow��E�}j�Z�ߣg�Z�F餥c�z��=�~o  �î�=����ԯ��ʟ���X3��;����~�۷��p�^0��D��=��Xn��\y��r����]��)�.��x	}Z�'�W1�2���vGf�Ttw�Wa��.eX��4�c�f�l�gV�r]�&i�WU��=�6�zϞ�v_�_vi)ՐSk����/rU͖��#��в%�W��B���+�_���ɾ�:  �zx�z^�yUS���>�ｺ`z��_�8^�eK7��q�մ~y�  ���v��$O4b���fM��A>k���-8i�r�HG+{��x䎗������_6�D:�
g�+]H���r��X�ɜ\�-h�{�֜Z��V�Kx�,KS�C*�-IT�.w�ʴ"/�'9$�H��ϯ�'e0+�m��?��uJݺJ��/��V��`�e��4���k�l����pk;���  ����T~mV��&'��@uye:3��$[D�W!1���ਵ���M�������*H,��S�׷�B۲o*iY�<�a���awhyr�)�}���u{l�-����oE�Bv�6k�E[��f��+���qʹ�qW�  @?_f	X�����۲+��� ��l���ZYU
��-�3��ҩL�C�  �'������qf��Oj@�����U6��L���̔Q�=�ܵ���ƤY�H޽:b�>�K�Y�Pn'��l�c;���#�9�3*|��+�l$'�tReΰ�~Cs\�4���d`�ɴ(�S�f.��P�A�$I�L~]�y�:���*dȳ�*�Z�iu��	�{�u+�Z+O��|8����e�k��3ڏ�5j(��a)(7�X���loF��t]$m-�[\m�!7	  � ����Km��RE��屆<�a���f��'|��R�R�*����g&{%������/39�=[z'��!�1�x͢@)�pE7.oB�-uw
6��ש2��L�MR����ȗ�� ��}����nu�!{��W�Qiߴ�(OA��?�����-��ʩ<6��i��-��O�"�#��f�  ϵ���L:��9���Hf�&���q7&)r�:Z��]̿��r��u&�:�<}�F��1���  <G��~���=��慅��c�2�ٍ��GH��h'�YԶP���wy?�ok�M�d�6\��o� ��$1���Tr���m�,㎬́��U�Tm��r������Z�C��(�Zy�=d��jy�Ǭz�{6�:U>-��Ķ�.(�Y�kM�^����׭�n�i�_�V�P}<s���Z�.cl�:�{T��m19����:�r�MF�Hg�.ŷ����|HmteǞ�34P��G�=�_ �1Ⱦ�����Kݟ����g�tJֆ��i-��N'�Y�Sڔ�m-�ӣ tJb+]$[�]n���|p���R^����:��<��r�'ˇ�L�/�b��x^-��Vu��ʹ��g��~ݽ&s,O�}*׭�$��A�f���2-z�U�k�w�][G��qm��{�i���6W�rH�y{�5R���wݿpt��L�	��� U/P�Cx�C̛�y   a�
�> 9�[sM���7|��s���Um��*��|KiQ�X�B��ʫ­���>'���P2�B��C�:�  �F�0t_��V�R���ȡ�!��,�V�3lQ�.p��/K�B��V���d�s:d��?]��8^n�ސ�I�����Ӊ�S�Fɦs�ls�ߗ��߭p`�u�)?��&�i�ii�,כ�ʫ�Gɺ�_�ɮ�ߑ&��VS��W+��[���'�����<�hy�;�~=�?�t��ek�[4:���viylk;k���{k�m|^!ܖ������l@{U�>1��b/� ��p!@�����rQ�8���)gh�:���rG��w��5�]p ������-�5S��/ۜ��l�h0�X {R���m��3��+�^"�[	�)��F���j����5ۧa�h��}
/z+��O˦k�-Z���������	 m�\&����O{�o����X�X�a�2����L�'�?����=���М\�  0�����П��|>,��;8���f=��.D�TW�ȗ  ������΂�zF�G��_U"G[=å��Sf�JX�pt�D�-��-I)>c-P.�i�e��8�S0����wte��l�-g�-�4���DUq�҄CN�O������/�|�Y)ҲS����D���}��̮>/^	r�av_�4��{����<��i��܈�m�M ���V����m1�0*�ؖ^�� �Ǡ��nQb�JON���
c$�����jT��wk��!�@?����P�4�*
`���A��`cz�)������)���)����ۚ��8X_�MoVu��n�������>R!��j�Tl���#�A�������=K�2�H�������=/&�&�S���$�\�?�"ee��+� ���E��3&��   ~�E���^k~�[���༳Zc#E�{#��\1i���[]�  �:ߺ\^;�/�Q�Xq�:k0��.Ö]'>-�7�y�|�l����O��kDM3�bbV�N��
��CDG���w�a^=�5���KY��蘸����|�qQ��P��ze7dW~�~�#m�PM�/��V{^E1�ivo�R��B�����!��0��;�S�ڒ槉��t6 �O�u��,�  �۰��䂾�o�l�����R��1�D���A~o���3�������oio̤<�s�$�,'m����L4Pn�q�d�x��{~����u��*�oK7���j9�O��"�=OUv-�vGK�jZ���ݗfs��B>�N��_������X{P�^_'�$���H��߿f��n�<�^�òw���2   
�d̟̞�fvm�R�����.�m�8ӗ�SE�Ǖ&R�����3j���7  ²�g����k�V�{-����!�sk4�'��Άy|��9gU��'dqU�
e�N��%1�}��j3�X'>�f�%�L�g��{��,ʃ�$Sv���Un�p0[�:���r��6W�l~�v/'�N����hd��2�._,���o.���)y��|Mg�z�U#�'�����h�TV^��ζe�G���t���V�)˩�к���vz�Z��C�_�������  �پJ�8?(��O��<���)�O�<���z�:-A����:7�Z�4N��;o�78T�IJf]��_��Α�#�d�Y�,-���U0�x�-���M�E�5�#�c��^�;2��I�Ɖ벚�hw�MKv���]�![D���O���쭺]�wq_Y}�g�d��;��C�M�ˏ/&���-QYv��k�}Yk{d[��t�BG۶݋�c=��P�*j´>�w�  ��{�Ђ8ֱG��9����a���9�/�/I�O��1ܵ���#(I���K��}�����e �?���I�� ��B����k��bq�Rn�����m��z�+"����c�9��-�5��C$:N��8�z�V�����Am�S�yb�c����_��b��<p�s����3Q/ڀ<wX��FN0�H�d2�³ŎI����DZ�!U��V��Rv��m�n;e_M��'�˴���iٳ�D��t徨޷�����Y�]�C���߆��ݶ���_�C[�Gۃ�����UPd�|��4��d:���"I����wY�������  ��l�-zd�
��ls�������M��*�+߲�ܚ6��Q�T��qe�xC߻��L���-Xs�������U���Ry�-Ez��˘?U��\\7F�t����>HV�����x�Ʈ�����>����k�u�S�ϤaOe�)2�/-M�Of����j�Z�g�2u�� ���b��͠�Zҳ�{I�լR����l�5�H���&��f�,�m�uY���_�K��Rk���d�
�j}p��Hct�3���ɼ�v����� ��YjA���a��ɚ�������_¿�r�ɴ)G�P�^O��߼�/ص��N�6��'��G�q�:������vcƚr  ������=��+��
,��J�L/k��9�m��,��Z5�9kR�mܿ�]%J�Ӕۉ�Gk���L�E"�5��N[>�^D΢R�y~98l�����V��7��l�?&e�Ym�=s���[M2�:.�Y���?�X
��F��^5����J������<�OT݆������J��ng$h^�+�,{�����ձ+/+  <��}�8?�����4H�ڂ��G~��'H+�|+O	��
_�OW����y�j^�W�)�"f�Q_a-u�D�~���{y>�LM?�?��OP��L���׷l�'W�k��l�,Q�׊즒V�m�V�(i\�n{��{�n��C���u
M�'���O����=��O�?�m-0}�[휓���?뾦Vo�ll���'[�  �Td���i9��������o������,�"r��P�s�#Xi9AknT�   �!>w�O�D5ʈ�w�����t*泾���ןSj�<��"��kt��/1(���c����c���m;S����R�LY�yZ=��ί��7Ҵ��d^�Uvr�������=��������ݮ�iL[��Hm=���dK���k��2.iķ�������$3�  ��t:����R�� M>)Fs�i��ɴ=��*�{�W\!���^_�f�ד=C
�Jk�B@(��;/����R�c5={Ew7J^F�[\�ʓU�f+�d����2-u|�Mg�l���/Nꑽ�[f?e�V���Q����h�<�ƥw��� &ӧ��	� u�����3p����i  ���4�ΫI�f�a/�� �'���9�m�Ü󔋙���~k�*|ң �;X�9/.n�ʱ�f�?�?�ep�Ss��쥙��c�惇/nY����,��{��� Oˇ�m�,e1���{��������NQ��T
:�_ǜlE�i";^��24�o��i잹|�>�4����S���Ի<?�`�=��~��)OW��5�-V\}�F�T�@�c߰�F��S�t4�&������l �Q$�p� =@pt�yv�Ϻ���:�m�.�����֬����j��� i��bDݹ�ҙ�,8��4�]D>�LZ6�	�ƀ�~��l�8\'�%�͓V���V~�z6�n��Y�i�nK�o�>�fN��F���i���ii+��@�=��)�I�<+fl���F�3�JR��4�;(�����P�'EX4  �H�1���v�ѭz������a������Z�U��bZɝ��u��C�(�v+|#����u�%  �I����6O���+w����{���	sn�+)�(�Ƀ�1�#���5���"�=B�*�b�6�+�ч�w%7�c�/_-D�3�')��yhC^&8x����*�rGf�۲�+iE���fCi���9�ԧbM��Ӫc�_W�	e&�Wz��խ8�hu$�3��(�e^�3�j2��Z2�.�<ɑ��x)w�g���@k���ġݛcu�QV��"�le��]a�5���:��ܫ�������-j.��x�  �	)! ��g�5r]4���� 肂е�
)�~h�Y��|�����I�N��ڠ3�a�L�n��|`v�ym���C]���ʙױr/�x��Mzb��]�\�#�}�mmL/�v=����r��k�H7��!��R��j�����|2�C�Z^�]�>�|5�MG6�4-�ZZQ��}��A�Z%�b�l�}��[����ifJ5M�P=)� ��rr���Y{1����i����rF�N���]>�s�G��o  �������־Ґ�}�4����4���vY��7��g���۴��x
U��<WfM1�%z���9JJ��7  |7�8�����W$hPߡy�D�>�F�GЧ�*�:�o+�6TwX�=�����G��?�#��H3��w������-9<Vڬ#	�UĀ2����eI,�xЊ�\=��9WI�d��Wq�&�r]���h�=���4��*�(�;3���*ޕ�\���<J�(�)��)��*�Ta%������uƺ
e�,����m8y   ���f�/6V�(.0��Yf�� [���o��jw��T01���'\���jej`EJ�\����vMPΒ�<}�	r���u$uc
:J��~���͓�i���<_��k:x��Y6�:�5��v�i��m�iu�S靈l�&/Ԯ��^̈́i��[�y���B�YQҖ�l�<�c�d��좋bP6!E�j���M�%  |7�I�Ԋ�ڹs?��x���w��w޵�dz�b�ko
�س�X��o!�h�N|B��l����   |q��a�(Z�' \��#h�˙��ɪO�E�;)MqN�q��� Ǌc�<c+w0���F~sd�sgV��f?�wJ��0ZU�@�ꋼ�㯖�ɠ��F�h���������UҴ�-�X��)it\���u����>�ݘ⽐�Za��M~.s.��K�w����W8$��O*�����������  �SRJ�.en<S]�#�<�i����m�AD�C�o`O�W�zu�vn�?����4XV��R	�dK�If'#'�������1Ԓ��lnˈ��@u]��4�����앬Q^���d�a2P��MR�]�A�����J�7�d�鴴V�f����'��sz7+�)�O�ޫ���=��5���~�z��k������W��N�)  �����/zy��f���|'N|fl�B����	i�:;/��9�S�r��-��V  �-`�R��6�yO(�!9��1�;Je�0�{~sHr�Qt��5����<@,.����Ylw�m(R9���aU8CZ<ߚ�ye*i�ɡT`*��Ɂ~���(ǶdPd��:�HӮ�d7�����Øj�B�Rv%��E�6�k�-]�}��)LQw\7��f�IF/+�*C�]5qs����yS��M   :��3��Z����,�X�t&���d�H�<��z�mu�Y���&��/N������t�#�Z��_��F��[�6n��#&�$��+u���l����&Q���1��]�7B�^�I�}�{�M[��zl&+eg��ZyR�paa�u֭f�E��r�ߖ�Nz�<����Y�[�Z� �"�6&}%<��a��ńtc   ���M�)f���	Mk|64�V��ǅm��=TNn�͆�\  ��,d�3��!OFO��-�/k�3���~]:�������1��,jeR>�o����Yk�d�q���(�e��q�;&�@��JQ��fmv�:r�4�~��#{����O�u���{5c�����Ǫ,�{ǜ��<Y�Z�s�TD�6�۴��tH:�Rg��l@���M���3��`�e"�&̻���0�̍�  <���[K>�E���޸��9��?�J�����o��߁�٭x==[,��9�6v�Ҳs����Hp�WL��RV���.�'�&��L�=U����[�.��Sk��r���r*י�9�@�m�Ĵ�������6]��.�j����cb���"Oa�K�U�V����$�acp3���7tp��JA�2x�-�K\L����۰3;v[G�1ks86�� �_���7�����1����k���~�ʾ ��_�K��Я`��NQL���/E������{�Sykk�1  ����S�~j*R���Z\ʇ癷�����2� p��ڇu�S�;r>.$���c�s����d���g6�Yc�ߌ�Kӌ�%�?��G8��ے잣#)�0��P�V���[��S�#��c�$ߒ׆���TE2ORn���S��RU��\{�솴5cL��i��Z��r"�2h��L�ܤ��Z����*��J�&����/K�so,׋}D�P�m/ri䳝�)X����o�BE�`#��Ϙ�$�4k{�B� ��Y��q<�������\���v�:������י����zC�����x̅"H���Ԙz�^p�}zDХf;�����\O��?���a6���4n���-}�b�D=��T�X��>��>/۔��rH>�uS��t]~]vǊN�p��2�^Gid��*�q��W�:י&��/ͦkɐ�&��^�&iܗ���-˨�n��V��^Fjc�ɘ4���s�߁��=�c�c&���mK��K��O+(���l;εs��*�*��߆�+M=��������'���҉���e������~�]�6�;zX �u�Vc\"�-�}��鸡��}��*��O�O}�q���֖�x]%m�p�����B'���y6.h�n�sm0jF���  oD3��4*��ɼM;�э�V}�^�Ϫqܚ�,x"8osqG�M1o�=�SG�,�-��(�	��1X��w��m񘢣�1����f���4UE)ю���Ms�OMv�ף&_K���^�ͪ2��{K>�ٶ�C���	�c%�d���� Levްr�7�����   ;�8o�i���z���G�}�ƹ�={ja�<H�$��'��b�p�)�,,t�q)P��U������K��_��f�б�����M;M��z?��f�4�-��ʰ��S�Y���⦭Ր]�P<{����T~e��|*��w�tb��%ew�'ٕ�e�|�L��;���rY�f�<Vm�"�v �3��~�9Q�n�{�D�Ql��ߟ�`iZ˜V;��#���)�  ����isg�q~Z�D�
7N���Qz�ug������F9�_,ܴK��f�i��sn��
B����V��]�.�Y�X����(�H>��͆RgJ1πv]v/��M�LGZUvWޟVޚ�F�#���݃t�ȿ�2��̞u�#Ӕ��<�z�2�m.]�8��׋��
��Q�L |��g�L�!��J<���\4RjN����y�[+�c#�͎��P~<���
�n�1��{���1��=+p0���8SK�I��O��.���K����Y9�=`��N{���ɮ�'�j���)e�ו���j׽v�S���n%2n2UOH�>:�����U<���B�"��C��c2߅l;���   g�c�]g}��P,�!O���ؘ����_2�~N�h��^!  �~�&;���l���a}����#��	i��{����-��j�)~�y}���
K����$u\nM��4�-|ϗ�&��8��L�j�JŬ\�����tn�:��f��l#�(G�)e`�u��-���JZ�|�r��_�u5'�*;�wS��J��_Hv�'dN��W����匿����O-�;k �,�HXF���;\O�R���g��?齦�Xڇ�^=b�l=��}�<f،�01���PH�e�l3����f���>���Pt��2S(-�`!���J��6��]˞��ݙn,��/��<;m�=�J.Ķ�:"���,kl�9�����B��N�v���D�3l���Qs�  @�j�ׂ\�69Z����]\�{�����[��Q��Ǳa�g}�2�  �6�fv�z���[[�O����14��_�u������d���t]���׫<�ϕ�amŹ(��������A���L������[�X�T2�Q�Nτ��yVx�B�4��X_��>eC��蛍����4�yUUҊ`'^�(ǵ�X^�&���#[.�Hˮ��J���M���JS�V:4���ɐ� =0�rE�+HS,>g���5�[^��s�G��[�ڳ;�*���{U����c�/{���:ڞ��R��g[Lk�/�d����������#�  �M���?]�M;2����'\/������'өg�����|��כ��e�e��3��+�O�����4F�R�Ez��^	'�Sb�8ӏ�R��W�_ʊ�R�-�z6hO�jK�/��-
�Ĥr�4.��LI�d?X�-���4��u_1i�nw�>J�6�F�[�aٻbYZ^���dyT�5?F�~����;�jpژ�v
m�Y���Dˍ  ���q�X4��&{el�2��+;?�� 9h�ݖàK��
�耝RsY��9�  l#�A[�o������-���6�g�	�&?��A�r^�p�?�&�L�_��Ǌ�g��ӊy�ȱi�
��S��n�HB�[��ŴJ����ʂ%B��1����K��²cV�҄�B.E��T哲���d��'��K�3�3���z����-�S��bEv~�>��z��;�����0��>ҵ6��tյ�#w���� � �)x��C'� ��_>�O�o����]�}��ٺMM��L���`�e\T�-�(�4s�R�.������>���!'����	�`�Gq76�]���饔�b�dA�	Kˎ)����i�X�F�j�&CK�-���{��R��i;�떽%��S-O^��^���|iW�;Ț����2�P�|*?���)���>��,�c�0u�  <��;e����!f��B��]>� vn�����=E�i�1�  ��4&��2�L7Y�}P���~bk0��>����T�ͩ�˽Z�o�b�HR�)�D�Yi��һ�\8I�YN|f����ڠ�zOՠ�������M��b�h�[^�X��+}�zk�mG9��5dh]�*��^��y����U�:����ߠ�nq����" ͌��u  ���{	އ��@{t��|㊯���c,���aoc��p�N6��߇Ȉ�;�O�◤�?�q�")�G���x6��ث�w����y�d��Г�fO����W�q�f��\����fj=g~��/W�d�vÑ8x��쮫�}�	+p؟]�  ����_cW ����v������e��Z9�p��廊���!��+ �n4���<4ߎ;����jK7��^�}��#N�Z��NH9%g	��Yc�*Z���U]���i�}�c٭A���1o�Z3<����1�����EoS:2�SΚt����NM�k8V�&_M�Z^�|<O��L�Ҋ<�{u��ƚ��5�,�����&{���.���}yl��;�=�"Qa�
O����O�����=ǛL��OS+V  �	o����ę�G#_�+��1�YV���9P}2�
�3�p�I�k�^d�lR�j�+���Cz�!�9�g<���m��D�f
�bi3E]�g��0�ﬢG;���Ѿ��M���f���J��W5Mʷ���#m��MgW�ɧ�[v�ݙ���7B��ݦ=�����{S�v�6��b��*�`]�M�~  �W�[��<�=y*;8�>��Lx����F����lS���j�+�J��H��jE�,��  �fF�e�	]���Hs~�,����kn�c�S���ҟL���ܠ���,]�.��ژƶ����Џ�O�j��i�-�,&8�H��j�.���Y�Y����d��ZyF9VK���L>.��H��Tg�i��ʷr���Z�vCZ�}�e�w[�IyU��HR~0��\Z{8k3ʞ�`k;����P���Ѩ+aC���Z:���c�*-8  ��on�ɭo�A<?�<���#?ۏ�8��1o��kq#�w��r��z�1�`6�c�+!J6�a��ÿ�� u��+�-B�gp#"��D�&.�:��� �Z�<��*R��6�IQ'n�>����e��zm����<)_E���Lg��gU����׭~_�����/���Z�Q���`�^ꥵ"�IuKk4��  �Zh%&�W����d�QAfͣ{Q�o��0�B~��U���ջ�0�J��AhȀ���^[�c>��&  �j�A�=m�Cn	V���ʹ-S��<h/�6��}��� �U���Y���3��4�������w���=�&r�6�����[ç���R��e��?a����X��y����Ǘ�ɸ3�菾�C\Nە��K��o�Ҹ5��ׇ<�����@'�z�:�.���iN|ji�:꬏H�YHL.{V��&O�_���?���r�hm���8�����bZ JMv:g'_&��)\��
�g�#���?[�����L�:����ɬ��  ���0~�ŧ�!]U���	v��I�[e���]�ޒz#�m���̹ð��1->�Y��?6�|4Lj����"]�������i�VZ�镫Pͪ�3�'\����,/�1��xϦ��T$��d3���Lie�XvOI�\?���l�Fy�l����t��ݒ�菤eqT��6�Lgڊ]�O�i�i�+�\�ܸЯ+��(iE����֣߂f?��6|q���}ټ��1���u1K���� �SoAvO�IO�/ӚV�ҩ�w�O������DG�{�[�E��"zw�}͉�O���5  �ip_[�R��+p,�4
����Sl�2��C�����x�9�M���&'wB�ԫr�F��Fyag~*'J=�&9[�r4�S��O�K�(�dL��4��tb�J~��+/�e�SI�f�M��4WK�����i6�mK�j��r���Bͬ)����+�+�HGj���Ѯ-TNm���4�f  ���Ƭ�ԃ kC���O�B�~��Ǌ���>��z<c��L?K���2E�N.�<��8V�(t�g6S�=��)^TǶL�.�E�ŕ:�}k��|��}��S�^��J�|[&�b���m�WxZv����W!�J�u����z찙���T3 ��d�k�OU�V��oK0b+٧��N�vlL�H��*��   �o5�d�*�QW�B�S1��+���c��W7���U�8�K�)��ڋ���	  �a,�l��3ˈo���g�]�9�B�?.;?}�����1���i6��_����҃N�+�S�#uTk2G���D�^���4Q%Y�m�E�+�ː9@���J[��+�Ć4�ȗ�UK>~|�W�;4c�O��n�]��A��;u�)��u췾~�9����8	4���� ��-�F�/q@V�̡2�~��P�'(���r�VqA��U�U�E�� �5@�M�)3ݾeO�3H�%���vM7��d�z<�l���z=�7���m�VZ���i��o������D��y�9��FYs�+�,�\�=��Π�jk�Q[1������l� �u��r:��F�-�@;���8��G>r   ?�l�Oa)Ə�z:Ȝ�'|�Wg°��R��;�}{�3����G��Ԗ�eg�,ʂ�I+pԪ8�}�<!?��� ˝H�j�d�B�c�Iv�x�������T瞩W[+-��cUK3{�,�x[Ժ-��4���Aʢ�C?���S�����	���JG�[9QYgq�٭%j�َ�nz��}o^Oxo `�Y��r�Һ�0�����2�c���6��}�i��i�����h����IͶ�O!��D(��F�����K�-�B���qv��awl���U5�F����հ��l~�G�"^�"_,��_�N�����E��̾�Z9F�_徤}��pc�-�h)U�l�2b��V6}C0�Q   �z��}^�^�M��T ��P�!4��|ؒ+˫3PY��  �_;�q��Џ3�ܱ~ w�}h2��O��gKY�v�ε�f�����1&�Y�N���ryR9����'�?�!�;�GI��3������<�l<�7����-�������[*�&w����L�Z�WҴ�24�+i��ӝ&�ۜ�SQ?��HO9���=�u�<M�a�}݀�ڳD�Z��6�x�A�ډ!�~�����OH�LZA���p��]v~?R��Ϟ���y�  p���3������op�?v��gx���aO��&Y�\�"�e~�d�H샷�ދ6�z�3��N\:���b��f�j�J���e[=f�#��_���c����mR� �װ��s��̒K����6���um)�k���p�&��6�E���t�	5D�s��+������e���+���!?��s?���+?&��V����s�q���*xg�  x7.���{$���I{�+r��)S{\��l�3*�#��w��FQ���  ��XV���נ,��&ui���Nw����JҖ"֖(W�q��\���f�q�3������;�ɭ����S�Y��y��"�Yrp��o�YhrF�eǤCMsw�W�P�9t�;��y��ąR>h������ٚ&eߜ��C�������+��Z���|��e9yy���h��_�����e{l_��'T/s�Qz�v]�M  �Ã�v*ʙ�|�Q�u�O�}���I.0�m���Rd(?vJy� ㄶ��ŔӤژ&mm�`�н�d�8�~=�,p���DD9Qg%�b��tq�>[���v�\š��v�ͯ�4�/��U펖|;Ӻ�"��S�Θ�=��=S9ֲ!�"�i��w�e߬�>�����&iY}�gu���7�gd�yO6%��+   Ёs,`|��Qj&=����J��$(�:���[�(��O(#>st.1A� �'A����pCإA�=}�Ɇ�t�]ɚc��/�L9��ɩH�]���sN}��N6dpO�eyGG�a�����g��bI��j�T��}��pt��҉Z�Gi��JǉO-M��ʷ��&�H���3�����^�w��v�{���jidP}��)�Wqȶ+��u�9��<�I?H  x*|���v*|�S��f��gN%ו��	h[�͜5P�jɉ�.;�R�E����d,��qi��*lf$���`��y�K?LH���ua��R�t�wU��Y��j^J�R�>b�ԆdPIUvy��s���v_��I����2���>�-�w����X�\	��\��U��e   @�5�d��2)��ݢ]�ɟ
� �h��0X���)��M/5   ���N[uX3~沍+�_���c^8J"U��A��GC����%Gg�&Ql�r�?��o1Ȁ�(&sfY����d��f�J��9O�2�<YQN��k8@���v]+�BYZ��
8~�<_�'�Ӛ|��\��B��ˢb���-�3Ծ��V�8T�I�.}��s+��� �`zf]���c�'�.8�2|�
�<���l��}ș���J���d��B��܎u��E.�G�������S�B	���y�~^���k�yV|���0�G��q��i�rdZ�&�k��vc��Mg�����,Oq�&{Q�ؚ��w��V�kiO��  �ב�l��w�L Ǣ�Ƙs���  ���/����H����\\��]n������Tg|��,��%W�����+Ău��&W18nI���c���$#-s��óg�Kۅ�Iu��>r|V�+�:�U����^x��\'�~{)���V���^M3yZ�|��峯��RvC�����b���eCv�{J�s �Vnh���A)�<佮_�.�=�fK���ooc3�ɔE���Y����]�!�9�	u6�{�l���t�����>�@����E�y��>+vQ�^��.j�ײ��������%{�gyX�#Y�R>��UꊿO5;F��9v�.���W���z�٭   ���e�暽�� �i�ϫK��EZ��I��byucL�Ñ�:�ؠ�+Y�(s   ��	������>��sحY��9S�����0Z�2��Rļ�ӧ����3��Z�ӳ.��Qt�����oEy�Yn�}��}�ns�c��ӏ�r
/U���O�(�SQ�j��L~>��ϫ�ֺ.�1�`��r_�n+i=��cZ��F�gy��
�jC����6��ǥ�S�~�Y��Xk����P�>��W���������1|�{�q��
l�[�Y ��q�������稽G\�i�?÷O��1V���+����3o�2���X.�l<7�2��Cr���s��~>#~w0�]L>�I���I�F��;)�=>��^1t� �7�,����*�2�2:+ٚBm���^�l
a�hv�}���^��"�"�Ҳa4[��ֲ����E�f*V�٣��Ώo�WV��M�����Z=F�I�5[h���i7@�u  �j�e��c����k��L,��d�l�o�0)UIa�\��EJI�k���	EEj0Ȭ5P�  �Y��;�:�[��]���5�P^��$��2��V�`tᬌ�'��ך+�iI�`Y�Yh�����/�ƈY���Z���{Pg�uZ�L�bH��D�,GK�k׭՟1����h~�� l�i2h�C��Q��Wm����|�� ���q�A���~m_)|�ިu��:�����1��ric�\��&��&������G{��c�Z��!��V�0)�5��ǆ���u\^ _�AMk�S�r]���1���A�[펖͔�@m��&C�f���9�[_�]��{�-<e0�5��  �K�{��,��������m�@K�'k
��-T��;�Wq�r��H˨   �± ;�r��#h��X����B�����;G��l�-��-:@�V���4�g����/�=����"g�r+&WT�S�w�5�n�yȜ���Ҕ�k��%�ZM�� 몧��C-�iF���R��K�L�k��Zy���_��"~������  ~������a�k^G����훝�='k⊃6���M[�,ʼr�6:�En��h�л��cbFYQ�w������o���m���m!mS�i�l�����������c����.j�(�/�3ً��VFI����8�Ƙ�L��   �NM���Nq�Ŕ�o�y�
਱ϰ:?>�id�p�s  ��X:{�^�{GNαm69P���e�`ں���J�E.80���s�������-�))�#:8�9�J�T*�D���q��wG��e4y��jR���i6�̓�T+�)^��T����6�gj2(u��YS�wQG�uY�x���.��L��̫�+�n���X�ۭ����A0  x����}���<��:'��5xuV����Jm�+ۤ��}�-����� ����g״�  ��IDAT}5)�^�)[I���r.��dc�{IrVu����Oq�G�����JZ�f2z9��X]�{�v������f��\~Z�@T���7��G��ۇ��g+[��W  �y�߶q����q�5���8\�J�+0�y�Eq���.�$����;�&���e�>i�w�W�VT  ~ �����^#W� GWt��~��>y��{���d���og�^�����Bϧ�}��
>�����g��@&�	�3�g��]LOY�H��ɝr����d�P���RIk]���id0���������oPq�g�X뺭��QǠ�~_���Ώ�5�Z�I�Z��8��/��IE���LI��|�޻P�w�`  <��j�B�e�Vҙ�����9�i����SW"�����=mK�Q���j�K�¥(���	[�#|2��-��+._�ûC-���/�fr!Ve-m��SeEe�a��_M�u�?W��H��ciW�L-�V��U�Τץ�U�do�7[�FS��7^�F��J/է��   @��<M]}�7�̱9���o�ͪ�h̺�<�i1����aD�
����KN��ə��: ��Y�?�Wఆ�����|@�d&C�����0���h�mg��B�^��sK����,��� �I�(Ntx�Bq�?��I�H������%qr�U�`�(��\�l��CK�8�����ۍ��Zu��_%m)��i�3)�c��Z���y����[��ZG�*#�<@B���Ҟ2����րI��\��>�s+�Ub3%J��C��sT�?�#�7Ҋ: �_��x�+��c�7���q��3���5�3��϶`ŧr�
����b)��w�����P�Yd���a�Ja���A�f�
d�p{�$]�m'M�\7NB*��[V��U�6��>ݯ��y#�����Hk�L+z�V�H�m��}iu�c�h�E}��Lj�2Kc�h���	#�<�8c�m���1{�0���    ��Ӣ����ik���~v�]+p��V��̾ua��<Ł򞕻��Am^Zo  ����|�~@�����0V�9�(�N�踴l �y�؀+w�i8�IK"G��rƹ�� �(G��r/w�ێ�[�X�u��%n=i�,!��q��iI�[�)�eV�K�F��7��4S>�"�)i�@�����,�󿐚Ə�4�� ���m��V�0�}��z  `���3�g� ��u��o������s���|�޹�x=��>i��޻��;&ì��>���\�%{��g�6+*�;�x����S�+���h�6�0-���fR��Ǧ�b���J��m&�uB�X�}���NȠ�k�uo�������=  8���ӭ4��-T��L��?K`�H�?��
  ��2��f2�2_���Q2� ��^%x��r<?f���z,I�;�©R;I�eY�N�r�6�ɯ����#d�N>*^�8�Z3�2G�1Y H5ͤ��;c���˪5w0���IsB���R>Ӓ��ɇnٟR>�.U�+��(i�X�o�y�px:%M�_v����� �+�Ճ���.����,�8����V  �%��iY��WM�<_T�u-����d�͵�n��g�.���쓨��5N�&̈�(R��.�d�=��#t�L/z�Z�S��tci�rdZ��+��f?T�:5�@�EY^�H��춊|-�[6]�R���J�n]�G�8���U>��=��;��8~�  ` ��|;��X|�~k�/�y';8���,9�i���(di؅dڔ���Xr��sި�H  ���O���@���B3|V]<uG������oԇ��q��p�g��t�/���U
_N�d�|m�+�gI�e�q�r���FU>�����$��]�����Ea����<�xv]��t�<��Q��uTgQ>�]gx�.���ъ&��h��P�+ӭ\����ĝ�P}���(Y��a�9Y]e�2�q'6���̨>қ�x��Ub�eugL�{"��`N��~�6'O��6��j�Ůr��o,�,~8ɥa����� �o�/!�L�/����64�e��1C���c��m��M��/�v1�;^3�4�3꺤G]�[ƙ��%#�ܞu�2�>ʐ�XZ9�4ߨCZ��a�w��tX��+�3�9)����䘗:8�S�&�5E�D��S9R�_�;�7<*���fO��f�\�Ci[�c�0����(�����h�W���SOuMvUnǻ��1���{Mr���'[5זkH.;{��I�}${]��q�5;�H�׳b�����w  ��6�7�h�&�+}�� ��z>L%�Dy-����� ��h���S*3V\Ɍ
o��P�fg�<�y%����P�|��  ��k2���5�_��d��w5K��/O�f��N�����=���J�>ȉ�Μ�l���	e��UX�r~,;��a#Y����L#���LGr��<x��)�Ι�ڎ����Ë���s�ipJ>����޽��d3R���8����'=�,���C{�s�������{�4������x�f����}�$+��"����?>��D���L~Zx'�;L�G6��wZ�291i���N�W��J��F���lh��7�R����}>�O4���vM֦�zx{gͿ����	��Or=<8���� �r�p�s�O����X*�+���[�P�s^�^�Z�GP�u���9���y/��ް���]�R#�<ҧ��Urԣ)���������Yq>�SYQ״EYA0.dn��������fz6�g~��/��M�x�&�Sf?p�&��=UL���>e>)8C�
��#�pυ�aR��ݑ��\V��,�T-�˚=�ȇ�ﶰU�,�QG���@��β6N����6�1��Z���������1�<Ph,N���z����3<���G�kwO`���7Cq�����  �=�1��H}��/�5�ۯ�1������c~��+p8[(E�s2;w��3�U\�{����X��ėy���,  �5� [+���zrg+?ű<M<ǆ5K��>��s�6�s�j�k�Q��sz�J��{�2=��U^�:|��K`2

o�k/�w���g�=fF7���L�}��|�nz�g��4�q��� ����J:��cC��?s�O��s�/V�1���JU쌝��uD�U6�k�TW2����=��<��5�z�^��4�S��(N���δ�[{G����)� �k�g�d��O�m�  ���>e����0�k�\��
�}Q/���(���*O�x�L  p��˗=�*��5K�y_���>�}��4���� ���AGE�NH3,�.{���w  ��N�~6��-�N��g��oŜ��`�3�1>7�>�����7��L���9���#0   x3�x��^�H��}˗�[��kK�1Q�
OX�8��.)J�x�A*�ǧ�  �v���b�3�t	;�E,���?��wP����n�bq��̳�2ch��2��Zy�L=�����;�ku�|�{c�L��.}q.;   �	,Ψ\������K�a'K.������!�3�:ÿ�Réݻ�N@g�g����Z>#��ϖ� ���[   �#^>?������@3/��\�����l���UE8FԻ,��1���7dh�2��/�  ��2��ߛ�����s���Z�H&�@���@�+�������>�I��N�����^�C��N��g��*���F-����vM�2�k�2G��2k�nt�Uξw𺪝��I�w3;�/��Lg�  �YY����XV�[�M~�_����WL��;0���&���$�VO���g��F�MϤ��U?��p;�g;��vl��1jeKy�l!��^�<gT�{豹�f{�b��r~��zG �Y� ����@w_�������&{�Ʈ �4s��>��qjr��f,�*��b��`���~�P��2�����=G�A� �[H[�lX}#~�A���ux\c���s�g_YO7�epZ��kA��yνN���y#�C:㾡~�� ��V���I͹&J�w��n �z'���9�e�ؒ�O=��/^����!�ch���8��������Ě�Mp���w��{!�9�����J����_�i��>YԨm���8s�=����͚���   E9�麶��O���?�c��_M^es ��=�/�2`�g�,s�@�7Z  �D�]�7���Z��l�mP�W|���V�6��i��[��#8R�ZpG�s�X��k�쑣UFOڞ�Z+���o�Ay�����:-�}�O  ���sz��������o6��б��
�6i�}�0F�_���*=:�(���^�kO���2�Ҷ�c[d��N��p��kio���a��  xW�b�G���kV�h�p�8�̢h��y�-�  �7����l���06cc��8L� �     �2�{� ^�-�AD3S�����%�g��{���UQ^ſ[��r`�q  �rB��X8���]��8�<*�2���g���  ��1�X��2av�bl�YVow�?Ug�Y8 ���}�G���V���҆��uUl��|К�~���  ֩uC��0S���v�H{U5�5&�m{p��5� �3���5��m7϶W����Y��hvQ{  ���^��o{G ��Z��?E�g3��>Iڅ
3o�p��7�~�;	���o   G�4t���3�k�̩cm�[=nգO���*wH�a�־���3�e�[� �Q��O�s�2��=^Y�l�z�'�oyo��O���`��	�5R�]k�m�tS��Λ�S�D˸�� ��@ͻ}���E�5�G�l��4��&76>=�C�l�r��;��� *}�	Y��zNL_P��k'|YB���s�F�+�C�J`�7�3�.��4��[���'����]�ЙT�k  ��Zdkު�/�K�|�%�چE��{T��٫+D?an\��Hi�?�䠗���� \�a�,�3�@M����ӕ3  x>4���T��*粆1��9[y$']
a�Bj�w�7w�h׶�[�A��Ӧv�V.t���yf�+e��_͕3CG��9�>��Y��U��l�^��(�˞���e �;I:�a#a�.7������ �+aC���K�̉�d[�� tiX�m}&��������kvK�N��n��>=�,�l����3ʖH��;8Oz
�n�  �$�6o�:��/z�'�㘟ٶ~_ �K]���M%c���^�-�A�s��uaV  ����k�v)v�)_Ea�G=ū	3�)�t�ڶ0{�n�ҡ���e'��pt^N�3�u�~�DTU��Z�1�X  �-�5أ���O��1����y�`�ݲ_Z�w�uԑ��ZOb�~�u  ����ӆYOa�#�¾ ��-�`)4>t��\K�0P  ���-��RƗF���|.�Wh�e�����-�ϴ�_[��>z�j��Ske��_˻%O�>xy�0cj$W�±�Q�<�3����  \��>���.}$?kp �'[�ୋ&�'Ы�^�U?����V�c?��J=eԮ�j+�s~_�<�2���c-�hٷ�@�?h�v�ie��?��
џ @�ʘm�����B%��K�i8Wq�|���E�J����58�$  \�o�������oςA9�gϼQfpG�n��06�H����[�K�y�M��Ϥb`Q����P�  �����o��Ǥl�7�5@����L���)�E   ��%��v��7㘽�#u   *0���KMq�����*��5/�(k�*+'��Q��1/���v�����Rg��7��  �H����ذ���.��%�X��f��YG�}tW��ל"{%�:���<9�\+���=��ʞ9�~������U�zx��n?���e����Ȩ��|>��쾷!MY��X�S?����zC_  ��4�6lc�[�O���]�#����t��|���7<^�`�+��g�u#u�=�����J��,jm^�}8�n���?�%������>/�%}a���dRy�Ի�Ň x������p�VN]�@������S�^�
D�W�o�*jQϦXt��82��=���+ �737������h)�{��򆫥��������p��kdY#W|x��l+g���|��y;�¶���꠷  �����"S�E����P��M���@O���j�����||r�s~|�اȔK  �^�>��9�e���%2 ��c�?���+�3➥� �y�ŗ��"SZ#nsuJcH-��LM)�O���h�5	�1*�ܾ���z�Nۻ���� ��F\]�kH6̨��[���t֧� q��-j�R��8g�ݿCK�;�i�.   �	���_�������&_��^V;q��V<�c�uk;�+  ܈��Ǿ���6����YvND�Y�,=�׻�b���8�����S�I�(_�`��s��˲V��>C��6����l�H  �(�{�Ea�M.��&?�yNo����}>p�Þ�����msV��o#~�'V�۰R�_��?��M  �΅�)--k�j���Z_�u��)|�}�N7w���mN?��MKUV��<~o ��7F+?'�  ���q��a=�p�����7��D�o�1>ϰ6�^���V�.���=�ܡ���{��%���s]�|?���G�-�$.�υ���	t,km�t(#=3�d��NS�S�z����� AwJ	  ��8�,m���������'��[���f{c��?ws������s�!��9�!�wz���Ȳ��4M����45_�&�<����,�I�Io~_h;�g�Ç}�ļ��	���q0NE��2����ue����Э .�)~Ä�v�����'���O��*.���]D�(��fl]�[����0�� 1��\ �/CAs�<���>:����~O��%��=���6�\&�y���T넂�x�k��{��Be���x*�U��[��<  x� �I��q�\��s0�l����p�a�l�ۡ[=`�g�6��iɢ�#˂���<iu@�C��?��r7�
 �H�囶�K���*k��	ZWQ��mm�� ��_�q9��Ƞ=�$1{���w�R  ��ЪK���qJ9��1pV  �Ph����-T�[�>���:X  �&���|@s�
mK���}$8��U ��y�cW���io  ܊�{���*��7^�+pta���֥=rNRFl(��A��-   �;#��F����  C�SWd��<6�8�\֖��͑�ri   ,�mT�3����e��l�F�!�y��ȳ�ڊ p�[��  �,�`���+l�xo�D'�;}&埜�s��Z��I�  ����;5�8������}��+>�1 h��F�)9:[y���\
<��ڹ�(b����t�\^�n�E ��9i#,e�F���1�x�L6M,ry��!T�h�{![�	jG���=��`�|o|�c�~�`#?Te1��  ����̠���A�*�� o�M�t /O���4{-��2}�Y���9  �6֙�m+�Y�g4�h�<>&��a����v5�>� ���M����v�gL�ϭmw��`�+p,9�]G��s����+�|xx̛��ww��3�  �dilϛ�c���q��h}8����M�M�,m�A�uD���<�¯����~�{���޺��_��d�]�����?��ȕ�{ �?v��B�h��ي����4�:��;[��jq��gt~�C�o:y �7pxkh�ˍ�mu���^�U  TF�h��d�Zp�Ө�x��W;geٜ��m��YB5���t�-  �*�ȋ_���+˹�C0��7r��У���3B��{�#����
���3������=7 �wX�2�ǥ��Uܪ5l��g�q�论K�{k�Z-  ���m��O�\oLXv��6M�Y����V���>����w}�ִ���hz�Ґ���=�b��jp �:  �a�C(�
+����g���
��3 ף��1"Ϸ�?��t   ����o��V�v�%��z��u>�s�$�L>�d  0�d��ֵ����!n,��d6�*oU+ȱ�w��_���?miU9k��YD{x�̜':ϸL�r�3ػ|1��Z�ˉ[d��������ZQ��k��  p/i�^�WNRf��~Ȳ���w�����%�Ӏ;@����l�'!}
Gd���W1�.����  ���p��"ʽ��h���8����� ���u�^јB0ħk�'O���1*����2��7��h�j   #p!�2���Sy���84?n�������4�$��|���̽��|���/i����ӑ�O�>���iJ��W�7ju����w���5��:���(�m��-�\^�V�{eړ�4� �s����P���Ė�mq\�JC�b����g_�2&�cϽ�E-9���7��f�d>��L`{��6�� �W�4��u,����Ȝ���V��7M�Q>,�ɬ��6x�R�o�M�}�3�or���K?yO&�G֣�FO���l|����g��� �(��<��6�c�i�-{�_�W�<�^h��[i�s��b���	���Sk[�Й�@g�j�'  ����5e��6r�A�V�6�dX�;;']��`���w�x�,���^n�
��x�s�X�'�p�qe^X  �$�Þ;{jp�gA/���=kG�1��5�1�w��%z7O]��`�+�:���|�O{Z<���B�.)�j�5�zn�-��;��n.�;�� �r�  �nKiD����[��Ax� 2�?i���^F󵜬��$`�ݶU���&ߟ�ө��ߤ#�x�=��o����'��q֤�a�6~)�|�e�)��?�+  x$��-��1ɁUNƵl|e����O�ׇ�R�ߺΕGp�c�?���/���Ċ���7��w�o  �È�.7��ᗪoΐ� ͸�� ����`vm���y���9�y���ڽ���u��h]�ͮ㹺�f�]�B7s�a,;��3�#	  �I>�47�ԅ�n2o�B�H��=`q���Ԑ�쮻���tK�
5ۤV=�A��l�5�r�L[� �e�>|�v7	  �����b	��MGrY �R�N9v4�^EgV�&��������P>  �S�zܔ]X��o��G�����@��~jKR�6�x�����䟡ds�s�D��i
��Q+m<+�  ��dS@ǲ���c�� �4�{��y��'͚Z�`m����~[�����V��h=_iW�=��*  �bl؞Ҙ����*� w�;h���<Ȁ�Vx�_b%_j����  <���
}_<�c���ۤ���ϑ���8�t�r����C?���9�G�v���N��F7����y�����HI� ���m������E$��ݞ�t�����N���>��
���>#9y�������l x���m��WJY{�O{/o  �xNm[eƳl�_]�?_ը[�o��׭��'�$V�����<��PC%�Q�G9:  �@0��������/����e�d�3��qGl��gZ��l��?����9���_�6H��Z�ji�@m듭�굕??�u��Uo�hx:F:�O&,��;ђ�}L�E��w࿿������aہ�v-��' �:���ό_���ԩ[�ݰڟ.~v�
����@{y�Z�(����ٛ�>]�^����=ۚ^��s�B>�\�k�����Bdiu8r�N�7�z75�Rۊqm���	v��_�w������)�`���w  �&���BØe���-�ߖA��<���$�<��X[S�� �����9�ϧ�JV��ϷPʌ3�	  �a�8�{^v�옼aH}�������S��&ӓ7w�u��|�:���Q���Zvk�[���O����r��4� Z~  �Ʒ����H���d�=��呜��͖X�fb���ن]�_[�a�}?}u��V��R�/��� �g1�]��m��b^�v���� ���֬"��Ii/z�  �gXf����/����H�2�sm�-Kv=�q�TG�ֺ� x
{�W��:uŚ��k�8�<�l.�Pxr�  ��h�e�0���A@�"Gpn���"5��7W(���#VX��'ߞ �-�]�9z���so�gXK{�������7  @a��o���"�ozK�W+����ug G�U|-���ڵ�⿜'{���  gA��Z�n�i?�������@���3���BQ���Ks_�<`��m�w9^*��:�-*F��7���s�݉�9�k����񛸃�y="ǎ>�8ŉO�t  �8�\-���rY�q����"���v�sq�Y� ���Q���ׇf�?���F�� ��B�����kہ���VZ�$l���Z��Uhi�oy��.�Ү���ɟP�%\�o\U�_��  ��ں�/���}���yaþ}3�+p�E�~{� �+G>~1~zC�a��K�y���Y��-��   va�g���M����1���AX��:��n��v�IĘ��)��n7e��V�O�ۑ3�z!w��r���tv/��]V��|�2[η���3M��*�U��Y������s�2��%O{
-'0�����o��+���Q��Y7(Xp�������2��Y~����3������n �����d�9�B��t¿��?85� ^�A-�� A{�:da�%�(ߡm�G=7ql�0����b�B&�'���n��j:��(��
��ד��i4���K2?����#ϑ�p��Ժ�Q+Uhr��S���=#��מ�YvN�����lS)����n�q;K�4n�H�E;.;��ȣ�'V')셼Tl  �$��E�fl�����Ʊ�7^�*C�q�k��`t%E�����e�t�B  �J���������{���_�c�3��As�����')��{	��Mk��F�Oem�n�3�W{�[Ԩ9$�֑�f볔�&�{��l��B�\Y���lCL��3v�����K����  p���"����4(Z/�Z{g*�!�ǈ��5�]��ũ���ů��,��Z}�x�Wi����"m(Y^���[i��/c�Q�����y��|�o9�K�E�Kc6�]q+G����u�l��\�� xoi=�؍��Ka��[�����I�q�mOcS u��>eZז�	�����S�R�P^�)E���N#  @	5�eS�aPې�ә)��c�dʗ���_��o��9uV_�7?-P���'9��M���wA��+�Z0��N�L�<�  ��Q�A����8b�?)cy��_X�ivpγ��Р6��\�����v�}!H�Z���w���޹V^��G����jWx��  0��;ZE�wm��6��1o�Ǆ�Ԣ��j+pX��p�
2�3  `,�wy�e��ys� ;)a�m��["c�k�����zA��޴��/r��n���z�P_�n�  Bn;��T�/�Ƭ�yV�?�s8�x�gς6{�_Գ[+p��/i�D�Ṗ�Y��_�   ��������m��lc��.=S�ܩ�Xv܍Y�  @�H3NK�.[����U;�[p&�Mg���A�tk��q/PF�C��Q�{G�(�1lo�'�,� �pASVΆ��:���L"b+p,z��z�� g�����zA7��utt+Hyܾ��h�������ow,ڛ
��[�6����S  oòoN;ܟ���M�z&�,"Z����9,��W;]z�Sv���g�(f�R];�W�",
4  8���4moci��O����vc������Ͽ��e�����,���';J�^�k3��.�YaK��@:��6�Q��-������~�E�=~3��Ámî ����/��D  E��zg����6�C:�2OI��q�zXszW�,л�T&�"=�l�qӉ�l��z[6͑:����k:ym�me���wӲђ��{��Zv�,���=_Y?�sz�ǵg}%�F�D���S^���w_�~��e�bJ��r�c>  �Y;#���_���F���ȸɦ �#e<�:;T����[_
  �'F��{k���?_�$�ˑ��O`�S���z�ku�k�p���Ե�e����cd.80iE���1$����=V5  ��EM�m1����� ƥM�2���WtDiӌН���-���O��=A.g�#%��]�޴�ă��k���+g�3�Um��y��cksb���K�I  �[��b>��\��Vx�*�8��F�  <������љtZ���   Fq�,�;u�A���h�4�(  <��O�P4�0E  /E�n!���v�Z(�i�\V8��  �Z��`�+0}�ػ]��6o���_�׽0D  @�=�3���a~�o�7��Z�x`���?fb߲�Bm;��k�<�1�;[��d�K����2�t,�#)�v���gY�^�����u�sr:�V����y+q��[r�mĞ�GZ��iF��  _�|_��;����^�S8��k�k�l	����[[{��J?�-�/�m߶�Ӭ�&-�o�.�ͧ&�^�r�����=�&O�{t�r���qw!f��  �N����Na�(W��Q�����^�RDr�tޗ�%����	Q�n�]�=c�L  8��?�f�B7`�w? ��i�q��N|��P��`�4����wF(x�L5�]���� �����jjȼ�'�t�g��O�9[A)Z�[�3-pC����:G�G:���y�����l>Z&/�`�,�ɴ�,�L�c`cX��/c����Kv�1� ^�l,̆��?�w0+����~!�e�s@��|�7�m"�,��֙��Y=!��㿿2�&���lV�r�&��׀���.�G_׮�Q��{���D+�e��m�����9�A��.ܒ�&�ڳ��$�_�|9��v>��c^yO���gn���`}PW�̒.�s(X=��  0����ÐO���4�Y<����rp�'w�������L|�5��g�ø��R��E2   N�w��N�����87gCp�J��|�S�2�(CoҟF�Ԡ�^�T|k�`��߫��t���|Oϸ�����R��͓���~��� ���31b?��=4�7�shpԎh;�����X��(@���������W�����E��F������<�v�тT�L�.Dp,�-]Mel�llW)�-��S����  ��[���Y�(d��[�+���?����g���[�~�d0�����8��  ���ae��L�h}o�	�L�NE�����9S捼��,��)�90s�S�3���X��X��  ?F�k\���ڲz���tޡb�����wrvl5��3���U�8<	=<�����W�	}��U6/�U���V�+�1?�  ���\�N�sp��؛��Z�H�k��)�|��|�D  x}�2a���>KA~Ǘɍ����n�?�&�|�q�)�G� y�#y��D�J��7��ݕ3���a,P   M���V�H>��e�y�
�V����z,����6�؎:�]a�*��W��F  �r��	~�oz<�cc���︵�/x��^r  �9�������iKЅ���J�B�༌�{J�D�ˑ��<mO�5�K�^g��s��~�>����������uOrti[���-K�ɝAM�J�N�� �����l����{{�  ����sW�*�6�7���Ime7���~w2��8��:��'���:Ǌ��U��z���� �%����F.-���pF����r�����X��Bt8��)w�]��51�� �P��Mwi��N�We����]���Bzc�9�|����ud��@�4��=���s�tZ�����s��Z��u��+�<�1��;d>ZW[�?{�'��`b���2�0w(�}�.  ���Qf-�>%�g9V�#}�5b���-܉�.�9)ņ?������34ɫFZe;[V���5t�AO���vN���^��f�o�-�{{������nZ�����~Y�����:-v��-�Y������l������  �Pc#^K�>�K�(n��Cu4����0u�}޳��̍z��ڞ� m�]  �({,�d~�	�L4���}Σ�,	����8�����t�ܽ��Y�#����z��x��2H�H>�+��-���}v�  ܂w8����yn����
�l�BA_�\g��3�*[6�2��;���)߶�C�v��d����h-H��n����� �WI�-f�
�� �1���b?A��c�  ���4O��\�������oB�S��.��}dU�o������wx	W-ܳ�h�[	�F[����  ���ʑ��F�]y9`��/�>���n���g��і���)�g��   x)�~��g>�u+p8���MW>���im�����Մ��l#  �c+�+̽�����3#�ֲq4+,���A,!��-3�����V+�s��_Z=�[g�i�\�U�ٸ�%�ϊ��jD]��I��|�  `3K���`�Kri;bda�y�ɶ"�w~���azn�������[ێ���ӫ�c��/��Y������Z��O�Z��}i�s~�  P�o�&�~��:���v�l�Ŧ �������g�lgmK�W���,��#g��&�0������r)8   G�;'�V���Fm���4M���^��ߘ����`�{��p�O��ތh�L���g9@x�As��s���g���F{����q6���Qۗ�A�S�ult�Ħ�k���4���}����oQ�U��$��������v��.�@�A�Ҫ�k�QU��%W��輤q�d~=�cUY�xѿ]3��\,W�=�B�p@�
�x���/��GIk���\^d��cL���񫓗?N�k_�xe��Ħ�jP�`��(�ɯ_��fpy�hdn�)މ�g�a��p��ns����k�n�n������rA($�k��~N�)
����6�:���8:@��~7bm&J?6;�T�ـ� s�츆���Wma¬
J
�B1���B�~<K`��AD
����i�_�`�Qyݕ"����h�d$.�S:߇w�ՙ�?>�3zF���ƏQ�h��P�|���R�܁�u��n�0ͥ�
�Bq5�2�!ߋ	���Oj��Q���Ƽ��0/��F���>j�6t�L����Be� �G��;�gn�xz7g,�p��}�:�Z�g�`�1���9���cZԇ58�x_G>E�����7��n�~SA��(
�⁈�X_\( ї��ۨK�%��A���ܹ���S��B���X�;�e}6c���F��B�P(F�ՑC�>Z��Y	���Y�(&�=�\��lH��2�:?���8���
��N����Y��d%i
�Bq'���]�#���f6Ѽg�
���G��!y&� g��ڡ�]��9��\&���o7�bt��=7�~QH�P(��s���}Cs�Q�Ύ;p܄�hA$�q��!�`��U(��c!����/B��Pl ��g�X���`��8��],����&�y��P���ub;������ڿ�:�@^G�yR(
����q	ܑZjغ�
''*��8p���Gc��{y�=��W;��F�|;E>l[��v�B�P(�7̞�y�8�E�{8V%�Ale�,	�uv}Fo��
�B� ���������^����₅,����>t�I�!�+B����+C��(���-')-�����1�l�gOߏ�ϻ�Y>o��s-�RW(
�1������:*�pt0Ҫ�wQtN�i:����W�<����x�f�y�(>����ର�nR۶�yB��G���[���:�[���[��E�w�V(
Ei3+���3<��Q�o��8�7Q�.��z~r��g^zG>���t
�Bq�I��[D�j��J3��Q ��fcV[�\��3$��yћ�`�.��4b�I�W�r���B)��ٺ߈�y�z]��+��^����~i|��sv\��ߡk�.�vu����~!��q��>
�Bq_�0w�FҬ�#-��<�h������7>F��P���qp�H�EM�*i��<�Se��sl��2V�_���'��$�����g���\.?��1����D�//�g�s\-�k�d
�B�x��E�_˷�f���49mڝq)��[(��#Tn���nC��́P&}Įnu�P(�V4��/�m���0籫l�swߨ��V<ɱ�yN� �\�mۊ�r�"���Ȝ�@4�)
�b7�H�G�6 �f|.'2�|8:m���a�T��欳����wE�q��m���q&n�D������3���
�B�L,a���b�-�Y��&lK��х�	Y7��
�Bqc�����������1?��]�
�ɨ	�N�H;��G۷��J��#�� �VG7
���NOiVJ�@w׷�G�h�H���ޅ���2Б�r T|g4����W�Ң=�P(�Fԧ�s~�a�Aڻ8^���z����@�{����P^�C�F�P(��p��	���P��W|�V�sE3�a���;�N�9m�>�<$��}��Ecz{��NZPz�P(�p��%;Rc�s��4S�xR�>�e�s\E/��]��|�#m[�\x������m�B�]<����wX!��ySQ�P(>Qh����^�b(V����{��?���0;W��PB�!�6�#
eǐM�K
�_�_�U��
�B��8��.
��г�MN�וɦ{O
�`�|6���rZ�Iʤw�֯���ؚ��yy�|�R�S�t�Oi���X^���enh�2�K����g�N�����̵��Z
�' �~���i�2���UnS�v��2L��E��cF!�
���5��n����)��?��p�v����En���E��	ߊV���R�ois����O��P�9��Ϥj
�Bqgt��ጒ�ic��E�r���|�0p���z~�;Ҝ�u��;�tGK[���G&h1���ʲ&�+
��Ibc��e�*���ۅؠ��pxw!q� ��!߽B�%�swWo��KIA�x?J��J
��s���M�ƙ�9�
=�&�`i�ߧ`	���]ށO�h
�Bъ������d�uި8W����\
�?�B����P�Oљ�FF�͛:��F�=���
���z��	��c���JsHڌ����ξh�3����O �Y�J����C��1kJG�	��L��?�gS�P(�(��
��|��zpF�m���+�����Kޙ��TP��G��1��PY����� ����c�9 ΄a�{��m�V(��c�����q4ͯ�&x��C(�Co��0b��7@���j
@�]��z�ڻ#p4>m���u�P(�^�hI"o�kk�	�MD��8�H}d�:R�#x?}#0bm��]wXk��NqF�x�G�"u�P(���%~����0��|���#.�a�GV�� ����9��&*��=�}���U(����ew���v����;>k���HO��=;�m(�t$
Ǖ�aJ�u���p�Q���9���~����Z�frf�M8X�,���}�
���(E��DZ�]�}m�<�a�����w��_��F���)�<�5V�<�lk����7j Q(�7�m&�����d�}YY�;���vC[.�n�ҹB>�0h�T(��n+�̾U�D�P|#�yY���6�;�����/���b&,�5�Qh���J�T8�菽aq[�KQFG�Z���A���
�Z�k;�J�,�BoT��|J�Z�yZT�w�B�Et�?��+�B�PȠ�j��fgv���O�F��8�'���R]��'���i�:��N�woG͡��[|�/|!�e�;;��̧"��caR(
�`C���8���F�H'�w��{�Vń�K#S���J�-�n�g��cE�������VG#p(�o���L�g��V���̾��GQqG�9�'W�!В(�ˮÁ�"�@��*'��Ԟ�+ϔe��y���������<R�
zoiWmN�����븠V��s�k�;���m�o�br�R��O��;#p�|�`���
�B�x#(��ek�x��Or�;#Z .ޑ�>g�˳A;��� 4OG��R���YS���v�{�H�<�������uT��_,��.��Q��q��V��$�d5d#Q��l)�-G�ydn�H���j5Z�`�6��礫�p�<cݏ��֨,�P(�D�7ЎeE������Lr2'n�h
�n:�n����e3�h��/"zk �%� ����^{��+
�b/���`�W�Sb�8�y+�oߕ#��?Z#ul�����=�w:��c���B�P|1ia"]���*��!�M2�;zYup�@�o	{#��ց~��Þ����sű�i�Kg��t��;�2�I���J�p���>s�B�P|>�1p�)�.tvo5z8|��S�L����w$�;pY��a�{B�)
�Bq2�2�p�t��f8t����
�B� ໯G9Or㷵�:���C�����������R��M�i���B�P��]��#]p�J߭x��B`K�	G����=�P�!r�
<��U(�
����*3+
.�?�}W0���܏w��[�O��P�#ދ�|�7����+
��f\gBi
����#T�I��x�%�\���K'�+wA��_�3���G�w������}#��g�n\�<�Gm��Z�Ώ�T �wj-t�W(�P�3�0?��1�ٱ�~]%b9�ğ7��u�j� �����p{�l5�g�I��JX�C'�)�#�O�I
��|�f;ZVG�2���T�y����9Kp�72<�_�����p�gx�ҝ�X�޼��u1?^�S��߲��߻R9V�O�~-/�7�Z���:D�j��m�ֱ��c8�έE.S'�B�8v�:�4 ��~�u��F'	)���,!�$�X���p�ڮ��j�N�A�����hHr!�~�8��Q���wAjG��ȴut�86;i��c���=��%a�j�#F����q����Q�ט-�B�P>$<_'L7Jό��)��K*
]�˗[a�wрw���+�{�;�lʌ�[`e�>ò� h����Ij%�h���v�ףA� 0��PB�P|&,�� ��ʏ�e�g��y⎶�'_9H_�`����U쉎�D����pEĨ]NR]��SΊ�0ZY�@O?�f���c�%g�Z��ڵQu\�^�X������|j�W�������<h-z
�ۥv�F8Z���M�J��P���׼2�1��+
�P8��ā�8���IZiG�< S����lͯ�Ƶ	&_��ā��#K�,	�D��u�r~��׆�ơ�Ѿ��93����������6�0��>�i�C�����|��y=���~;/���z�eޯW�\�i_���%���E��a]�u��8:jQV��E���|8&���X]f������!��@߻�+�;�\��eg��rY��ڮ#?�������z]���v���w�ʝ�Ds
�È�rٖ�{d.oB�a�B�P<�cs����')���̅�S��
�+����~���v�������Lc-NIZ��M	
�Bq �.�0�w����c�s��e��\T��|l�[���|�������Q�T�����M�����Q���H�g�dڷ�����y����΀c��X���\uӬB�xΣ?�������H���G��>߁�ԙ�+����3<�
��#ه����P(���q<�ê���T(�~�T�.�1F'ÿҕZ��v�:��{�J�/� �/>��(eT(�8y5a�,�	��n�	��vMN��U�*L�QF@�P(���[|�J��+�B�P<#�\��ό1
�B��P�ЯI-���s)�YE�����)�����G�o����N �Y	O���;Y�Cq9Tc�P(� �t|ֹ+�B��lS`����Dm�v�x1��9�"��pާ�S�&���S$V�P(F��6(~�N_F�Ckg���S~Nu�dl�,UX�*��>󙟻�?��͋B���5����{w���H�g�g;/q���U/�-F�K��"Bձ.��\w���}�}�:��^���n�XOyܮ�7��J�P(�A����&�� -����$ixі��s�V̩�f����v��S����ƭ�����$9��d%�<<C��/�:N��I��TVO�ji��ګ��O��9���Y�(sI �c� x�rK�K#�+
�졅1=5v\�Z��&�|�9��o0���g�4:G�7	�v�2��1����g�)�1���T(�+�Md))Fc�Յ��P�>��7�џ�0~\	9�M��;���E�ׅ|.P��B�P|6zh}�ܚt\��ŕ���N��3�nY�S0�Yg�8�i̞$�D�Fp��eܸm�Zm�Bqc�ǲ-���j��<�@gК�V���1_쨧P���Ϣ�	��u�Nbo̸(
�ǡqF�½h���P���ҧ�\�������U
�C�v��@#p�B�P|"�x���G)���墁�Z�G)����y�O�UV�#F#���T�D�8�1s
��;��8��A�d����wf����Ś;�KMJ�"�1H�@��V9�>Ix�$��e��[
��0D�3Q�y�8�LH㦻�O �����s�:�$��4\��a�P(��#F�3IWr6_�r��!�?�@�Ƈ����4w�I��){'%�]��p~��*+ǈ�����?�~|�|£ �/�(
���pKy���u�6\�����z�19��z1�1��� 6R�ڶ�ȶ�e7�\�͓��byR�P<1����\��a!�Y�Q�����*q�Y�w �+o�(ŋ����y��B��ӈ:m��H�8���3�Pi�F���O�A3l��;:y�����~�FMZH��Yxʜ�j�E�P(��K�����j}7?u%!�����ru�>ivp��Z
�A��vCh��߂���+t9�?/�;�V5G�-�՘-�Lߊ��o�y��ao9G�)u��y��G�6;�v�g<�%��Uy�Asx�\��x�L�P(r��ǌRB	n6���/��>ǃ�ح��9p����\���1�ȼd�[�h���@p6*M <���^��@�>������4MM�H�6��F<���P(O�گ�s��V1[�<5��_YC�'0+�*����1��Q��+z���|��B#�R�G�ՒO-�@JcH?�W))�P�u:Z�~�Nӂc���6��բp������U)~$_:8OJ�B6N�w��"/~��他{wFJk�5)� �2�;�[LZ���;�P(o��MA3}�a^LП%]��N����}Y�g�6!q���_�����%��]m#����� ��K.�ǻdB��$^�ݰ�>��l�|^���j<�;e�R��Z�;9np�k������Y���{��,Yv����.Σ��q[|y�oj��T���Ay�-2p�,�2ƣ�.��
��Z*��3>��ynp��`�ف���B��Lt�`6���g��5^�^�,��V�����܁���ہc�7Qr���<��Cc�;�(1}��P"�^UC�P(����_n�"N�o��=
�wi��w헫�ep�@�\K�+9=�Q'F�e-Q�h�w��B�P(�ֻU���H�Qr/�4�~tsM�fn ��OwC�~�'��{~ekNߥ���mq�)��N�1
-��[��Ȇ�6��Ѥ�'t���M3���a]p�0
�S�P(���W>Jd�s&x�b�7(W)��#T����R�½o��lY�*�g
�⹸��*�eZ��둈��y��w)2�f��4\���e��`�R�	���Y8#O>����w�V��$�Ř��K{X�P\�k$��}����8ƶC��B��p�b~}T���s��ȺÇʎ��W��N}}4�"�U��P(_��?�u��U�9B��� g��w�:�K��`��K�B����Ւ�ɦ#;�v�X�2�c�zwD��q�.���]���м=y��%��^�ͧeG�{<�H���s�T�]���U��\����,6�9s�Ŋ'u���kw�P(��0����CE��Eω�#��dͳq�؝�_��.�ӽ�ܽS�qt�}�������~���ծ=х���F���cSJeIrYK���8����f�`tCl��ƌ>O�.tB�P((j2��C�-[�uq��v���}� �x�_�8�C���Spщ��"h���w>��a�t�=��sg	�
�BQ_�")^��:�Rd�Y�FoOZ��#�D�#�Ԧ�kv�o�~U:Z����nB�T��J~�.�,)�x=r�5�댭]�F�~�#<�B��s�#$�c%e�V�w�;�U�֜'$�h��
)�g4�n�)�Gw�iZڷw������N��:0�R4��ox�R��6�:��w�1�,d�})�mDY)�k�KGS,:���E�������W��o�fPp�O�"XpNv9't^�8'��*05+Q1�LR�c�S(_��tƜѺ���"̓;Dq	��h���x��_�Mr��;���Pow�!������d���K�d�+#p�n�Ǐ��x���oM~����~*�W9J�x��|k�6��\J[�ɝ���T�1��v����ӗ��yG�-��V����A,C�{�;Q��Km��pY�~�iCx�߯��|]�g�^��=#��,�@��8�NN
ʾ�o��g�J�P��������@�.g!i����n�I˼H���2����'��n`��u�� X�����=j��KSS�P(΄���rH��jy%�F�u���`�x6i?�1��z#��_�UR�`>��[IY&��TFI1��R��3�>��N�`����t��iQ,��mԻ�[&GiK�m9��|Kmܫ���w��k���v�E��^�;���7��f�S(�����y#8q$��m��$��u؝X(Ļ��<��(���&0���K�Е<��&��ZF��%����LZx�=�8�!Kr^��8�%G���.Z�yCZ�Z�ze���f��/�V�����4TK�6 ]tN��fr��ѽ���F�3]'N��\���U,�|W�B���ץ��#_k��l�ܱ�9zd�<�)����iQ[��n9-=e����8��h����=X)�GD�0c����P(gcĺ���
�u�$�>ڒO��a�~��^�d��ߑ�se����h:�,��j��m.�ƶt�'�=c3�F���v�(�{��W9�O���Gxk7��Q�P|3 �Z�A��u1bMA�egO�qkZw�r'��H�Ҕ��3� ��q��kȿ/�q�SmK�G�+��-�߽e���<=��H0J�j��Y��·�7���c�?��bũ�|�����S(�"�7�C� �D W-Nq�P����g�e�v�x5�y�����D���< �&�v+c�P(�-;_RS+/�\�4`iE��C�+n�F�xީD���>S�Z>��v#�u��M�;����@��2��=%�c���cbt?O��Y��n�7�y��*��@�7|��g��T�8���|_ۮr��*Ǖ@y�*W�b]ۋ����J�
[�B��Uo��$�5�xz��F�𸝓.	����~�*
�?��:����S���,Ҭ�<ە�e��S{ސ���ʲT�����)/T�a�=��9�Ͷɺ��e�n\��y6H6-c��w�#l�|!��Y�
�jι�.0��A��P(� �O��C4��'��Щ/�����B�*�ĄN�$kb�4�Y�k� ����F1޳xχ��J��ˉB�P|��p����#p�5<Io����bH/�9�nw��3W��J�@Q)ݛA0.gZU�C#F�Je!��ӯ�T���x�R�Wt���7��杞�%�5�-���;�g!��1�QN
��+���*Pa�6����v��!��<5��W�D���/]̟rՙ:�@(�8�{�������y��[�ޮ��3��i}T�e��l��ͧ�B�P�m��Q�%��7*�}E_	��ϑN� Y!�Tk('�3kmK��M�n]�Aŗv�Ao;-�U��&`�$a1$vy����;�ɮI6��A�Ubi�\ ~�ԃ�}�����T���4��{5�G12g��%��r���`�eq|��#�[䫁ʻ[r��x��,,ɷ~���Ke�wY����N�W��[�=)]�8n��!ON�s���B�[�>R!?�4�F�x����/�B�P\���1y���'>䄪��RP�|���,�Mk�5����aH�;�{�4�i2���'�yDk~��ڎ�(0V!Ŀ���́������ �C��d7��Qv����7
�B�I�#m0@�,1�����,��`�(�O&א���k*�JRH�fTH	4ǝ#z���l���U�Dk�����څ��ӭ8|&W4�Ta�ϙ�ibY&K���M4��9yg ?O�|�<#�3����_���˄u²J�H�X��w��r���BgG�Z��	֦�X���_����+-W�[���+�XQ���
���W|_�+Z����H�%c���������Y��p@�i�����?�[���Is�(�1,�	<�P�e'sq���ӉLt"�����"��k�����}5�A�w��Ay��-[��f�1g
J���Q9�g�_R�^%�ƚK��ۭm{]�gBa��W��u*�i7��E'u�f9zk~M�n�u
}�ŲXn���
��S��g��!��Fè�1���J��ژ��\�:�Y8�`��Qyǯ�sX ��:*�x�n3�=�������n'P�:��ц+�%)�^d��"=�<����bb�s�=#?h�,��1^l1��l κ�V�q��&Cxq�)��f"Wx[�Ag�	y(�y������:�o����?���t��Ob���Dƈ��~F^�q^�[�8������!�w(_��$ߦ�+��5�yNך��v������3��˂��88��3s����e�I�(w��(ä1����!���SX/���w�J�'c�QS����kY瘢��tS|�����_� {�9���L�hJ2���������u��*�h[�3K)�m6!�b��P@)��7�[i�,c�G�i�l�I
��;���*�i�'�/��G�1
"���mKsGYK����V��۲�'�QGG�����G��~|�����L1��a6y�I%��"C='٤2���y9W';5(
���y��*.�:%#��D�ctzk�$�<�o�t[�Q5��Rg�z�=~K<+��/�B��z�O�����j~�u��Հj>4?���4`�&��Sj�.枧��J�jM���\��˙R�>[�')~s��@��w{�S��$'���u̜��h�q��#�`���Z���Q��n�)�eiG��Qz�
��0 �k�{���[1s`�Daq���A5��o��r��_*��m���-�4����)�+�_�2C/�Q� �d/I.��G���������ٸלOm�Z�ʮ^��}�?�f�(D�2��R��<P����ؘ\N/��?�s��-惼pi=�ƴ��(Ӭ|��k�rKWs �d�;�L�XK
 Ϋ�@Pxi�r�'/D%�Ȃ�ޕ���#v��b׳-�
�w��zv�js=����k�\q����l���F>}?��A�X8g��D��v���L��$�	�ES���K�ǖ	ُ��U(����������w�|x{�f{V:Ha�J)�H�f��#Un ]b��a�sA�v�����,�;[� Ji0�
\���g�9(-���]���԰���rD/|�pZ�
��8��k/g/=�OQ[��6��P(���o2�ō��c�r<�1�}[��M�㟣�C�ݫ�1F0�oE�)5<���.�߹���U�ܰJ<�����Q�!��Vd�q��I�_S�j�,�$?�{ٲ��ސ���ao�B��d���z�]7���N��\�2��R� L_b+�t�3�.����z������6�.os���K�P(>ܷ�_+{�c�Kw��Q\���2:^Q��ɨ�j�;�x�f_ʻ���T��͚�wע���N�-e9d
Ѿ����s-�����wh�>c��Th^`�o�ZPl��0A
�}E5���*
��U-:ߙ���i=m�"}�G��,�u��{�����\��D<�m#�Y"�ӧ{�xY$���;K�b]G�x�jX�A��>���c[ޑ++�'D��x���CEv_��%����胲�3T�ّD�2��8B����7(|.�y"�8��8�N��<[��9��!���2��u4f����U�CܸN_��:/Y�ip:8^$��Bwo����r���������ZA��3 ��N@��3G����x9oh1�����E������F����^�6�P(��B)�qA[r�g�yF������Xr�U .�����c�5���O�k�Ac��S W�ݘ:zk �b�kɯf���r!\��)#�fM����d<�o3��������s��^������+4�#��!��&�fB����T�d�Ƥ]�ȊE�#�|ٵk��*��|���43o�I���^K�!��Y;k�WIy"�H.^0��a9�|��`>|\�ڦp�}Yn,�϶���ټ>���y
�m����9i���D��� d��W]~X�����t����?������,���6�)&3�<p�<2Nq^X?��]���UY#p���P(>}JgB�MZiK�j�Lx���ZCw��)0�^Z�ڲ{�S�oZ��o�N��o����Ʋ�����c�F)Pߩ�Vv����9��L��X�P�a-#�����#�6̞��Gԝ�������U��Z).�Ȑ��E~�d/��P#.���w�N+޻�lF�'�x���JmMŲ����%D�C[�-�M�:�s����]8�1Qy��̖P�ۯ�ײa�8�m���B৯(G.t*�Q� ��������Z.l�%@EDT*�-(����o_͍���~����	�:��Pp}cp|����}5�h��WJ�T��ԏ,��Bz���Y�q�IC���)���R�%�8; ����?sZ�����E��O����pܶ1�]G��x�G������9?������#T�q�F�����X4�tա�e.�[��`�+�g�	S 	�"�BqWP�{����&Ը(�%��,*����Q�V�wKP�y�E��t>]t��T�K)�Dr�����`�v+Ȍz�3]$��Q�C�B�f�3���#Jm�d��i(8]�����N|u�/D�Ig�'j�y�4N^�H�l� �|%��/K�DG�L;��!Z��5~����΅�R��`|6*��6I�ZS��O^����螕O�����P�e����`��:�$�}d���`~2ޑbz7ֻ�ͳ2�嬻�{�+�.C
��n��:y���k"��5��?�����p?�`m�j@�{%F�#��ܕ$?$��M���^�G��{��-��1W����(L�<_0%�~�c�TF�"@C[yۤ��}Gxgt��|
�;P��af|N�.�����|�>[e�uyLv�b۬���&�.��F��Ɋ�;�d{i�e�s�"�q�.�_��&I�8�>?6����@H2f�g�ぇ�&��\>P&���3&:d�&~٫�����H��;�|�,��
M��YC{(oo�w����� �����!ӎ��в�]�,Ӌd��:R��iEk�~�5(����u�>e�\�i�� ��UZ3G3R��t�+�k�n�|��Հ��Vԉb��yoI+c�] \�|���c�	��L��x�vk=[�T�]����d��Z�t�Yr���agfsF�V �\�P(�����>���	p�qB��:-D!1	$�A�^֛�8������bzӪ؉��6��mR�lЄ�Mi
�.	ȫ4&w��D:���.�����(8�^r�)��0�V�z�9�_���7%��*G��J��>�52&\��9;4͹V�>-yp�+�I�I3΍)J
�z��c>%���T�L��d�	e�AYj��>o��ak �o(|W(���N������.�т���`��4y�FV�_�d����<Ŋ�e�
~M����O̧%CD-=�R@�~�VWQ��2
�Z+G�^�ե_����)�?�\�]�/�-�A�^�w�C-����7-����{��&-��(+�3<�x?�>e&�CH��{��%��_��4PyU�LNx˺ޒ�POb)���?T��n�9,�*�����:?��w�֭�zF�0��~VkH��]���am�	,O+��{tl>��x0'����5�|���g;��1���U�`�J�s��޻	�w�bh�X)X���q��{^�r�sW�k�}���H+#�.]�����.��G��#�U\���.P'�	r�Hg3��a"�+��L��)
�"w�x.f�b&״nc�ǵ�>�f|0Q��yM�w��JH��y� ;�K#��VT[N7�\f5�ij㳕�t���J���jU6g����L9S-ig]W� �.P�bL�8w��4��}݋w8н�a/�
ږ���w�I#%#
/���
pI�]<�j���&[
�Bq��&�j䉺*�`��{�~�|'�>�b�:M���g���0���SpĖ���C��kx�{pVQ�5T�4�U�QI��Rz��i�n��VU[7���o����z��x�s�8Zflm�2��m�[A�<�Fyc	�sn��Q7h��<UZ���^�ff�4��6�t��&"���H����*�1�ө>>$�;&N��@��m�����Q���aB@mΕ �M�;���1�׵6c��ѫK�"�����@z��=�l<��+��ٺcR�5�Ƶӝ������*X���> @�u8�
�p��"M�<h5D�0�"M>���\�2��b���2���!� ��8
��sq��M��{b	�2ɐ�^��~
�8B���Nb���֎�"*��-?�̸�xs���{�c5!��P&fJ7����)O	cxfl���=��Gj�J�$|���V�ٺ&2p��fZ���x������O��]5�/l��u\K��w�1Zdh�p��㡱��h��ZFT>L�e��m"�!?���e=�q�����)
�g`�J'���BZgM�}@��P|z�e/VV�M�z��g��*仁�\�*�L���g_!�Y�p?A��#L���W��߇�U���6g�I��$��ɦ+�ݘ�2g����C�g��Ѐ��}�ڵw�U� R��|��^����P/gݵ� �=:W�6��_+Rp4m6Ɍ���բM��g�]���y��z݇]��&�s�N�g���U�EE�6�2�E���<
�eV�|;��J�|���Y���Hǚ�yGcl8�9�k��$H�����>�Į������k�hB���~�X�-��������y��]�>k��5C2<����"���s��D.��y('�C'�Y��/���P1�QMࡢq:A�R(�a��G�^Ǹ��������
���*����L��Gא���=�������vkGwd���ݓ�;x7����:$������z,�8Y�� ���F�o���ź$Eo�mM5B�^���cwr�M��hi\6g]�?V�^��'B�W�l�cP�CR�-�����q�
���bzJR�~`W�7ѕEw]Pt�q$�V�����jOR�\)F�#\�-��=�����3:�����	W&��6'*�	��a�N��5yO�����B���*={�l�/[���yf��E��T�_���ʚ_;�5�zŴ�|�:��k	<8�Wz�z�+t��O>����	Ĵ��n���$��:Fy�/w?�,���'������OA��3�c�<��'��������њ��{٘wz�p�̅W.Q��w�R��~��x�,�vh�VdQ��b������8X\��DI4�N���/�x�@�|�x
��/�C�b.Xt�@�ˠ"�&�m	�@~4��N�H^l�da��?�"�7��|E~�e�1&Mu�Ü��F��˳kce˜ؓ�G�z&}�4fnZ�3�������^���N��uG�6pw�X�_G�m�.�Ŋ&�T�^P���u�Ӓ�x�z���ܮN�lw�jo�d��� �u����:-�k��c���G�	���B���^�����`�?���v��H��+pY��>�@0힢����H�&�܁@w`�k��LQ�
-����w�J�S(����}�:%JL�uz�XF.�p�D��a���������fr@Μb*�}�;@F!��ie#��ے�Z��g��i�K�B-�0�S��BR׭l��%�HH���4���\��ܳ3�D�����;��=8�oA�����u威�n�ۖ��j�Y�'(�3ş))J
�B�x#FЖsW��܅`^��꽘w���V�J��Ȉ�1�3�7�k�h�~|���+�q^FY��n` ze�]�0������s��i��8�<lZ��V%���-��e�h^��D�Sq?3��1p�y	g�fZ�d��j֍�7~4N�4tl� �$�gfP�-E�p�O܅C�a�JT?���4��0'#wV<{��¯����I��+��-�l��i��OI-���4%��}ۓ�l�tڧ8:��v��tylF�*�H����2Ȧ��=|:8bQ$�D` ��Y@o$��KRF��&p�=*P�s�p�N�0F	�B��d�[�Ʃw��@4]@ː&�)W��z��*�����+��2^+(P��BbI�L*���٩/f(��հ��Wٖ�v���K1��1�6٪v�G�}R;�6A����P�]kH�"�^u(|��5�5��{��[�ӝ��8KE?�<
��3q5WF5��q92\6@>��q�lF�S����^�z{�C2J�"wl�}}��X?�����?�s��8c��`Jr�) YKr��QNOu�u���B�K�n�B� �s�@�oX���G9o����r�$o�pQ! ���Nq ������Iey�F��Yږ<!ӭ%ǎ�Hs7�v�B�� 
�b/�B��� �n(W����<B����2�X�p���Ș�<w�������X���"'�pg��y�}]���pB��ќG�v�B�<����=նz���$D�����c!jKe��M�6W��6�}�X��!��î�T�m�t��yUU��k �nT|���]��AjO0���Ω+�j'Z�5����2�)�<�Uu(cK����<�k`S8�Bz�B���M[�nw������mt�0����� �R:�*���4����o��	|�� 7�K���Q(E��[wʸ�6m����(P���쏠G���rLT���㋳��%��
l ���z�tܤO�M�Rr��93 ���2Κ�0�B�G⛎n�.m�{��PP"P�ғ�M=�X�9��@�Z[x;�eK�l�����S� ��f�>e :n���WX��< ��wHw:p`1s�����(1+��ŋݵe ���ʿ(��Y�+�����rNvN7X���̂�o2�X���;|;� d[�o���\���> 
�Bq��}���X�)k�~?��3ˎz�_���a%G��7���&�Ɵ�G8�ӦS.]��V+��C����5��/�g�<O���oQf(5�;Ar��t��?kg�����1�;*�f��7(<���Y�&�mԨ�H<��PK�o��{��d<^2��g�J
�gc��ങ�&�5~
k:8���mD��|:��6c�Nԩ{��F#g��g�[s��_s���g�!�I]Ֆ^�<�{�so��;�d��d��@�1
j���V�����G�@���m7�a�k1z)��9<:΄���(�����ds�2ZtS�D��3���B��vad��,���ΌK�P7V�R`��"��ׯ.����G�9��۝N8�v��C?�׃.7Y�%�ʳ���t��'�j��9�z3�C^��O�>~}©�̛i�}s���>^fZ���]Ż8��(��I�؍M��>��D0Ȁ�2i��B��(��_@(,��]k����X&F�P(�D�
v�Œ�q�w9�A;��<ԹK�"�4N�k`��:�gg�^t�x�[�B��[ʋ�QNY(�J��ﾊԜ&F�����&��(Ն��8 ��D��?H�G���Ge�B�mhټTx���K1	��8\����YB�h.)ӹ���(��ס&���GCG�B��A�q/9x����'������(Ҧˤ#����r�����;$.���9���'�P�26S8j�<��KS���%∯�N�m�F�`�����߳mE'Hcp���}��
����ec(;�D��a��X�n;��5�V��;�vtԹB�v�if��	G�Q���h'�8��!����`��=�9�� �����}l�<���2n���}��E�yV�����+���EZ?p�92�,1���|�wh�#��~Lǳ��՟�O�}"��wU��r0Ι� ��cy?��c٬��޶HeQ.�@�Ji�q�<����l�b���sK�P(v��ksꌛ�;�.��Z�����7�c
�.�x��c���0���F��\̝>��և�n���$��"?��<
�BQ������"��3;��go���P|6��TK�s��T���2�O��B���ܭ}l$;��ͨ{eM�M����Qy� �a��	�3	�N�h����bx�QZ����!Fj|бd�3�v�iT������F��h�']��ӈc��d{h w���3'��,9�o6����ot�=C�#�~-h�z��^>�U��_��s�x��l���wL `��t�H��ͼb%I��������ޤ�ƞ���_U�*�{��F��i�z022��<16�+d[:���X$y���
�s3�}�fi'�U��I��{�x"F��tTIK~c<��<%\�+mDy([���e �4��C�3��K�P��^��^�&m� %(
���8�m��`/�����9<A�W��{4Bhʢ�%�~$��;��mQ�=|[��3���埆Z?�iGץ7�;���v���(F�S[(Ej��^9K:�e�<�okA�m#�m���ӵэBW� ��d��,�q7�7�w���j�i��k٘���1�z�pz���n�n���u�Z>�t[���(Ƴ�[-��\Ь�`��#�l#i��`i���K��+.�1:Y�m�c��YW�ӏ�<�?k�7g��u�ȠC��K��tsD�׾��9p�%"��<)��?�t��w�i��3���,�μ��P6��6�<�k���e
WõP���c��+�+
E�����T��<'&W��;&j1|[]6�`ICf�ӕ1���%�G���.֘1-�^��ŷ��f�"I�ԢX��S˛�'�'aT;�*��3R���U�A���-_ʷ��\���B���h�6�W,�?�$�2��)X�]���Z�􋺎0g��4��;�(
ŻQ׶����.j/=1d�o@���"�Tz����Vi����Y�׈i��h[�jA+�}wl��\�\^O�j�\U�j׈<�b�;Ճ��W���̇ލ}�m���tS�m̸�;��:�����Xjh!�E9dK������L��;Qã�X���TYe��챜�9��#0zr���nu���3rN�D�Ix�g-��]���nd�-�q-�������{9j}/�.��"�l���(�u`O"-�t-ezLۜڞ�,gX����y��'�����Q��X�����u�0�ﯟnH|��{�D����?��]��D`�w!��B�g�NՍ�+���s���Z�3�3�x>�'�ĝ781��K
E;r�ZN�ߣ��s��<!7�Z�Gb�D~(\���%uأ����H��XTvޕѿg���^�������{�-y�>�T�Ũv��X�\�u���){q���^G�9k/5!� mpƏ���Լ(:w9J��i7����:�ΈAi��ѥ���i>V>�
��6��S�)���o�B�P,�k���Q.��g�A}Ҳ����U�)ѝe�2��т�M��(���ˊ�k�F���|��3d�M��E�`<��z�Y*����Q�r��)o/~�:��Ϸͽ-�r�����	�c������4����}Q3G�&� �kg�|�M��<!�Bz�0�ċ����3�w2(��:9o�H_��������Ƭ���1�?|D�%����W�E�\>���>�����F�$��w#�zKK���̞�9�eA����#�������&�4�x�^c��s}�^q����j���#�]�!K3>�[,k��7WDz�n���`T_�g�#=��3D��9����#p+@Ü^W�pqi��`�k/B����gWt��(����S��X�E�M)�Ad
֘��?��x��܅��N�Gq&�?3���=�>�d� �Y[ӷˁ�v�sw���oZ|��n>M_iq`L\�m"�4/|�ױ@���ЮW(w����rA���MP[ʗ����i���B�P�q����f	���#֕����t�&;"��0Cɖh�bJ�Z�J
ŧbK�C�v��Q^f�*�Zo;�֬��ُ�P5۲H+Zv�])S�]T�dd*�)������'`m���"�^�S��-���5%�Q+�!�bg���x��I��xH�@9�K(��Q?�G@Y��c4��P2��Ύ
������6؎���V����S?� K�Ց?=�����acA'���w�:�X�[J�$�BY�u9��&�V���O^�e^���wE�(X7K��*)}�He��B�1���^����> ��@+S�@����2�Oyɩ�k�IHu��������c�h���?��ǅ#��K���+"��5>4�}`�'��l�i)>�G��b$���>\��`};��N܄B�P(.��_��@:`�2��!Is,?��dMk�1.7��>�;J�
��Z�]�{e�5�u/9Y�DƖQ��������Z�.����^���o�yCq"�L�^�Q;�ߎh@\�Bg�O��<�5
�6���<���	 7�B�Ȼ��NC~�����)�eV��3�LɳG�����66��GF�2.K�?��lb̎}�ߞ����̺ �7�y�$k�ʏs4K��o��7 ����zTE����sX���3��]���ql+KK�;L�*�G�z�ˁ��A~zݏ��tC��C��ް�_�i#*d	��&�����T�2����Fj�*;����^�����؅uh����
���K**1aM>��)�w&�>]��5���J2�� �@ێ��B�/�*�@��R�7b��7"�R��S;�Bq5Z��ۨ�%�!l{9�����Y*��׬��{�v�箍Ƒ�My��޶)?�x�2�F�S{�u��cP�K������8n4b;�˶���a*FPg<M11�oK�k�q�xue�<��>��+Gޣ�YtF�mM۳�cMp��2��"i��Z�h����C�Ξ�y6�{g,�+���������_�n�ޱ��V��q:t��'Hsf�!�P�*���>[���bX��Τ�[�ˇxj4�ӻv̶����,ZO\�o0N0`!ʂ(L�,'쥶���yr҉/`�׵^�c��oBɏww~l}��*������rܗם)w���k|t��V�u��AVX�o,˟�h]y�9MX��n�N�ڹ���@�zx�G귕ר|��Q����gc��#I>ǜ�gvg�Z�שS|����$��)5�{jE�������~G�둝sB�(���K?��ʒ�w
	2W����;�����P(�A�:�$/�۪͞���E#�~�?�E�� D7� $�9>�?$?KV{�X�R� ���=�`ġ;�%�p����l9�|
�uw\��O��[���zz��=i�;Y ��D!RB��4�q6ϩ�pK��#�r�euY�9�����^'=K�Q�S�f�����Ir�j� ��.C��%J�9�4\9	[�-G����>k{Z]Ik0A�
a������E�B�n`�K���c��cT͇� ���D��b��q������+��4�r[�y�*a�]$�T�BZMT!�����ӰtG=Z�\�\�7�(̕�[�$zS��?,׵1z��P�\u)-6���$��:P���
�5���]��8�5��V|�E�(QY�[�7�
gAf&��(E�!F�:��3���e)���%�֫Ƥ�@��K�x����|Z�x"F��u<8�3�ԎV�e�u�M�z;�OkN~X�.���&�L������\�1���$�U��L��y�D�Heb}��5�Q(���]���-�;�%��%;����PtTv�hDuU��Q�T�Tb����&��^�9�����?*m$��Զ��<����ϻ!�k{yڽ8�7�p1-��HY�nso�;�[�.^+Ea(峀Σ�c:˔F"��͆T֙P� > �=E�[���f
Ǳx�Cbc2�ǝ@��?����uy�r�5tC�ZV�z����N%=��w��3Һ3�&�i�i��X͓Л�P�E>r�-{������P]�'�3C�B0��kpU�r�X��Iӛ�����6�|Ӣ��v�2C�6�BV�������.��ԴR��t�|:��W�0�+�����=�4K����/	Y��ǩ�>�Z&��$>��o\󶱔�c��9u�5&�#�"O��#���"�Ls�uq]�0\{x�#��\�9ź8>����KP��Q޷�^P�^��$1�v�+������}��fPZsm@��1��9Q �R1�4��nJ���$H�J���m�Ӓ�1�=�qVF`kA���O�lm0�Q]�0��v�ح(e+
�G⨶%ѷ<JѾ�L��b�q#���܃p.\�K����V��L^>�g�-cOsf�ʋ�������c�Z֐�z_9������32�Q&���,��ltL�kY;ZD���O_�ԗh�,}��(:�1E�-�Nh���I�y�D��f_lJC�ydK�+9�]�_6���g��RS�ef���밑7d�vZ��ߴu���'3��zS(397�gªgG�"��2�&w�1�ˣcutPK��Lޭ�;�EF�K�զm<{�*�^K��,y8?=lS{���;�:�Q8"�M�㞮�Ɉ��-c��)��V��<���@ע=LO����n�PM]Q�bAцJo;�&Aw��C
�B�Yh�>D����ad�۝�
��}�����sE�+��μ���K�<��s���g�}�|7����H'�IH� ����lp`fB��a���]�w� �P(w���iG2�-�1bT�
qkp4�ۨ��y[Lٟ�S�6X]��V�O
z6�6�S�X畞�8[}����.%��f���BX_���N��z��q���R�e���*�Ii�Y{���}A��+>T���_J�~?��eI2����sC�C���+U`�F7�n;�#������3p�E��U�����?�[s�B�F��=�HįB����b��\,oC$��zDѐg=��tO����Vn��ګ���{9�CVս'j�%�%^�� H��q�`�\��º��I��ICKo�Q�P(���+�}(ߖ��s�uǧ,��}�lL��Ӵ�L�{Ԯ��Gڸ���w��@w�K���V|/��}�'��a������d1l<��q�}4����|�z�L�z_��qie��.lU�Q(�èo��ò&E����<70��!��Nv>��-N�a�������գ�`K<�Mj�5�y�#�L�K�b~�S�9r6#o����������[�=1�[ p��I��v7��j6�{t�
>g[.7m=,�j��[,m����H�~�WM?��-��nҵФz�U��z_uG� d����e�.�5�%�~[�Os�����6R�M��jJ�}�f����ZHZ#��G�:���А�鐗��h��;@�����e��.����N*~�J�K�c��lL�K���~�w�����8�!h"y�r59vX�6���g�C�P(�c-s@��U"�i;Zp&����/ ��1��0�5�����ˋ��	��5�nn�X8gyl��������gO���ŵ29�P��єA�ZS�f<��/���CO[�Οy�X+�b��H�ٻ��E��Eg�����+\�M��к8c�����`�3��������[���x��u����V���8
�Bqy��
�mܐ���.�@�BI��u[?>%�2���
k�u^i�M���.��<��5�t!�
�R1���Z�H�$�%D�:ٳt�����g��?��%G!�g��Ҷ:޳$T&v�Z�� >w��5�Y��^`N#�&;w��8��q�����Y�-H���������#o��.�r��'t
�t�6D�)�RF��u��2[}D��B��_��5��H`�%��R�֩r�|���fi~K�6m�k�OVG0�<ͯ�������q�anM��� �: �-vo>.�ׁîf���\�}a#1��8Qb\����C�O�Ok��� ��5��Zc��F��^����a�ؕ?�Eng��3�mWC��J�P(U�΅�2u��*�yE���{y3J���>N|�&�.�$�4c�Y!�Ti	� �W6�:�	#p3[걻��\���ikI��'/�wc�O/���Y4�%!��g)bB�AC���q��ǣ(
�`	��ܡ͜���L�]"��Q[�W�)w�&�����V�d���]Q/h�h,�ue�D�$��mFO0�]H�������|阳�c���t�9��X�b����ϑ�F���g�_ھ���@��һٜ�규O�}ٌt�n��ğq���Qr��j���gZ��B��w`ㅰE���
>�Ӭ;��p��坓fsd3�I��@��gG
���aԼ�a�22E���ň^��nV��\�T(
� q��d��4�nd�R��Isz�
�T������.�k������rA\�,`�L"�@�r=*�(
Ź��h�䪮+V���*��9��3�X��:��Ы�NBY%TM��,�#EX([��#]l��0"��[ �sO]N��]2;0�w:���!?Gu�5ǅ�v���ny_�e�z�d�u7�6Rg�Z��9Q���>C85c�v�{�d��w"<��mJ[%��O#Ӓ��ʒ��t����lv����<8ׂ���05{ �3Ԑ��E6�x)<�/`xI����-
AA�g��*�c�CG���B�P�xgD#���a�M�#Ko(q3r������l�cJ3>%y�p�=�y]�4��N���q˱Βe����S���P�xL#�2/����l������\��2�3��!�;"���&A��TWs999�ԉJ��q(X�f='���,�2���E�ѱ��Mj�̭loqĨ���/V�b��h9ƣ���e��gO^�7H�����no��H�F�vR˷p]z�Pv(�����#��s_��Ι6[Ew �ݵe����b=�;��8p���gV���O���-��d���S�Bx�_t��̠ȭ��'D|����/�*����� ��Ik�t���'�eiC���_-Y�����Xf4sC�)��(�l逗R�F	R�>U�)
E?F��@@�������>�ۋ`�3�K�w��z� �"�˭�I.�l�]ʟ�^����PH(�Z�P6W�n�M��S&&7��O?�_��DtN�Qy$W�Ղ�J��<�oǝ��
�B���2O�w-��4�v�R�]NV
����|~�ZoM,g^�L���A|��66n������Y1��I��2�4���x���z)��^��?��G�A#oм%=%7:��Tw^?)��fOy��i9>�%����h�l�ⰱ������dU�ރV��>�]$3E�>���1�䁱�ׁ�@_���˿�'D��2N��$܄�ҟ�-�9�pZe������R��ᷓ�hj�5�؉�;���<;2EhXH��BTӂc-��NtDo��9�ȕ9�[!��G�u�g!���
ŷ!� �Z���~ZQ`��^���P7��PҐ~�J���LeB|F�,1��� Lfa/��td}���ؕ�`������l/ӡN
�B�1"�f��3��ĻK�]�f�Ӈ��գ��Cu�D� LOi��\�պ�:(sK�c�{��'�:�m�P(�]�Q��Z&�n���D�r��G�w���1 $��|�3�@�1M�g���D@��٠�uٻK�}e�2I!�gN�
�������q���{Sz酗o���S ��A~d��0�hlHgqn��`1��:@���h�%���歞�a��#��,��hw+��ԩ�QDjMӪ_����&�+�5/��̽��SVo�W=K!F���hX�ۙ8�k����r���g�[��T���sڌjq����G����3�X��i�vx��`~�7��(�Y�Ǡ��׈Ċ�]��J9BS�s+�S�P���"���7xGO�f��j�x��5o�kn2)�wȫIhIe���BY�w�B��\iɅ)+�k�jB�&,�D�$�+i3���S��Ƚ�X��~u�l����˸sB��
�Bq4˓B"�k����x8�s�\3�����J?��?�B �wIi
ŧ�S6�����i�g�ES{�z��L�E>!#I�l9D�#9���Gn���G�Q(�O@��'/�1��;�R�]���0�� 7���s�.�#I�&J Wr{�I�sшY0Ȣ�F�[���7����w��+�=��#y���3�BFc�G,o@i���<p[i�;��γ7�x�͇'6��Ts�Dn ���S8�эQ�EL���ɓ*�eIZ��o^�<HS��HZ�V�٬j6�q�|1�=�h����T~)��k�|�
}�x���5��i���5��1gz��ڋH��\��^1@
�B�e�~zw
����"
�!r�����K9y��s�&h���IX�Iǜ%�}�[���f��!ֱ�čÊ�:�mš���������R�ո�_D�,��;��<�cr�B��╋+��ƫ������I[�_��M��Ú�Z��)
E+j�Z���l�@�RZ�5F ���������'��ZƧ%r�B��,|�.�G1�O �%XX�@�֒>	��>��Q%�`JΛ���Ʌ���3q��a�o'D:�6�S\|�W�\��`1?����< ��F�+2q��n����F��B�x�;��Y*]����UV�Wx��s�R���35BŤ�����s���9�"y�3\��dfQ�P(z�^���(Ȃg7'O�l?�%�8f��(g�5����:�P��*���Ar^
��L\�H���.�Ǟ5��~����l��T j�\�$���=%�%<_Al��c��������2j��>���P���XY�m�+��;'��g�X]�r�ef�����p<hD]�#�bu�P(>�H5��Q��Un��Q�W�q����U٬t�%���Á#z�$-�P�8oR�QCY<"�EW�dF�0���z}��,����z�
G���9� dCs�ifS^B-S_�9�����+e!������?���� l��籀��
HE�&�����*�p#}�
/��1y�[,pJ�-�	��#�Tn2��AT� �E�V�E�y����J{�Sșg*
�8�S��Th��J�fb�������.2�YlT��ٺ��ԅm�;������ڿ�d_��?�AFY"�)�(��k@!ޑ��UQ�d���8M?Ͼ�l\h�(G.u��N�ʚ�䤖F��LF�8W��}�΂�;a�����sؐ�����bV��jS�(��˭�`���8��ª����V�
���ۍ:CtO>]4�Y�����=��!�:�Ѻ5V=�5:�
�;Q7�':��.Ք�q�A�u(Z� F�Q�@�R^n��I5��`~��U<$��(o!�L�O��F��Ou�P(��㔮�/��Ֆ��ױEV�����y�7_���� �&�x�!H)��1zpx}���^��nP�8B��y�	�ɚ�i���^�O��~�5��3��C�銨��+4Q�I\H����s�M��Y��f	|־�fb�b�1Ă��)��H���-��1x�~�vW��w�:���bҎ4�.	%�;3s�@�_N�� �-�S�������`��/TcO���#"p�ЧP(>��G��S��po���'�"|iQ�ew����
}>Š)t�>��a��
B�@��y�XQ\�=_��S��h�O��⓪��y��)2�g��BqΛ`�`B�E��-o��aMS�)�[d�V�w��1�Xe����)��j���V�H�m�=�*�<:n
œ���bB�9�A�7�+Úe6����v6���[�d�G�i%�T_����B��k���(���e��l���O��	�y�j�QG��pB����8p<6,z�ؠ�tǧ,N����{B�<��c^,��a���*u�I�7�p͂~�M�9���l�;�^܅!(�yY=���a]j�����������^����1�����,
p�1�����" �����A�3=ܸ��qhtA�P(灟�yLIF�� ��(o�WδD����e^����$Mt��gV3��I�� ]tG�Du��ڎN�g���;�����h�0�O��C{䩖����i��B����ـ�ՂwVᩞ�y+�ϗ��6��6�^G������ޙ�Վ��L���:쥩��X�P(��u�H�s׺�i\M�Q�,�h��;-��ۍ�/�(�Tʇ^W�P(��Yٙ�9ØQ�[^.��ɒ4� �(�w���{{�=�99�'یW^)�x������oN�QXf[��$2�����Q#�����:�7�L�����k+�Sa�]ˎ�zI/��Y�����+��|��c,���p$/���y*P6��ōr8����Vj��_z�x{K9��"E��.��H�q'�κS]��N��@!�}�y*�.Oٓ6�j�s�N�Ä�ꘗ�>}����ɬzZ7��+�v�mғ�~v�$��khK��e�����R�FU�*�� �;G�O�����#S0�S:>%�5=��Rgm'`B�'H~Mm#E/������?�	e�`Ĵ���y�I��kvޗ#��ݖ�}�H�1GO{f�s�n¼�>m�3m����F��!�|�JMz:Ji���Q�ș�����{F�y�GdЖ��#�m)��$0�:frEI�`6�lT���hhWr� k$\:
����mѲ�~�6$I�	a�_뫋.���z'��E-���(�A�P(�*��X�Q�񳡈H�H�T�M'�f�Y�4������>�T�F;:+9��,�@�SqW|7���#�p���r@�A�P�o�"YP��U�����M��B$g*��-���8�8i�4 m��5��(T;%'�(1_|2����6(��M'�V]�`�o#��
�pW7��7jJ]Xb��X��wJ��9���J�s�����٬��Bƶ1u�)�x�bz�PC��PUك)Y��Jqw���@�R�a��j]��|����3q�G=�B��bϘ=u�s����1șM�w|sBn��q��0�@���g�Z�W��0��}̖�pI��q�Cq,}�|_�����H~_�
yg��}��\�R[�tF��</�'�0�V������4�$���_��x�>#y�]L�B��Һ�m�h(�y����K���w�S-Mb4*t��~~���ׅ�_x���S��(���և�X�i3�����i����A;�9��i�L&�'E��_4��Di' '�D9]�����S��A�`27v1yu�G�߽e��tO�=ys)��ԃ��D.+�ʠ{ڍz�����9�E0=I~{UX���'LC$f�5{D�^�q�e@�>���3��C��DgV���/�h�̷#�{6���`� [:h���:��V���~/$��h�
�Bq7�cu�W�� ��@�-�>,jy�͒o6��=?�i[��Xvm� Y��̩��7*�_�s?�V}*������~U�p�\)��\G5(W��!���<� /�peI&�!Q����'ׯ���X��C� �cB>H�*����7�c��婙9�5w�q-m�h���	h$���$o̗ϟi2���^�n�ڲ[�K��	5agv�FX�)����'*"�<��&�X̃��z�<����hx�f���L2����|�3�\"���Q�L�a-�//�j����4ǟ!��]|~Xk|}\����1���;�o�xs��9*��ӏ�����ڤ`�j�LӇr���0��n�r�������:�2����3E����ٚ�c��NN��uC~��Y��'�N�lϴ�Ư�~���h��vA|��yCV� iHm\�%�ɏ��V�@	������]a��H�?�5ܚ���g�J�����X܍�$��U}���7�(aZ���5'R�%�r�[�a����ƭ��i���|#�P(��ٯ��]r)+��VƔ��Oe��I�'�"�Δe���E����E�)ZK�rX�٠S�̏����z�o����B�ba�[K�N2S�(KI����W��_�����3=�4����6���2V�`\�md�U֔CTX��HY`Ʉԡ�2���Yi�׶Y�8�rC2�8F\��|��.�'l��9o޳`��e��}��>L���� o����îб�w��? �6��.<?T8�Wrx�r����$T�u�ɺf�n.�_�����%�tk̙B�Z�r�Kr�%�6tF��¿w(3J���Sz�t�e߂�,y�W/��MNN����Q����Y�ir�>�\dY��ZB��h����h��|�&C��9�B��m
��8��>��e��D�]��lcb���m�Lk>1��5��e��ȟ��!��N����V3_^���}��5h?*�@��<�g~/�*����[Y�	eS��g�g�
!EN��z?�/��N&�k2+�p �mj�M�}G�Fu���=�ْhh έH�-Ӭ۱f��� i��$1\��?VEԼ�[���T4H�Pi��v���4׭0�f4^��?IЧ����Ģ	�Z�A�a��K}�
�R��c��յ���U���&�e݅��Ҝ���ۇ}9Ju;^BI�_k}K�
��uv,lv�;��P`�Str�
��W�]ɀ`+Dw]_��H;��1��+���I;�M�&Fԫ�?��9����#��mHk"}���.xmK���q�.FS�P(��h�>�
��3�z�96�qȁ�dS�u�r=<�c{=pF�9DD#��X��F4n���X��_�i����Fr�����hP�6�3B��G��a����{�1 <R/�|TE� _^���>#)����v���K�Ec�4
�(����*�&�S.E\���b�6����7��Ҩ^��B�N��	��{f�,�af����ZZbB��Y֥i%ѵ�f���F���&�����%Ǐ82D�#�8&��Y����3������߄p��GEЇ���M�P(�:S����Zx���g�^?��^������}�	c}�b�vu�L����X�Q���D�[�վ��6�H�8/�i�|��:Rޥ���kJ��-�i� /�ygt\6�fAf�O5�}F�7�1$�<�C	�� d($�A=&�f��3B�d 8�Pg�4�6	��ù�° �ǤV��A�^�ϼD��w��|$�L�S������K��[*����v�[6:yX�o�����|
7l�gv͖dM_m��<�;Yڟ����e�tjqp�}4�K�����}}���;����ShV���)�޲�6PEgȼ߽������N�ԗ֬_M���#0_�>Y����J���%�3^%���E_h2pL���ǟ��G���C�� kR�з.p���t��%W"��*M
�'�e͔�ҵ����_�19�K�Kd����G�z�����D+ '�z�f�߰��f2�+�3�����zl*���F2���耟gğ�k0L�\G���Sq>�M�X9��5�.<��wFf�O^2N��4��t���s����s-��yi�-�����vE]�5+���s�Z�m�_�V�fy��Ne^�S���	uΈ5�E�%�_2�dqm�u9�|�i�,���V/y�.�se���DN�����$Ka�&��\5�����_/�.ĩ��ڿ'��~�ב�TQ(��(�2{���u����B������@�l���`96r	�����7�m'<ɾ�����DZV��\7K���RZ�(Ϟ*�
���Թ�����7�-a������s�L��O�]����.ϣ��yR��Q')�,��$�Az.�-/m�y\����TK9�氵8���H�(���}��c��!X^���3�u�h��q\IP��0�^�,����c^P������N�ܣӒl!N,Z����eA�J�� F�j�tu���v�I2-�?�ܚյ�*Wx��������>�T¹���#����H����6�S�ѧ�� �U�n�m2am��fd�.g�y}��#��;.;�%͟Z_�����H����,���NB*�O͏���@a-4&�s�G��S'��0�c�[�78^� �)������?�1����D�Ւ<juX)��~.z_�{M(9*��P(�[%\��Ik9_5L��$����!�ǖ�����q{�/�3hAA�����lYA���+Ű�S>� 7���>�@����/�o�z��e<I���2�KY+�j�.o�No�)�̶UG�YJ3e�e/�ijy�x�Z!��m���X��3����{��Ǌy�>��s��\�v��i�B����U�	v��_䰤���~���� ��I&Ls��#�/�MaF��~"�3�/̍�MĠC���7������"Z�7��T�]%��%X|[�����TQ(�^䫵Dg$t�FBJ�6(Ӄ�eՐ����T)R���/F�I
�3qVdN�5��E`F7�,y���SQ�_�����8mm�M}��7��JQ�:�H�ﵬ����:�)��mڼ��DU�oh=���}�o���s �f5����J��rL��g�������W�<Su�s'�'������K_r:�(��\��<�CX�F���kpG�@�c��@��p+:�tG����9	��.����Iy�1x�L���FaZ��������6�����?��ϟ?��<����d��暃
ȱ#vŨ��-T����{�Xے�<lU�sν���� ��lˎǂBk�,C�G��@J�N��A����! ����� ���2,Î��r$��$J���%��D5�&��f7{xӽ�]�]k�U�k�Ͻ��~��E����S��Uk}kժU%�z��#(qc#]i�L����p*�;�J����t��k�-�~����PU�V���e:e�h�2���zn${�N�t��t9.�I9�ư<,�<VM�2��Ft]2��v������rj`���;��t��eu��;�:dT���{c����]#�+�d��Ea��5R2=�(Z�֍v຋�6�eē��:��=�]�"D��V�I�8:1���Us�FSN�X�"�s�ux�v��V0����p�a��]���r6`gi��B7:�A�S>�Q S�.��Ø�xN��y��w�</t� Ʊ#�[�|��D��u0vl[�tΛ�q=��:]��3���xOKv����m�.��r�n�Ձ���:�ߤ|v�P'��0��	���h�@ݤd�~�[���{��=�@
]:��HN',�0A6�:���8��ɦ���*�,����b�3^$ف��;�*����>��%�~k�a[��t ���/�����)ٞ����!�չn�UK�rJ��vP�S����� x&���P���~�Ԋ�W;�ȸ�y��Gưܸ�A=�)T����\0]��nP�k��Y�1��^0<���?ؒ3����?r�N�Y�ҸO���5�u��|`�Ʃ��dp��f�B�I?(��I�3*vB6���6�T��m���~k�H���qwq�L~)
S$��行D/N��мW��"m �Ә��4�X�qi\�(v��:�C��X�s��lI���׺�u�N��qN�F7�=��������
ɳT&5��g�C
)J#��d�,�T�`�_8q�3��A��J����Uj= ����9N��D����y��x�r�� �����x�����5T#K-���Φ��##�z����)ۢ�-�e�R(�K�jZ/�)�WX��v�y���2	Ι�(�q%�8v����˘".�J�Ͽ��{9ve�$�F��� ��T�g��<���t>j;E��ݾ@QJ��?�Sgi��c�Z��aښ�)=��1�n�oY�����dJ�'��8O���iO�"m$}'9����y3`�AǺ>�p�o��V�kzi���_+�Q��������H9p�Mxa,���A`��D�L����E��!�>-`t�Au[�w�Y7��������r�����# qhd��܃JS�6el�Hc3Q�/ey����ZhX!.�ey��6_�p�ADvǧȜꏛ�3M9��峒��Y�0~���S���2E�@�ɂ��Yw&�nt8�������˭����[whG3.h��ft�V�5V����M}Ǧ)Az�I ��1����W�Q��m�w��Сs&� �c�϶�JRr%{V�|��h��U���@rI��M�����y��zm�N��:=�4�t1�w�-�J��\T�LVodH�.�����`����;t5ت�͠��A"pY|����$o{=d�x���u�)�7�x�y��܃L��2��vCq#˭����c8���6�,i�|�.W�m�Kq�|��.�H�cs9�X]F�����C�w;_[/�wZ�����ud[G����u�[[���$�*���HAs&50Ϗ���wrЊ�TY�yi{�/XMmHv.;�W㓜�ְ���@?�3����~���f�W4k�i��Se�de�(c4/�=�/��x)��F��D7o��N��:]�G=��1��v���.���2�x�,�&�AUmĎ&���5*��7�lt���Н��=�����og��+e}�[%xdB'��1Fr]��b���X^��w��G����i�C2�Qqv8��غ����ҧi�=�#���?.����>���Yw�ԍz���k>���.m(�\Sc���cH�R�ߓ6�=��☶Ρ4c̀<���ڼ} �L��w�z��o;U�u���nU�J��������9�vj�2��8�����#��|�D�l�����}�Z *au��2Ϭ�^*|�Z���u/�o�5]y�9�g.��v��ز��)�Cp)��D����8� ��>��O?_��?݀���޳(��"P�St:�����pb^�1U]�'c!"If���}+�̦q���t��.n\�.����_A�z��.���qO�O	��Ъ3�o5a�}{Lz�pr����z����d�n9f�w��8�	�qߦ��%{����2��ųsvy,�ڢ�3/��D�*@[��X`�S����,I9���);��\�$ذ�Y�36JFC4���l^zॻxo4L��ù�S
J�s�-o.W���tY;�vm�N��:=�4��_fc̞�|!��✂�����Be�x4?m���#����ܳ�-��t�sV����tB5[�7Q�m��ETY�,���L�U��yP���2lƭc����,�/��<�JM+ J��b��`*��l�r.����(cz���h<��E��ԗ�p�v�l�� Sˑv.o�{�kֵX�������~�2b؍�VE������x�M����$3Md2:�'(�m<F��rk.��|5�X�iBn�'9�rk�c����p�����C�H���%��Q�5_���m��t��t��k����)�>'��u�NW��:�sU��v�/SΡl�}w?(7��������ͷ{��
qL�f��k0�k{Pi�_��Юߕ�5�`��]�*��5��P�xi��d�J��-���6���	N�}��)@��g��W�Bl��~�'��4�w�ޥ=�Y='W�F��[[k�=-'�q��'��s6��Xεgi�:�<��si#A���t��=P�˵ޝ��+������Q3A��P��<�u��xyL]�>Ny�d��l�ѩ��Vgu'�,�f���y��z���b����l?�əi��_�L�t+8�A����i�����m��Y�r�����q<!gP%�<d$�Ds��<��;�f�?����OO�u=H�85�P1�=�
�i�"J�%�lDصTT�O��� ���h��R�gR[Ύ뺊�?\�3}����
P-M�8]L����b-)���J��A �"-+'���|pd�_8-�8}�~w<޺!R	���d$Beb�U��\^tcOum����%��\��ދ�G��F�X)!�p���ַT������4�/rB�#�,�v�Je �w�y��s��O(��*;y?k�'YJ��S�\����,��߻*#ek�\@/��)���:]�V�#c���os�a��*��6�I�ji0*��4b#F�Ý6S�}ê.��1q��5��	h9ٜ�˟�c�;w!<�����9BY��xMN�%���9#����b�e��gZ��ٟEx�ߣ�e�v����!`���b�q�#�i��S���F-�3��DK��9���s�Č��5Pey�Jv�㕕�NK�^�?�A�l9��gYg0qƐ��y+o��8�4���ݒ�7���+b0F:w`.���2��s��l�㒗T9R�=`��]|����"��ʎ;��r��aS��5����S����<�}��*ߓ^ꑟ�����^���r/��d�梆�9y��.	/jA�rS�2���:}y����z��L��-Y?��>�Ջz.�����u��#|�E���Nn߁/~�C���쿀�tMdX�ۧkْ#9�;֏p��nV'��^sW�a=�Fw=�s�2���x=o��s5f!.���;���@e/�l�P֟i����ՀuA���8A�tJ+I�<���IZ:{]6}�wj�Ȧ9��4�K-�ñ��u����{��5gs�.��ʵ�k͹���Ó5��5���m����uJn�%e:�2���N�I���B�x%����T�ϣ�'���Y���kG��^Ck�a����~�^Ϩ�����2EKG��5��������?�4l6k��+��O��������t�tk`D�G����\��w��`Ƈ�5�=��8"����:xᓟ��>�)��-�2���W��D�����������/`�����ȔW�xh�8i��v�eJ�,/�y�Tߏ܊WZV�#��װ�7C�/�T<83�3%@����tla�03��ܐ�!l��fh#���]�>:��_W|n�S����zb���l�v��iT&�4�.5��s<����H�D���6��w���N����$���<Z��)\rd�^CK���p(wdy�
�*����x�:U�a�;G��/5�F]��:
?�έ6d���o�>��߄�>�~ ���\'n�M{܈��h�� �C!rTR.�j@�*��Ō�.��
�8=�P�_�骔��t�����ڤ�S>��}g��qɋ������N��;���̷��#W�Ƅ��U��G��b�{�6���߃7}� ���ՠ����9���R荼�T����W�F�H��U<nt��(\���![3M>W�����f(���Z�P�f�(llAYNRbU�xU��}!�r+c������9��'WMs��x��!�G3���N��`p��f�m�y�UDϻ����6��'�\��<��W}�U����d��c��JO�/5@�Lw�Ns���N@g^=5+*m���T���`4}Ol��a~Y��"�1f��*�e���B��N���>���6�5E�=<����/B\��Y=��2�e�Kub@-yK��B�12��׍>q�^j��p�r�����#i�vgx�?~#�:]�/Ǵ���t�ٲ���x�)dY�G���9�qV(m\�~ o�*wx�:��n�O�7����?�,toy3������ALﱈP��o(t6����S��m;y@�N��59A��3ޭu�zL��H�d��b�7\1�N�0���d�]�[7D��rQt��l�֖Ӂࣚަ���^[6L�����E�e��j:x��sN\�{�4`�҇�<N|.YM+�~�����?s�5M�ޔ�]��8^:Pٵm�V��I��;ivV	L15���hu��<�J��7,��^���F̃:�f�v��x��3x�SO�~}^�Y�u��c����1k�*��t}��=ց��V���m`؉m	SkL�Lq�����A ��[���к/� �|��໿�/w� @د=���t�Z
�=�!�� G�I�z��*�}Y"�r�B\�ol䑍�K'ә���MpE�U�S�� ��稌���&�)*����1F���ĈeP�ԸQ�J;��jEW^��Y ��O=^&�4��IU2��qoec������s�0a��m\��������dΜ�![�#�7��_�L�J�Jgp��`��'dI�~���ڨ�ǋ�x�=3es�`���F�Qb�Ϲd�����ݥ�
>�7:7�֫l`�����?���߆�m:X9���}�,{�L�Le�h1��j�a�V�.7�A6��
z�J-9�R>�-��q��� ���QR��uz�R��[��w������u�����DJ�fV�Yn�uj��Q��'�\e�绅������A���䌸���m��?��|�w��u���Y�8��fdz=�$�����1����_�#��>4�H��X#���K+#��Z�*�f��k��	�S����l�������9��.v]T��"�=c6BA��lY�^v���A'
��u���E����0���X��,Mc��������r>k�_Wa}t��t.Yj����j��'�DC����T�M� rL2�E[������ �X�r�M���17�g�t#c�4C�������Z�����Pox7�7>���Wp��_y�L17�
�5�K؁ÚCB����R}���A��X!I��?��OK�+��-�@KY����ܮ�դB���ߗn2��@�u������90S;^�i�6?��[<r�٪�d��%�>`�� _�CE�b���I�����������|FG90�:8����?�O����M�?�.��N��� 綻b�.]����r(]d,R��l"�캵#��佌ه�,.[U���:U�� �u����N1o�t�\��)�ZM�L�ޣ� ��T��?���'c�M�7v�[���J�xzI��z|K;�����`}K�����J,=L���9}�4�rYǍ��m���W�W[�u��jk9�fOF��P�χuS
����ÇpAʛ�;��&}Ae;�8:׉x��oyG�6�����O�7G\�d�p�[D���t)K�q�s����uż��K�W"f7rGG\y����$;<ڸR�Ɂ#}^�l��q�����~޸Y�&�Ë�z1⣹�S�os�*�֗��@�P�$wl[��X郵O4�N�unO��!�����.����u8��?'o}3�����=t�5��C��i��j4_�&2׫ c@��}�f�Wmж8ݠl$��7�_5Xp���e�Yko-�0��Y|�ţ��9NN�1D�
��B�ŌlR�2���S����Bpf�r&(�3�粇����C�/F��^<��ܜv_�*�c[�tSpr6r��l���C6n�c�\@��N��1v|��p�L��L�.kH�c�oE���g�\֡rj�U08��?��U�����Ƞ��r?�F��_
��s��z��n%���v����>��?	���B�V��' �@�9&� �6�g�
�jH)
�2*�T���)%|I9K~?���9]�7�T��Z�GaL�c2�S�9S����?W^Ki;��������ul��X�1
ZeW�������ȥ١��o��� ������3F��}��'yH�� �Q��c;�}nG+q��� �7���bGż���8S�k�~���ꄇ�u4�nqC�#��;�S]+���.�W��m��Yt�hrʳ��(́r��K�Ӵ�Q�g��5��E�8b�G�}l�^a�Ǌ�O���f��$%� ��uV�2p�g]vu��pw�볦Ste���1٢�qQ�,O�O����(�%�EP��8�$�+PɛNjg�d�LS��'�5���;�:�/��Cp����֠��n�oV<��v�T����L4�r��J��}�G�)��)��[5ۖ��e
��6�{E?�:Z�<I��j��KˉO�����N��k���O����ب|��T�cj�rj��?6�m�F_)~�\�F+�8v[}ٰ��D�p�J!�d��7]	v�~��W�اM�A��9ץ��=_�1�:�m��:�@46_�P��O�T
�2�^bve��`kgppEF�%p��*�˲i����z�6�I[���}�XH�m���u��\���.i�갶Jȍ��*�9�߬�Ͷ��n��3]��{W�S��e�[�^���ln_E��CN�D�8�l�B��c̞�o�_��b�{���kB�#gT�K5���^$B^�Rw�~�{�̙�G��lW�a�>�#���ì��N��ɦեK�����޶�[{��w���=p7�K� ӟr�oI&N��W9��s���l���4�����A�_2�a��@<��{����G����������n"�n7`3��;V4��O������{Ry�B<yy٘"Ȕ	DY�d�� ��鸀�e攛�r�(��gf�g�t�1
�l�c+�l9U&�_�Ο��Ʉ�R�)��.F0�%� ��B_#��$O�6y>�9dt*�*�9{3s.�#�$,`;XPQy�^��%Y&���\�8�Fs!A2d~!3�]�ⵈ9ݸ\f���su�_BG���fܚ�pm�S�v�Mk9����{M�K�9��@9-6�K�������pAV� ��t�q���N�>���qx�t/t��26C��·���=������۶{ؼ�&l�	�t����FVQ����'(~j!�1a��Nq���sFG�����W��V��a���F�/�t�Y�:]�G=]f�c�0i�O�g�amn--qZ;�N�է� /���v��`"�M������� �>3`�.�D;�?|����9�ƿ�Mp;��c?����̚������"�X�G1���R�I'�}�Nb�1���j�l)��1�}�"�iYrz�#�A����t�� �),h�MOӞ �x
��j�����Z�'��j�`�<�ՙF�?J���{�T�%M��\F�\E��j�Ee;�Tқ9�u5��R�c�uZ=�m3�]R#�I4 ȫǙr-�dS�=,�ɚFK��SЛ��E��*R��E�p`7�ڛO�<)��8��kAg�6b�N�%��4�Z��O�u)�F���պ�� �t���={�`s��n�`���t� ��s<js1��9p��ǦB�^�XZ8��Q�3������e�T�ݩ��0��ɉ�9�����:}٥��b��]��+ʠ�&˯�1S�g�v\4��Ŗ��,r�
�'�Rd�v��f�.��(�����y��r�xr�`���B������>���Ýep�Az�}qtݪ�'��\EqCdG�F7�r27�	�#�!0�v׌�~2c䋤squzD6�@Ǻav	A�������A`=�v�V<h���FJ����IѫXt�8�--1e;�8@i�hʮyU�����H%ot�s�s���^����Ĩ��]'Bw�@Q�^�F�gW�Δ��g}܉�S�|�f�����1��� �ˎ�ɩu>>�.k�^7ϊъ���D���Ԉ\�X=����Si���hfԅ�挎�%ǌ�#ٯV����G�c?�.x� G���Z`ÛK�g�x\���8^c>X �����Y�
�~5,�m�O�>����
_���E����6�����=�V4D�Gq�!��S�x���C�U	�OX/M�y|��t<Q!��H���"��_ma�rЌ���*�������b�%k/�o�V�81^��Fb��~WBF�Fl3Q��D����g�cd�(k@KP��\I|3 ��<Rn�D�~���7foA��F�e��d�\�Yn�퇀L�~��)Е�G � ��v��Ok�\G���8cd<��Qg��rQ�`0 d�f�1���`rG>����t�d�rW"��|�צ�x�(;-vV�����@a�6s�.T�� 6.�v������џ�9x��_��jC�'�5�	_�Q��jM�Lk�,a�ź�p���|�s��7��e�,��n'�ʘK�!+=����g���p�X��}�r�t�p�`�k�^��^�qޘ�3-���!��s���Iul;��ο	6��6��HU���ފ
u�ɧ��t2}�lx
�����}�_�"�7��c��=ޜR��0������'TB�Gڅ�9�k��κ��)e�G}?����%:h��rG�X�������9QJI泞� �w#��PT0�e�I�`��
8;�.�S&��x60�┉����lc̵�<5V-���{���ǰ�Qs��C��_*�f5���U�f#��>���N��b쨿�nCNA����C����LEUez��b� �B�����83�Q��$�x��ڲ�n�ZZv�v�c-��!�R�~�Ǒ/������=K�<��;���k"1�A}ٮW��
~������.�<���ԅ��13](�h����g�j�+?�Z�}֡��l|K���-Fֿ��Sx�u?��Rtչ��uԔm�Jq.�NW�����:f_��%��`U�s�b��U�^�]�yHǺ���jJ���N j��@N���˙q/���'`��اo��~��FX�+�~�S���|�W����pc���
��:�t�N§�@���:�r��rs���:'C��\Y"��g����X�}���˶��`�\Ͻ��vm8��E7��������쳶������Ys;@�����%���$��a�L�&����ô�Dk��G�Hjt�X�7�0������3�h���v���[�k���>	d]��u�uR�ؼʷ���n��F�C���e0q���#dh_XG��u�n�H�p��i�N�I�C��'as{���[1�1��#��/�=/p�ʸ����z�Ik��9CH�"ZDm��y�Eq��Ja��cN��}i7�p��/�/��߃����3�z��ܑ�F��{�nP�lz}
��	�=2	��ʝ O2<�"�Y��G��%��V{���ф=2<�<�o0�xQ�aHɂ��H�W��9Z���J�������`�/��C��2�-9e����w�Ř�@A��^-��XS��^�p�ⱽ]z���EF`�Ϡ ��1X
��+3��S 9�)'Q�}���E9�P?e�-���`
F��[)(u�V�������
�i���	�+/��Άb����� f�y�]A�F��Z옾C�vt���f��*H��,�=/0�NG�.���|�ZT�rR��6�R)��.�v��v*Y]���B����Ra�|�V�z��'i��>�s��e#�f�m6�����s[i��� ���]nb�!��@��z�_Q��n���5��`�n@�����=��O�W=�V�$�=��R�����x�w�� +�1]*�0��%Z� ��c��NG���"p���Q��I���^&�z,h,�� �z��u��ǡ�.2.��^Z�1��(�ߗZ���׺��omh?T�!��9^����]�|���nø�,u"�PzI�BT-� "fp���w>���N:DP�9�)^�W|;�#(i=��u=*j�?��tu/=�|��o���/&�&ʸ��稣��0���;cl}�M�����	��Mdkx�f���^@�$d\���}�T�=��>��d�\&��:�bq���=��tx�Qj4ێE��X�㝵fc�qZГڕ��e��%��&�c�10�r�-�!��q��I����r9�?�м�(>�ޮ)�9��d�g�{,�
<�c���P�4�n�k�*M�&T?`UW�^e�J[j�G�T.��;��f�<E�����
���(ԫ����6��O��7�I�$zk&w����8�}'����hG�z\T�Ӄ���8��;���W�b[�(A��$���rn]b�ʮBϪ�K��/4[�����#_Z�W������%��#CY4�N������F���`��0�5��t���0�~���M��+�w������:x�
�A�I�SI�uF��{jw�Mf�K`�&�I����\��a��Q��:��m�C=7��S߭��x�7�R���O�8�0�$mL�TǦ���:�=j�rJ�haB;�s��K�Et�k]�j�ei��\%M_t�kݧ~.e[�S�5E�s4~4��4�g�"�G{ h�9��8o$��W���Z,$i?��|ޔ�
 ������9�ɩ�("�����s������>���/�+o�F8�rq���~E�;����$!�Q��ka{[�cf������@����hw�����H���A��RU/2���g�Q��{��r]>p�xǕ%D��'&_��^)zS���nA�bׂʶ;�i/&J��z,�{د�K�5�)c$��4JOf�s�/�>9��G
�}���c���Uw�~/�(���b��2��X�|)f���5��q/z�>w6 ���LM�Z��*ʧ�ua���#�m��3|L[l�R�U���c�;5��}]?�~(� .Kߵm�rv�k{��F������>�~�"9��7���2�1+��S
��>�~�X��j����N�����z՛/F�S�~9.�<�l�h�{(]����L5 �$�mֈ��o�%حX ��_����'����Wn<���ݵpDP?��=�� P�dS�I՛k�8��)/0���v$h;	���p����C�#;'"�? �ql�^`�'m�|$CR��<���4�w�Z�m�s�����81$Bƌ)��Յ�..�k�Q�_2�1���\8��Dbb|�8�ż"d��.�8�[^�7l��fj
r!FU�D��z�m����bc1f�M$xESWشc�cR6Ʈi�*�A���(��G�hT����B�J+L��D;^���NV�3���k��qn7_�u�Gū��2^lB��Kn��%�(�kY�D�1<�>@5�{.�h�/�:ޑ6��i�<�7�R;|�k�tn��A��6�����?��?�܅����N"���n��D�K��Rg�kCx�����2	~ �;���8k�3H.���Bz��x�u]U�1_��K�^������~n�E��<(g�z��R�d�Ō�r�`_���I��7�FL#�'ZŲZt_�Jvs�N�xG2�d�w�}@��?���'^��_� |���w48���d��h�L�aY�q uӖd�4�����h�*��*��F�l��Z�.�7G�,����[�"X}�V��}�V����fz�h��'����u^*|��gtN��Y����A>��[�ٸ قj'�>e�<�&1����+m��7�;��q�#�D$ȸ	Mcwe|*�uɊ��<����,.)|&!��UG%��~�FE|�	��q������f��Ky�_L6P�ї@�>*x�s���d�Ef�ɉ]�"+�W9:FCvl�p�`6��t���������ָ�+%�|l�������|J���3y��9v}�,Fr�A�5���0h�93mƶЉ���$��a�8n�ꍈB�IT��܁���y}�KO�"��7��?��p��/����A��8�I��jH��Ďj!o'��~�W(����i�l�*��Aj�i�]s�Sxbjs�N�f�U9o��nm\_���0Sa��d[.3��:�k�����i�y��2ן�Wk;�rF����G��>Q!p����""~���B� ��G#d�'��eL��)O�'���k�9�V�{�{�g���w���擃�ݡw������t?<_�P.}�Sm�-������n���|Qz�F���ܖ��y�XT�hSy ���w��9^�-�!�p'��8�� �� 뇶�ȥ���!;���i�#4
�<@�t(���9(t^�RƲ6�a�U�ֵ⨜�q:�[S��T��Cݸ�gU��D.iD�E���( ��ȵq��A�����V���Y���� K7��'�Af%�h�_��
SKuF%pE�5�z��#���!�w��	Vp�C�ޓ���ư�ӵ�)�~�qn�ނۿ���������Wau3���7�K�s���C�{Zf��MO^����S����|��s�c�d�Z�ii?'��/I�M���=����������?��C���r��@<�p��|�,]��ہ��{6f����R(�2�p̤��0	����<��G����BFb��u<b����[�&���l,�6����猣J�"��yΞ�b��(��@@h$�M�/OO�A��Ǻ̝�N6T#y��@���W \�K/�4xa_�\����E������1i���T����k����F]�K��jV�c%�y M^�9��S �[c�Ae�㹷���;�Q4�(�Pp��voX�J�J�ۓ>|���.����"��2!H�5��儝L_�I��c�����b[�X1vi/�1����!;=�A�tth��_CWrtC�_���DKa���A��^���X?�,|���Qx὿��O�ɴ=�� w��:�y�!$MÏI����@v��2��ϧ�-�fǜ��e�����*�г��`��0Ώ=<
m=�Sk��"�39��(�N�j��~�Ei���F4�'9X㑃)P�#N�t�v4�Ơ w����>��u����»����"|����ҭS�}7	�=�O���A�;T���Zڼf��YFA�̿R�Z�8@�D�nGй|m���yә�¶�ROkʍ��V�xX�:�k���6j��h�(���+F9p����!G� Z���(�8A�Qj�.j�փF��d���C,���B����^�c����q��W�a5	��̖k7�m4��aM#:N�GF0�	����|:�~+N��\����#�a�I�6瓃(�o��(z�[��d��w�g
����cH��l0\�8��ӓ��e������\j,Y�z�kÈ�چJ7�z�D֤D�QD��j�Qr솂�X���d]�8t�w&]&�)�Oa?r6��'�|�}���/���7>��!_w��1/���3I�4����F�L�i�ӕ�h�E�Y}�ŧ����cY�7-�g7֎u"(6�*<YG�lj�Uk���������^�C�T=�r��q�du��o�g��a�C��J��ɹ�s�k��yۉ��v���F�u8���-%��́��N��Y�����{��_����~��ӯ��p����O�&���Ч�A\�	�2�Ju���=T�Xգ��
����9��g"��Ld�k��,=@�Q_�����m�b�X*�ڀ���	r Gq�gG�����\���#�c�W嘁�������:�`[>F[��h�#B���W��Ȳ��
A����V>+�G1�lE�5��j�T��5p^kQɄV�E������:�3c�m���?�8�)�)=���Bvu�h\�(��uZ[�[��N����,Lr���g�T�ݓ	q����[ҍ�v�3�UXE�`d%G��;�bq��+��5�����>��?���V�xjpMARt�����֥S��B�e�$�E���%xEi��M���� ��l,��N�`�؎�B�l��ց�?�c����3�m��+��v��BU�$�w�>�A�����w�1䭆��`��!Ӯ2�O���I_Q���RH¦Z��z�+��<�v��q��<�\7�`�W^�B�Qȋ���Z ���*/Z%5s�<�RW.��
l@��ȑ V ��8�r��
=��a��I� �8�0Ir$Hrs��U�cNnŔ 4ƫ����v���
hc��e	2b��eX�i:0SNm���mo@	�ӿґ\G��!���2c'��/��P
�~0lm��^
Ɉ��$G<�D�3��+�*��~� ���лtOi����7�6U�B������Va#��`�Rɓ�v��D0<�hc��.):��9զ��7g�?9s-Mt���+[��>�!�O��+�^��������Oa?�~����_����������~���܅�OB�Nl`�9M8��x�z'\#=.d1^Kwm��Sl��I����SmS�ZF�˴��Z}�z����k��S��m�*c��Hs��JS'��{��ֆ���,i�xM˩�G/�s���멹�����|���v��ط�:���ZJ�M���r�W���b+� I_w�O2n�� װ�{�y2ȹW��������~����߄��B��0����͊��X}@G���X�y�h�Ó�AO�~֐�bp�2*�J�r�D~���Tbu���w�}2}f7�E?iѥ��Z�1��^0��x��b>.���W�$C3�,4��+�F���}�21D6c/�0o��P��La2�u=�M�ox�`M�:G���`�o�`!�fSIt�?�7z�J�W(���S��䚵��b��u]��ݢc�a_���#]yDz��5���'�G���b#��E�A�49`�t�l�=cl9%%kQ0�"뀯N$��H��G������!ϥ_���3�},F�2f0�5�@|MWFy����_�cOK�
1�cR��5R9^�*�y��d��Nzf�B�3E��w'�����]x���O��?�7|⏠�l�>�٭�y����ȧ�
�[:k�.�%q�I��W�,s.u:�T~�xo9����p�[��i��a�Ci
ߴ���q�$�S�i�[<;����NS�V���ҾO�Y��.�>�����r����ҋ��ε�A����Ӿ�S�a?O9���dq�5�e�.�s�9ɂr�VE��Y���k[��c��|����?Ͽ�W�?�4�����[��[�� _Mgt��`�	{��C�9r�DCd�[������#���hLuy�q�chua}9j���APη�KE=ݲ��M�t�q1Ǧ��Gs��d��z�����/'�P�?���e8�u���� ��.��y&+UmlS/����$3Ϻ�+Ǔr����?�&����q<�\�� ϴs.��}}� �#OV�g��X���ܒ-@����<���.��ړ�:�/�XX��r:w���kq�0������{e%�ȗ�@���� Ⱥ���77��B��h5�[n��0V�ޒ!y����'�Ƴ�����?����D���z(tЅ��ѓN����{�0]��&_��1�D��E��8d2Mc�UA�ٱ���4KX��d#5G]��^I}H'�� 4`~���?�/�=?�n�_�8��?껾���]���f���0���������PL:��E�Bb ��t'�A�{���� �Ƕy�<�F0������g��э�'m:�!"F�,���\��*���N�8ƣ�����ΧT�~�Q�2i�z���#�&G��O���F'Ԉ�u]�gx+�I������;ǡSg�<���zN'Ŭ?G�� �fr���[���A�3�dX#�0LR�8}�H���?-` ��g�R<���F���,\:�Q �q�#��*�"WtLC��<��]
�,X������LON�&��I�A�0X�8G�����哾N癣���t��IX'O�*�:��k����"lS�>����u��9���#g� �����)GH�Y��.�4��^0]g8`�5�ͩ$��\v�
\��܌�(�'�]9>�6y=9�GBX���촡���IRlbm�� hCG�W4���M����1�~X7��;ф�����Ǜ��m6H����`��߃g�=�����p��g��;����C���=YQ���Q������1�5'OD���MU,"3�ԁ�nP:�1�3��^D�������JO�C�S�FQ��s���m
2�^���G},[�̫��p��ե�<�L2�K���˔�Y6�V��<�O�_�,��i]�P*\����o�y�z��U����r�#�I8L�rb���爡?#[ ��d��NO�f��� ��k����o@x����k�,��o�v����>x��~��o!�W�0�n�?I��A0�p?���!	�"�	�tүI��R܀��1�X�5�i��En���`�$���W��ɼ�{b�����:v>7���܁��������R�QE���H�Y���(t�G�2>H�b=�4ְ�1�����=�u
��0�9b�퀍�p�G|�	��7�Zu���&���11⑾��O?��A�h�����J�Q�ZȌ�=�K�ߣ�eB����5cuGV�T�Ǩ�̳�+𩯞���v��E�7x��,���l�Ι���('�p|���!�����8,�nD�<)��ʓ	��R<u��R�2NWtx����4�{Xu+]S�2i�`���x�R$����	�u�����b��>O!�=r��$��W��"K��n�Wّ���G����%�m��Cy֧� �de��J��>ґ"Y[2��7b1��ϕ�3+t�����+�����٪sp�������}��������x����֯�7��[ ��j��5���q�c}��10]��%U����f�>�%�=�����B^c�5�����F�}6j�;��%i�A����n�T���+�:[�~)�9���ϗ���}�m�_U)�Xǒ�"M��ό����uދ7��ƴ^o*�&t�1�S��2k�V(�I��*?�>8c�5����2C�ۡu$:`�M���7�4  ��IDAT���n��^|	>�w����|�_�~x˟�Fxi�������Ч��B�i����?3����H�����=ׇbLʿ��>����l��5+'^���=�V�K�gӮ���K��{U�}_�f�d�~�h����x��<2��� �%�K�+s~���qM(6�U���P_�8z��U4YEh��zy��x��x�-]�j�b�>UDc��'sS5a�_Z}�kZ�KsM�nu	0�%	٦cEʾ���6#LM����8���9������9
��4�>��/p��Q�.�ZpE��Hu�~��j�i���7sV�2��}��� ���.X<��}�wy�c@�4&�m"���E���f���k<8}�j�XGX����o�2�����p�c�o����|г6�"�lȩ=��l���}$N5u6������R�oV/��Ch�o��E���5*d �<��K�[rDCL���k�QGh��3�<=��Q0��-vg�����Ξ���g>��˟���������o|�����u�z�&l7'pcs���d���NF�QBN֧}Gr� �fC@ �6�O�"!c�X��/�wʓ�h#�H�]�� _��W���&�����п>����r=z�?7�𔍥�Fڤ%��S#����A�������_��#E	�{8��h|y㛾�gdtN��N���>���0G���(��4b<
����L@���|�Z���2�}6S�AS�'Ԥ��=�%�P�f���S�Ԩ��33�j��Dv��
@�'��z�A,ѳ�{ơJ��Jc���&�U����B���bbW���JQ֢��p����`�ks�AiH��랂�w^�]<G���X����~�@@a?���96��8�a�w��BB5En�Ӱ@�ȵYb�DǇ��m����\���=-�u/�!�sl{�uԛ��G�~�C��2��H�;)�?xb��'}ĳh�}�x�ʲ#Gq܈L���v��{��2���O������{6/�7\7nm�Q���Rح5�c�0	5�
�5z�rV:�z���Ƃg����0\s�V����iIESUiP7��{pL.�挭K޵��D~�<���K��T����E˞��07ԗ�9z�l��qr-��QIS�l�[�NK�*�^f���%����/6�)�<+
�� �p�P:`�~{��uR��̚��Z����A�q]��͕��6�f`7��;/=���3��_�E��w���w}7����sp�U_�A�q�>=Yc����c��������7Q){yc������9���ɸ����/cݨ��WUt���0�M2T��_[b6�.;�{1��S��Wp��\r���V���s�U���"�d<m�&�U���`��B7|���M_�؞oa�;�C<�"���g���xÉ�$z����<ɐ�O�{��D�(16~�:hd'�1Ω�u&kWk)��A�4㪸���k]B'}��I&	����!o�B�.	1��N����{(���ဢ9��f�I��n�v���Ԫ��(	 mb=0z�A������kD���ӛD��C:�5�j�#��b�'����O�]�'�x
�^}	v�-�7u��j�����@c�����k�x���֓�����i�w��F,'�T@XޱC�:�@^�j�z���?�Cd<��Eֲ:pH��u4���9�Ŵ��Yz������^,v<�Xr��F*�."'�3m�A�����9�y�s��~�������QX���0_=<y3)�ül�����Q� �Ǉ$\^k~�b�C�#��W:�	�կ��8��>�k7G[�X]�������a���Ŕ��\Yu^��,5�����5�f)�k���?fl�1����D��z~h��}N�y�-s�bil�Q��!���9v�j{�!^h�k}��#4����a��Q�;j;���9�hq�s�@ܴ��Գl&��fd}�dT�$o�#m�>���[twp2`�-�za����qx���=	����੯�*��)�v��z�@27�zň���#w�1�N�Б���D�ٞ0X��"��[xENC���;:�.����꼓�e��ıV��f���E�o��A`��A-H�",O���V1mP��E}(�/���b�܅�������Ox�z|�G��G�1�)>�e���T�諮S̏u� ��i:�7���\F1쮮�[�0Vs�2;ۓi�qh�붗�(=y�;�`/��7�RƳh��:qߋ1dL�Z�kAl��x>�,�^5���|�Fɪ�.*;����*�w�����Ik�����Z�G�k׹P��rP�}9*|><�Z⍠�T5z5�q�R缾��xk2�1ͺ)U�U�r\5s�U��~a�x��iFޮ$��G{�'>){vA�q�H�I:�ܹSX�;�����߅������{�7_z�Hk�$E��d�`�	:���<�v'���o��9/n'5:�}V��"���h)ڞ���s�)=�.���u�I�qT���k#�d�0
9*�^�� ����IXmNᩴ�ӽigw���<�k�0����!����P&�]on��wh��,�ٱ����OҒ�
�v[�3W*�.���P��x^�BT�u1���KJ��,��(��NDw��HT�|-d� ���|�
a2@��IP;2�tg������������ ���p~�l��HK��I~�x��8��Kx2�u��Eś�Z�A��$����I��NV�ܱ���6B��x�H	C�h9�-ـbi��HE<@�8�\�aO#ɜ����FN4��N`b� u$�DE_���I���i%P�V,��\�3��.�d��8#��{g��C��zg�r���q�p� ��plȧl��g�[Br�t�d`\�ƹ�;�
��O�����VJ����1J�VD+Ƈi�����hڔ��=���<p&���WE	�,cCs�����5�!�v2�F �r;�ׄ���]�=�q[y�G%�{��F�# �O��Ej�fP�z<����'g��<
O�q��_:����ݠ����z�������������>�5Xq�O�nM|�Z��W6���(v��Q��R���I3��s�t
�����P~�ˌ�oT�h��S�͹����VZ�,Nm�2�L��~>W�E$�f�Σ�����E�Z���4gl[JCK�?d({�Rm��Sjj#�ܦǡ:[�(�M���i:�O�T�n%C�Sq	˙��w�ix�N
���ia�YY���f!�B����ި�3ڭ{ė7��oƛ��G�
�����hd!�d2d��E}
ey�Њ������8���$�@�֘�Yn�f��G��MEQ��FRG1L�	���\e��J8Xt%q�Ǩ����|����H�T�6J�RJ學�F�Jy{�?=#R��y�N��=�����������߂׽�M��z��W\�E�D7d<��Z�@�#E��\Ƽ	��AE�E�3��b����W�<���Ϋ�V��u���P�9*&TgZū�
ō5��~�������
Cŋl���H��x��n��'��JQ3���XZ۫4�j�ԏ�s��wysD����J�k�K5w<沶h�h\P�
r�(�Q�i��=�7�$��������]��o��ş��[�iL��te��t��
D�g�c�,a3<�u�tt�OzΞǆ�d/��c�©'���cd���M�qd����z�r�)[NlE����=�-E�tb+�!HOHNn��x~0׮l��E��"Xw�:�$2#��i��O�9b��ֻ�Ϟv���L����P��$չ��t-p�&�Bud� ��i��|C�����B�F>��fdнܠwa?�g;@��Bz0�kPc��8�m��g�Mv.�l8�ڰDG���Q�)�P[�T�8���� ���*1�m�ݜ�it��C+�h-Λ.���hg]t���b)N��ک`I?n�z�gv��v�,q��i��%{Z�3�������6�T�1 2V���~�6V����i+�<,]��z�+BE�������n�"��f���� �ׯ����O�?�;�Ư�zx��Vo{t�
No}���YA߱�2/����=0�;d���R��[���V��Ts)8M�w��6D,�&�b��ZӒ�a�~T�1�ڤ鷠��b�u._��NΨ���7d	�
��"��B��K��P��CyO&�0���%��w	�E�E	�aQA���n�+�	n��BƕÈ4`e��<_��v*��G<w�~�{���8zч�Ɖ�#�:적Xk�9?p���6���9���M!�oU6�_&��h�X��2�S�S<�3�6�>�j��a�|�>�'0PUD'"�w�f5R�YW�D��V�-��"2N�b�YH���A�6 �P��{����-lb<h��-�T~�U����L:�:hKk��+��e���ۀ�.>eF�T�����`{���i8��g������GO���W���p7�5��g�VuG:FڠL:���?�'��'x��ְl1(�<��9p�(��U��J��l�%�pE��H6�h�"`�����^�����iON=Ftp=�Ѿ'n����(��!�Dp{��� Vze�T�z�eeI� �M�4٠&'�=zϱ��P:yPy�'R��=_y�����/�D7�_ߥ�U=����G)K�N&���[%��	l$KWל�U;xs����7�����08[�xG�=�]�
F��,�8hx=AH#�'AFxP�[W��+����&�Jz��+�Z���P^
YgO�$�i>��>�\ڨ�!p��;͜��cz�H+0�ʃ����lc�(ME�.�b�p�|�%��s���l������=	�4���Yh)�b ]����V�}����~�b��o�jx�?y'�/<�����I$aB�A脣���˖i2v NRQ�������a�$f�N�4t0�ql��@��tJKB��`$�|���Օ,Ls�����u�o�ҴD�F�9Q�������K4+r =O~�+ޜ�O�8L��q�6�oJ���M|����	w�y#
�1g�cQ#�$s�NBO��ه�� ܹ��� I 8ȁ:t�2AA`V�\�l��de�ޥ�M��e�8�=�6g�g-C�Xٿ����I�6 ^�l����ݾэ�N1���i���#K��=�LS�Ġm��s�gy[+�������5�Sm]:'�	�r�a*uc�,���<��n��� C7ka��P�7�/c4���$����8u��<�=��_y�ÿ�jP��|7O���Q�-"��G�.�}���`�T�6�/k÷tv_���ƍ����[F��ng��m �R)7�_ �G����!1�y�4�)<@<��k#��(���Wu>���Kt�L��jb�o�l�:|�1��Jه-<q�%��?�Vpo���was3���&}RB�T[T��^p _�����μ��Qư0��A��0:�٢G�I9�譥���;�LOo�N4O�:/y�c��a��'�fR��D!u#r~qr�S��uC$���8 ���S<fu�W�����+��h^����^�W���v���q����݈��������#C���+mVpc(����+�Р�|��OE�H��6KdpY�S�2/�Y�o����[-��1�u�N���E>YoIЌ�̨�t���.����(�A��3���е*��v��Sjcb�'ǔ��;:p�8^O�I(�TΆ�K$�y�D�v��S��1|X�a��ۻ�N_�IG�L��]r�����	�����%DB�h<��`I��Ȟ��ܻ��A�c����X69un��|X��z��f��ЗK�ӵ*<?9�������K�I�ct�9��ؾ6��X� ~T����{�ϗn}L���׫HS��Z����shLCˆR��l>}NGc��S��E����\���������4�бb��k #;�\�%PO��l����e��G�B��H8<�ޟ������\��3��'>���)��f���SX���!�/�A���t��r��oWE��2f6�~l��|^��3��8*�&q�a�:��E|)~���A�zvef�&8ng����1��T��?K�^I�n�N�����뛿|��'<��QH��= �,^7�M���T�]���	c��q<�M����^�ٔ��{8f�,�:- �n�j�~�Y�͟�٤M��G6/��}��kԏ�bh�Uݼؙ�&�,V_��K���7(��|X��G@��ԿUǇg�O����-��ϼ>���f�;�� �źE��=�-���ҌU�Q��a+h�C�~�#�6��+�ud[�U�T�+�E���i�ˏv�7�q�O���U����>�#F~������>ĻgC�s8���������6�j�${��[wx�خ��{|^���[8b�Hڕ�����F;oGV}�G�cXg~8�8�LVP�����!��D;Љ�ܑP���1�I�`�F,���ǰW!Sϊ;fc��K��S���0ؐ��h�C�ʝŽ3˃�*/:�922G���´�4&$4��5��k���׸f��ñ�w=���Eb5��^�u�?�r��CG�*+)��#9�>_��<&d�I|9Šp�{t������=�::y�����J�i�<���x�gOt��	@����Ȇ`(��L$��'	�9�E `����
f�ذ�cE��|v���&���Fʣ/�)9�'�M�	�.���A`u����,�1�h��1�`�@g�9���ØZ"�p��}���5�;X�
�RL孀A'�q�"�\�����\Ԓ4/�eX��C��{ђ��J��@/�Hk7��K@����EL�+�>�7O�9@�B�t~�yV#6�Ok�C�U�k��Nb=^�8��9��6$'�#���xp��sX_2X�^���֑�9vD���`<9��� ���#�K2O@�Éz@�/Ȝ1s���"Th���@��t$^Ą�q����q~�g�d�N���(i�����8d�&+N��c1o�T(�,�
��T���/����	��ep|JQ���������Ƒ�χ�Ƚ�_RN�����$�0��N�S�z�vjc��{m�x�DKӔѦ�-c��M���!��!ڙ��A��m�!���v��q�*�Uϒ���`���>�4�dݦ4�M�%F^1ZE�:�L�3�޹y�x����k'#qi��U޴E�N���;w�4a3�W]@���:�(�.����;��*9ƻtnx��w�o�^���$g{{�-�U+)s���O�� �)kJ$L���$i7a�q���e���bQ�b�t݂��d#��s0���`d.7�8 �l`r��N�3����q$;�S)r��]b���yC�����{u�&�LQ�R�{��i�"��\�7t�'���s89�Q���d��G��@����}���D�٪%0^mD�O��J EI ���1N��,�ov����1�֔�:��^�<�}ds��FG�Hz6�:�O�|�u�"�Y�"��bO�{$�5ӕ��|@I :SjOG�*�ҝ)���q��>��Ӌ�!�"�lp�֭��<�0VG��.adCv*P� _[ʎS.cl�f)��c�2�����ul�`��	;�Lr6`�UZ�c}A0����w�S��"]�(R���1f��g'���{�`��U�����NFc[Q9�� ��G勸~��/"��F�^s��׹���)r��_>��9�m�AY7_�j���|�yI	_������L:�ۥ�>�V�d���j�A�G�	9��'��N��4��D��80�CVr@�9�}�eH���p\Y�%���,�bD��BCص�W���{ c�\����dy�m�3zlK�Y�Z�em�~����r��9
����k�)�ȶI��Ni�vN�in~��sy�谗-;�%s�D?kb�zL��9��^xG4c� Z�HS�?g�xP�|�.e���JV��K����|��m�z^kݱ���g�D�O�ci~)?�k��f$�6�u����].�G8&�'Y@��{v>��=�X�rO�A0̲�^��l#�"ɉ1�<{۟���I�Y�}k�0Z���ó�W^e���)p��q��M4Q�i|���t�WBv3_���N7��(Қ���b�um~V�#���"�Mh�.o�ʆ���Y_�q��wAm�Nt ����O�Q���`�PtB	�>���?����'�����%���Cs��i;{�M�A._�]}�����ˡ�U	�U��
;A�T_QM �[�S49�2�4���½n+�uH.�O��������;�|��!�Bt:�6@���(�R=�=��z��ݰ��Ӱ:=��=隞�[�\nǸ[+��M�u'�e���^"<�O��������B̮�z�O�(��1P�1^wr�-��ܷ���<P��QU��畲��'͓�I�{G�2k8�m����_������=����=�8ִ���e�N���aa���s:��G�bW�\�����؛�7�4�nb�g�E�� rǗcB�tZgśӸU.O��`,>0�� H9���+0��!���u,��~�ʍ����N� �o��τ9�I�q^''�|�K�|D��\hڼ�]@O�D5��'�׹6�yf�<_�nn�F��/F��}�tE��0����˪_Et��{0�$�G�B�Yˆ�7�F:}*��'!�xh�r�΀tQ��3��r�"�
`�j@:
��L+�,+0c���2�@�Q�y�h@����,�����e�%�a��7�����E<A-l2�1o�8�W���m�a�)&�_r캿ځ{rۡ�զ����B�칙���Ye8�@IM��*����b���d�ruvb�
�ܐ{rrL�K�����a�/LõE�T�������u�����N�y�Y+R�#�5�CX^��g��LO�i��Kd�@�_�DE�ќ ��t�M����c�4�a!|յ)q�F@��+e�R9����؞��Y8�}-l1��'%3�&ཎJ��+$Z����r4<d�l;�bQ�e��{��b��0�8Po�6U� �"�XCL�w[ޣ�Z���Ôa�P��gs�)C죐Z�h��[#�DZ�����X��m)	Smk�?h�{�S��Sknj�T�_�I9��/L�}�.V��J�}����f[�¢��j�_'C#�n��4��{8I��|�E*��t�ee0�>9�faJ�����ʳ(��,�#��AL�s�0��+r���#�%rO�E��`���̑�s�,��j�hYyD����;�ΎO����]�.�V�=�v�[iFԃ� ��u6?�\g�1s�E��0!q�=�Ӱ�;��;�ѝ�ҧ�8�x��%�s��ޠͬ���9��+r ���HQԲ�m<r[7�u�bu�*p�d�+��̈�x�@��e�ฆu"�[&��1��sy�{��������?������˹F��=kѹ �W��D�����uN2��u��%zx��gʣ�"ߜ^��t� 9x܁<v=lڂ��ə{�۞��:�1O�Ⰱ�WY���hsU5s�u��q�z݆8�t�]㔕6�#� :���ɡ�m@�	<��lGp�a����&BSf���FHD��`:�d��-"��� ���c�_�)\e�Z�_���Qq옗K(m��򁐂=)O;@�#y/��D����ݶ��s/�M솱;�M������z'cx�dj�B-	�Ͳΰ���j��ԓ�M�̵�T���m�u"�>=K��Z��P���~3�sh�� �qpB���^ٗ����r˹�q��S�����X���œ�%���\XL3���]U�ZǾ;��:��f�5Q�nTU u��ce9�뚺xŶ��S�P�Ȳ�#{��n�B��W>J�?���*�9��߹�|ϧԽ�n���q_�dۡ��h�*J�l��N���ɾ�z��6��a m�N���M�b=�kWt��`���=����1_�ǣX+�4ŧX�'�EK k�����A����1�)�G��A��ӿ����wj��+��d�`�rD�s���B=����)�`r�ON}ې��5���cY7�"1�é�Ui���%T檽��8*L";�Fp��-��Ԧ��pdš_���BWI�l���J_�x�9_8�g�L� �?�GN4��BAb,���|+>��_u8�]��+�Rҭ��N�)9IE�w̯���$�"Q�%��~�{[�c'�H�q@�{p/�q��e�0C�P5A��r�D^DC���/�+�S�hA�9Q�	�*�!��{ə�e��\����#�������j��6~3�[���.�=�k5M��cym��R�c���hly
�m��8�tI��NZ�4O�E�V��De�
#R�J$��+��B��xMc6d�NU�}���J�BA�l�(�T�G�����L�q�w�c�^3`l��f�@5��?΀i��K�e�������  ��;i3�q%hu�E� ��f{W�����Enb�X��y`�T@':0n���a�&2���Z�Z��#�s�l?.���_���w�ÛE��>"^ò����?���(^���01����ev�5�qb��� ��#_����."��^����zq6c=L���;�n�p�y�[iN�1d�	:$���� (k��l�N��קsuNW2	[���,��������0�Ѹ�@O�h���60O0�S�mq����08�����Ҏ�#����}��3p�'1��WӍ�,�Ĉc�s���� +��\(�e:k�b�)tJ7��ڇ��)a�`�5����a(nka<�Ke�j`&!�u�H���`8/<jI�6:ָ����%��|-�(=��¸H����WMӛ����5�Nh��;��V;����N�T������z52
�� Q�}�LE�ebd�XG��T4퐲��T|/�����2��V^5L�[�
 ��b� ~�r�����̧�o��y�"x�c�ǧ��1L-�Ab0,�����v��-�}X�Z3��sI�EI)�&m�J�����zp90� 
  /�'��?&oI���#A�(�đ,�aH2$��Hɗ�����������LWկ��W���g�{%9l�ٳ�WVW����:���wL���si��WgqFgq�>��F��U0^E�m�-���d�۴ˇ3Ʊ��jd��7�g&�m;��ե�#g���r���7�Nn�����p]��e��JD��\xcQ�20��n)r*�FGXj�.����cU��N{|%����՘��ߘ��j`Y�2&�;�7c�ӊ&���ӎ4�^�w^�v�^	�z�݌�����${�q��F��(Ll|!雹=���"�ء���q��1�ԓk�Y����q';�!�s cw�&'X�!���+�:�L �ߝ��6�u�pt�������	���V�p݋�1+�Cł጑T1��������<�1��x$�j6��l����}�^��,�"���/�������#�/i������%B��` ��=f'�v�֙�m�X䍄���_�J���)t�p6����T���ES�V K9���"VOH"�qN~ƛ�޾�����A#}$;���K��7��z��oN#��<F����� �M�m4�#���iL�j+\�����-_���v�ϕ�>���Ku�V���~�g�~X���
3B��_����%�%t�Ӝp�o���kPr�L�ڒ�Pw	{����?�R�5Bdc
���:cr��b�������{��;t�-��0�Z_�����7N�!�b��M�zJ�ة���Vx�M���}�Y��w.{�/�E�o�p�h� ��6�y��d;�-7B�����k�%��Vqe��ܷ�����j9��m$;(�_?'{e��5�0�DT�uT�G����Yܚ�4:��Y;p�p��el��V�_��{�]�(���g}Q����XWW֕ݸbEַ��{�r��t	����/�v^É�����{E�n��0k�cD�X�Ah��8u	����'Յ*Ɩs7�{�)�����If�����ug;�a�*4�:����W�q|�Y�h��[��F%����>¾
/��!�K�6�['���_�Y��s��p�����h]r-dD���I�����(p �_�uͷT<<��k�9]���0�����t݀l���[�X��T^Y(�� <��0L�c*l����v�cI̽��$((��RI���64�NG�X4F�Q߽]<����\RhT���~�M�f�#���s��U��8���*����kw(����!b�K��88�Ԧ�p3���.��}Yͅ�ŭ|-f#����H^=*�3�?�t�Q��н0�6�3�6f�u��fO� �P�<��̑U�ň��D�:�&S\��-^铞L���{�����������;I������J���aO.�29�G˫Po�qz�w��f��LV�Ֆu��s�^�%�7�*�& bk�@�>��
ᤴ{��f�J��:S$�S�1v���Ӥ�}�mz��_����St�4T}�����ơY�PR,�z2$7`Շm=���3ѦU4`l(���_z9O�F8N��^h�y(b��M��F瓄�񽼋/+09H������Q�` {���y�^S�/wd��&5���\�Rz?��\߶�ѯ���U;{����&��x"���2�v��T��]߯ג�Bˀ3Z�OJlL�9��a��=�)�EL�'oһ!�e6%^t�Tl���X���]��6��#�>�L��$�V *'LPO{�I�~�M���o�3�� �$EʩCy	*�}ih�J3Y��u�zˆR<T-�lAx����sY�u�U��:f���X(q}Z�oY�;��0u_j����"��̞7�rx�l�n�B�+���{{0�ֻ�'���Q���ޢe��֩�R��c:�j���߄>+Π~.F��(�� ��QK�Ӭ�(�Y�i������S�]D���>p	n�ҫ=��]��N^�6_y��GJ|͏:%F{D�a�NWL���%�+��N0j�W�n'48�φ�sS'�QR/�g��<ho�˜��E��({�j5��$36Km��{ �%tN/b�3���v�Bi�qm�a�QO(洽����#�Q��IU�H�4&e���@܇w�Kw_�������ɸ����бk;?�Yn"dn���cD�1�Β�f�x@HɅST�/��!D�ȏ-T���D�6�c���I�n�a�D�lp�.��&Z��@I�΋^AH&�k�R���<?CY��0�MYx���]���0���Ǧ�2;L�����<1�a��Y�"������]ȝ��n�#��&�)�e���~I<g�ػv� ��ʺO6'�,����h�6�S�r5���h#�E{F�y?����'��Bz1	��Ɏ_����WN:�6�G�+Y>(%@���ٮ��cNCe�7������o �5Z�ض�y4B2�m-w^��~_b #�0?I�io9��%5�He�b�����p;xK了ġds���v=�s�C\ז�Q^m���+ݴq&5z��}�����?����_�l���¶��w>�_ҙg������{�گH�A�۬�ͤ�s�s��ѽ{�+.�7픶ȣ�u^p%fZ�'o��tEm��9>�N�kQǗ�{���AU�M)��;f;6��|��9�K�u~<Lm̹�'9����L�Ǵ�8�^���D��H��Rx����ۂ��uF1�|L���L��?�����xyy)���l�U���]Q���&^���Zy�*�N6�cS:��%��|��1m�/tx4.��'��ޔ���q�81�C�u�� ������<���$�����E�,�9�@���|t5�.p.��t���ncl��Q����@���8��2<��WI���67�Y��Cl�p�p}pZ{�w���$� �����i����W��g�]��y'�5��~G�no�:p���L�������<�ܱ��>!��Ps���<��)��7[��6�tw�>��p�(v}K�02�T�-q��x7ѥ��Q�<~*��e,�x���Iy��lT$�M��J�ʝ���.��Z}oO<�nߣ��W��>�>�g?G/�������z��\�Y,<YQ�:�NI�O�t��	�x�� �i=,-��,?�~��H�	�M��cm�]����F�@� ]�'1��ƺ�I5&w'�H�Yh�^����>�Wr|4dݞڴ6��&b���,��핚����j�l����u{s�ؓ�C[���vN��ND`iǼ�*�Ә�^ D�U+e���	C���Q(������07�kmo�Yj���x\JW�� $��uN��t$f�b�����._�{W���6����X�F>���nF�S��4��j,������:���?5pV��*�K�Z������oћ������=�	ˮF�|o֫�j!�����;��c�ܞ�m�`.����^r5τн&�&��g�v��N���Z��qu��C����F_&���S�\�uٲF(.�����$�߳��m��q�t��USNw:%�H�(�qX�Z��GZ�O?��r�}���#�U��:���C�@D{��Z݄W�7��;qBnb�'^Gi��`�U�7�d^rMj ��L]z=r�:�zM�Ԟc�$~|Ք����R�3��Z�8����k�&����t�YN��v7t�NB���<�|�c�1}�́cV
�kԕ6Z���@�����
�~	។�Hy�'=&˥N� Z�P#�pUn�cq���D�hg��4t`��s��Yߛ�	�1�;U���}*]4����� �5�.���:f5~^#��Y���Ro�ʯ�g~�?��qC��$9����"��]�AE������D�8�Vk&c	o���~r��ȉ/:�8@QW�-Qb��工��*������g�d���xs����԰f����U����e����?9������+a�ɮ�}ݙ�C8����ޑz��Pb��3�*���ڈ�<a�@�֩<י���gm��y�~�z�o{X�Tøu]��:�	\��eT���p͆I�+�MO��#�0jx�P��`>��k ���غшex7�Ǣc�1Q��~�������41��l)�&�:�[9[��d�+u�����6�3i0���KϘ<:'K���[�pP��v;ڗ=M�|����ߠ��K�%�����$��
pkd?-�g�.z��V�	Ӝ��K�$S�{�5��t�`h{��'/������!�9��Sˈ����������Q�`�1W�q\l͑�-:|)f;���'{7��'����ڔEV��������W��QY<���nlK��Xi��b�׽��V=���q�������������7
��q���E�)= �C�fC�5v���n̕!�}������*-�����k���=׏E#
&V�����,F�4Q9�g�_B��m���:�s����
�z�#_3�\�CO*6樂b�����ZHT�ѪW}8^좕5H
�l��S�����,Bή���&A-�ɭ������dxp�	�F����|�]
�D�cLg��O9�^b�2ފ���;�!�\�w'j���͟VMo���jGcQ���pf�ԕ){�u>�!��;��b�=�����=��g�G�C�I��2��8�8`_q��ӥĩ]����h�(�3)@��u��<�'l6�A�^�؈���>���R[	F����q�H�k�K��%�Np�����W&�!��F@����,%eB�ؖq���NTl|⡜O-"�x+�ѡ���Gi�@��sb��}����?�M�S��	�}�C24�Ӽ:���Q�!K(�Ϊ�N�:��;�#����Y���i]٧��,Q)��w%��FkXl�1@�^ �Z��嬮0��xӳ�%��K��v��-�9��z�^.i ��ֻM ��Q[�pN!m���gk�D����ɐ��	C���Sc�l���ю>�'�w��sc�KI��=���� S7�($-:m㊶�qD?�9˛K���M,k�oBιHm���MM~w%�x�7�&h�)��FH��������H�'�I~Ee��pCᱭi38��� ����`���J�Ɓ���kveXU�'D�r��wk~���������[��F\�P�����](�H�7�~�Đ�m�ނ��ǣ$�M^|3�I�������t��(��L��\�UCq9[T�qʮ��>;���^��� �i�թ�S�n
�Y��O�x�Z��s��N��(��tj��ᠿq�?�P�+^PoGDk��׻�u� i��r��֔?+éz\Z1��X���[i�=���.�Z:���a�M�gq�@�7s�Gf�Ѱ�U��Q]������N�׫!��hB6��h���LF��_�I8h���xՊD��B[	l4�#bj�,D;u3���.i;�5�c���DVt����)xK	|�k���f���#Ne�M�VO>�e�r9~z>����{׽����B�~�ޤw~�w�S?����������qG�p��괡�j��R���L��l����v܀���)f[Q��m�m^?<�e�̬��d�i��d���b�zp�B[3����Ȳ�E���}ƫL�O�Τ1��t�W�	W����E���e���?���X;~��?j<xZ�k���Ƙ����бr}��K8���yW�R���C�:6��O:'�$������z'V�2ߤ)Y?EF��tU�tul����.��b9J|���5�f����ۺ����n�<%�<��t�D����bB�w��2�ɇ!6'|��.ኜh�"{�#z�Dޞ0��靻��3���W���?����-��U;��ݮ����A��E��f!D��~��Y�$Jз�@O�>��}�XP�����Bf�%Z��}��w���/%�o�q9`��վU~%�{/�`[J�n6g?tE!7�e�ڍ?;�� �Ez pr�Nz<@�w�C%Yie�L�n+��	^��R�ꞟ��L��k8��]@V�W4�2��f��nĊ<��ͤzN�s��!�3�g�<;]�����(�l�x�ž#bE�u����.;}���5Wz�1���6h8�c�oa,�i9e�M/5�Ap�d�� �_	�
ڗ��γW�L��m�����c�lsq`�\J��o�&�Is�x�jtO�s�VҼ&x��`}�����8�o����uĩ��ڌ���izm ~�b��HAR[��Ŭk ;���ϩ�U�·�=ɮ�.��z����SN,7�����@���|�����MyH��k�r5����.�	Z�(����I����v���h�8*���	s`
X�Q?ۥ2ʱ�����g����.��HL��� AI02}A����
��6�r�y����Si R��C�9<���X�dpw",g@���N�$`q�s[��%�	�gn�V�A��C����32C.�}����a.��#��D��)�����>50�/w68}N'Ŗ�}x��;_�2}��}���,ݞ��ɓ'tw��ʫ�՘�<+�gC�BݱN��3���K��R�6�=�Q(e"��b���?�9l.�٥��9Z�s�L�5��I���+v"���6��Q�Ek1f0�����2 x|�q)]�[ׇ�^X�B�M�D+H��-) ��}t�Nc)�`���$���Vn�}.f�0��l�p`��������Ki!���K6�V��h�yh:%-�+z�k�����A}Y�S�$]�o�!d`ZE��5�פ4X4�[���4�϶���F*��h�"Oi��D竍_;SP2�.�]���+Y��jgȿ������h�*���);ox9��|��xg&P۱ltg���6�3�ѴN��2{ԍE�f����C�iGǯ~����������|��k"�l����K�s2��k?�;��&?]lꝰ�)�0�W�y�����*�Ȳ���X=(7X-&�x0>�S����d�hid(�P��7���7O�;�!M��1F>^	h^�P�u��I�Z��jXa�N�9�q��3��lj�~D���}lz6`jd l�;[��b��:���H���G�8�����L��t�����Ҍm[ Q��/6�ٶ/xt'Q"��=�C��WqX=4fY��8�7p��Y[�q:=�Z桁�v�ş�5��t�O@��qM���Tq|���eU��	���s{|t!��{i]F6N��_����kZU�i�ܮǬ�a���
t^�@�,���v%�B7�������|���������N��ߜ^=�f�]6���>�Cm�*wԕ�n\��.��5	��x5�N�`�"�v��P3K`���-i����1�k��Ś֘�m�N��+x7��,���%g�hs|�[k^=��1@�q�Je]F���琽���@Ax�H����4L��eA����|�a��Xϔ�k��b8�@�㰍L��W4{xQK�RUWh�h��o��#�����s��TF�t<s�T�j��K�c�]�m��G��,˜y8!������ĩ��m��2}���J@�ÑC'h"?���W>��0�U��ȴNE§��웲��P�'��	Hp8ΰۡGZ����dމy���Z&A����t���r}�<���nN���o�;�������A���F�ì7�c�.j�{�i��l�ż���bc��k4C7���Q��4�1*�q��L2#j|ج<.�+���.��gS��I��:�bU-����J��<��Q�Fh�u�<Hr�}�Hi��'�z��*��\�|%���d>���=�z�����s�<����.�v��yGTIՇ�0D�WW��=���q_�O|�F�k�������_�sߪ�|s"�rƴ:���i͹@�f~;���p1��jl���<V����a��1wr�{�Wsl�YD�%���1�n?s~��8�s��yw�_�h����I#���ʫ��%p�x��wG�>d�{l��5G�7R9��� ���ʅ�㺆�PL/�H���wo��v5�F�ѵ}zx�D�ï�k�|�0)�fI�KZ�b��%5a9�8�"K$��=5 nc���O����\-�˽~{�+��1�����@_�����>�e�Q<���U��C��6�AM��Y������r{0��2�-�7J�
vQ������7:�M�(��x}7y�hOǆ�9����������j��0^�y[��*#��V���`�q"���Gu +�����n����G��?�����$}�S?I＼#���;��̳ 1BW#�m�4�?xr~#�7�s�|�������J鞾�&��UrX��U�$��s�>��nu.��?�(ݐRc�Q��+�!K���պ�9�ʈZ>���,Z~���VR����z\CN��)�#�x�d3�X�����1r���_�)�P���q�W����������4ac(e��!�Q���Ů�܍8ϖ#~���>��/��{3�%�����44\f9�>���u�h��g,���t:��չ��t�w���~d���A����.�r%�ښ��K&��I�����i�~�c��'u�$�Ьxt��R��v��7�]ϟ�W�ӳ����$�b-���G�m��c�ц5��fp�R.Vd�y��K�9��Us���:^����6�}�R���*\�7������4m/���RJ����ءGD3��H�t���u^1�}ry`_��w�N�i�&g����\��S���<�'��zٹd�d�7�p#�{���d|6l2�5��5�p�s�t��ڵ���5�x@�ӗX#��A��¸|Wh���}���e���n���%��+f}ͷ�~iK����yB�����u���cM��X�5����Ɍ"�;t�Iu���{ߦ/�_�D�>��g��w��2��P��9�xz�ff�2@���[\Y\"1�>�����A͵��� z3�%J�X��	���� d(����lM��R��v��A9�b�?��>�b[�C��s��Y�u�r��b��[���Ȉ�D>��F�um��Y�;ɻ��0��X��7v��g���_��r2~�ЈhQ�4}�sҲ|�^	8����9��7`44�\���2^�׋\��AJf�H:�^+}6K��fb����T��w���9��
�1�����ru��W��@/u,|-��vݼ&�g�:vDl�����f�)��g_�CG�"�
�œZ����2j�`WmTG��z��|������+��i��Wi<��͜�k[/�Ā}��}��b��l_%-'L;Ɲ��?f�Ǳ�ٟ��{�����FkZpM�ע�$��ߘ��� ��c�v���&�/Bd�ۮ�p��p[���!kZi#$z�5m��̻���|tB�����0��ԏy�U����F������Mӧa��gt�O�s]ϱ�ß�5t�~O�4�	���t_�f�O��xi�e/wmĚ��~q �+Gd~^G��cs#��S�sB����U�< o�~v}{��.㕽\��y�955ɭסS� Q1][�8X����%�{��Ѧ���?<)I=�� ��9��ð���h���K,���$w[@�e��8��Km}ՄE��\�.�����ՍHe�z���]jx��q�.�1��<���@��kM���e���l���2T��o2��������Ηi^齀p�;B`(R�	��!̧A���d�K�u2��@���%����a�.�oVL�=.�:����~M�休�s֠9�_!��xQ��T�>�a�
�'�ŗ�D�8�@��������~�����?�������N�l9�UDm}V�c�6���#���Sx�>�`���M6�x�j���Խ�)��Ȣn,�5�x9�Ϊ� �ҴP����#�ir�H56�����_��}������+z���HL~��OS�J1�����/�2(R�4���7.�-�x�i}��o��K	�l2:ߛ;⸣����6�a^wǘFhi)Wr�0v�ɔ�ad.��[W�\�4�+i�slޕ����Oԫ�	H������V19��񙾢
t�8tI~oАK��Y�q��xN�Bs>G��*�s�Ygjnx���]	b���i��?��B�㺿�TO#���͇;Z����O~����y�|O���+ƪ�Db����aS�Sc�Ӿ��|���D�kE�]�����z��|��3%�?�A�1������[�M����Je`ŉ�D�1��4�FY��?U���(s\j�cE�Τ��
�	zH߳.�����0��r�G��8�)� �6^�ySo���<-�/�^��zy�fxrλT��d�O�.��	I'��Ovk�Ɠ/�z^P.�=��x��&����:��O͆(7�z�b��{g��[p)Ŝ�a^�qIq`�����U���'���W��?�w������E������-��� �jё���cr�����m�f[:3�"S98�w��x-̮�И��y+���=��;���63��籆f����X��j�Z�;l�/6	���`�H�@�H��Ҙ��r���hx�Y_)C�}��9-%}	�!9�İ�ئt�#�ߴQ�����#��=�M^��I9�i������*d�f��B�e�ZA��K��l���)9����� 65q�G��P����a��UzOc�D���<��0�m� Fr^�+�b���Ѣ�������%Z�]���������LӔ.��:`/��)m�����j����r���w���/S��A������_-�q�
����~j��z_������%�a��?j
��D�y��\�a�P���|"�u����	"pQ�Vcm�_�I�.��C�q�(�=�0V<�k��m'�o]�'����L�}~?�Ғ���AĄ��[Bo�b��e�V#��FJ+vy�dW�q�(՚�OCsM&j#���4�w�Ҋ�ם8��,�3o���br��4��á�l��U�9�f��?��M�V��5.o tX}���!s~��5uh�f���Q���k0�	5+�^�Y!�1*=N.:��-��)ۗ�ۊ����ki�)4�c��ˎ*��%�)�y9AY0=6)�����1��1�iC�&���=��i���8�_�DA�6Sfx������E�/�(���X�ߔlvihP�2��O�����Vx�KEOp��鯾I�M�M�l�`wE1:ҟ��]hQ�l�I�B�`}GY�=�8mJ�W'��h���/UU	/W�!��K���qIx��4*����
^Ù6��2�];9��n�u:�����X��nu/n�@i�z#e�M;*w'���oЗ��h��_����?G���^�o���rXh�'�ݘ��Q�2�clJj�p"���č��y9qR�����=��LUW,�oQ�-1��X(@zV�b�;Ҹ��t6N��������3v���/�,�\bl�_��ĺ���5o=|��Ն���LB��P.k�o`�=���8�'�a���0R�0���!xK�0�;m`nڕE�t�4YӬ��JZ^�:e��,��Sb����(�C�'jO�6���6��8Q�I8�#�*m���+\��D���vd�[�'"�y�n`�l4�2�?��&�vJ'�jӗ����}���&����,�$\mjd��$t���\V= �J�;k��w�:eC7�XY~���J����yTl��Fsz'ϝ�<���Y��ՠy,tS_x�m����k��7���ߦ7�o��so�����G"uÇ�!��c�+�X��d�J|`$�/m�����p.��!*�l�
i3��Qg��T��O.��n���]8n2(h�Bޒ����]�Ҩ]������WD�SKXS%N��t�uynf�q��,)O��MSѠ3���1���3��#�.��O�r���̧�V�r2��j���&81���F^ˌ�[S�|�N�����JY�
W�j�|C.�4���z���RLB>��:;����>�����sk�~z������?�҅�/;	���/i��������oSk�	8��%@�g&�Z̳瓜�;�r�.}��>}�_�����J�ԏ�;7O�E��(��Ѣ�:�l���u�P��+����`?��N!�w�W&��_�[�C��e�{�8���r��}�u�+ �2��WRL��f�f۠7\)�TR�N+wתSu��v��?]�,���i�/KMw�ޖ�X@�+��Z&��jF����iq������O�`�ϓn��sF�F���d(�M`�s>�D�ۭcZ�V/�4���!�3�ڸ����QB.`��&{��S��g�u*��Z���D�l�W|�Za�q*ֿl{�X��b��U���NX��1��/�U�6�R�9sh/�Ӕ��8ma��v\[g}�4�!S�p1`�+�g��P� �Nj�Y����ӏs�"|!�b�z���C2�u{����뀨	,S&u���<����|C��zvsCoܾ����/��w~���{���J�Y�'�C6���5S2�dt>m�)�_A�)��t�܀<B��ᇋU_ʠ� �5��b}��:�=W�
lR5Guqr$r����uD�V/s�́E��������~������Ѳ3&�~����ꂳH���lG�-�:Ф��З9��k����r8�d[N�*U��:}�Hr+̐#E�.�]x��~-�m��Iۧ�b\��<�����Og��aO��ճ����Ej����^[�U�fD�����O:VMy�9�)�&2~��m�����H���#�]����I����F�Mp��q,�4��@^�<3Z���4du�A�4w���U�F���>W �V|�?�4�)(�}�6�v�a�&g �����Zfo ��G���Ԧ�\��,+~��)l���g�%�𑰹�B�̍�� �6#X쎭��)	�m&�ёf�#�~�^����谴�m0z2jtJ��t}X�dD��%�ׂ+����i��wA_�i���Tu�}J����������j.1
���zپz��,�+���*;�/,=�A��Ŷ�hkݝc�[�i�.	�k�Z��u�e��$4'[�D��ը���ܞ�^���˨~c�GF�s|�)%E���fEg����z�F-b@{z��n?�;��_�}�S���~�3�����oP���F��W
ԻE��M�Ka̳L�����l��RXp��w�� �_bv2��_m��jR;�݂<�}�ǃ���ˣn<X��I�yN���1��@��i��|����c�*6��J(w�������g�k��=�V����alp�sTRl$E�d��Lf/�h��܈�^�{
y��r c��}�����1�ܼ$f:�l#:QM@2y_�o	'�	��R��yJ�-�����c=Q��D�Nf����-��R� *r����㽔� X� �7���
;����w,z1��1ȃw�<W�JŴ!]�З�a3~�pб
:g���+8z��K�"q`��T���L�;��Z��r���T�m��Ά�DKVc##�ϕ��z���5‰���im����uLr�	�̄R,'�8���/G4���$�O0DY�Ws�a�8��w������t�����W�N/��E*o�������\�u�aJ=��QM�͑�	.�*�o5�i�8�ͬ��e�_Ο֛�#����m+6�l!�Ѡ�~$� �lOv�y^zms�m
y�Z���l��y�-�[:�A�.<�,#�|-�}���s����%~�'������) �l J�ME��` �k���YZM0є$7@�g/�w +P9�w�s�K��˓����`��6y�!�.���P�
�&#��1����?1K�h.@5:Y��xS3�>7y����3O#�PfT�Җ󟸲�Q2��n\y��F��w�6l�9�G�ar��K��K:N���74���(&�c�r�j�V���Y۶�
�bn��b������۝$��W}��/_{���w�=��'��/ғ��(ѳ''5b'}8���X���j{=���PP�T�i/<�ʍ��q7Pn�OL5�_��v���	����Ñp�K}�{)�n2FS��F<'}aq,+����5kG�8�g�w�(XI`Xo���\k����
%�C�_RA�%�Y��ųg��>��+'��$}T�K K�Jy�+6\�Q�@�@7(�c&�%�e��x�A�kɩ�R�X�O}2�u�}60=�B�ù���#
6x��(�lh2������8�pj#��_��Tv��g������ ��w��(���c��~�ڒ��i��Π��A���R�!�	s��h7���U���צ⟠�)�>R#^��/��Dr�dǉn�@�։D'���kq%���U�Gd��Y�i'�ID"�|.�q*�F'���H�XE��dJn���S]oRYuS�b���%-o�n��mz���R�����o|���_���L�N�x����I2�b�D2��I��遢{���x�i�8���]lN&��,�3���s�~t��	̀���e�ؕu���?hJ�
�����/ImD��&rG�3q��cJ�=���_������ĝ3��:��6�f��6&�#+�����}J�o��n_{ ����|Լ��^���4U��S��AT��[W5�W_]�d�@
��CWޱ�?�c�y��8cM�W��|z��ַᚫSPGs��^���P�Ch���!�I�r(FL���^�}U�{+�l���
3��7�
���k�#�r)��H��}�F�7f��ƶ��"(���޵�0�T�o/���PJ�6��b��愈,	mR�V�!^����lZm��ɥ�ݗ�XC(1m5'����*k��Wr�6:�v�Ԣ��5}�kH�-kO��n޸�Xi
 ��Ai�to������R<<Nɬ�'׭�wQ*��6	�:��W�ה�)k�D��|2���ai�F�9�|z�����#]��v�S��m�G����	}���MvU@u:�{s<)�բ��-���_����o�����|���O~�>����=N�>��t??��V���R�'���PÏ��5�)ɳ����֎M�i�X�ZF�����ӻ{��?���������;��!��O]�'�R��t� %��md�ƴ����T�d�hg}�.Z�vb��i��.}H��jl�"�c���$D8%�rƬ��X�Ń����l��ԪX����s(怵�GN+؜�;@�U 6���r�]�LU���(ĩ��u0���Z�R�.x'ǰH��:�iD�j�ώ�"f�x�cW7�kD��.�A�}W�?N56����B8V�˙�P����
�9ͨq�P�	�g�O��a�h����ղ�K|2� kĒڷeq>�N/�}�QS�|튆,$;���r7������2�Sf�[f�+h!���A����hr�w������ޛ�lHu��+F�AF(��Ū��0��#��"�P�}$���v�^-5�g��7'�5�n�����](rϜ;�J	��;���^�,f�������������{���&=��7��o���zzxI�]��Dr�����{���4ų���4�}��b�m�ߗ�L.�yĸ��GFѕ4u�:�N�Sr4�� z����<��-�p>M�nԐ�-Q�"��oK��T�7����x'xT���W=�~�Qm���ڸ+�}hS��� +$v)�l���a�~�oh?��9� ���^�|���۲EX4���|�{{��ھZ��Z�ѻGPs���E>á�[-F�Y_+�`x2o^P��\��](���r�S�z�uI_�_c�W�ץ�\4��ʊ;_1ZZ�!����JjKො���ԙ�ꍜ��O!���|T@�$~ݘE+��gz�?};�����>�=���IO�������'~��}�c'��#D7Oh��tWՍ���J�C���omʱk��ⲄbCܧ��#!lj�_�F�`��8������:ޟp��Q"!�ꎯ��b��2�ƻb��&��>ʝ�ɸ���#�Ţ+Mn�qY�,��Ĉ��F��{��ᄬ��Xz	l��O��+~e6�!�Ah�OKӯㄨ�D����d�?��+��":F��'�W�,�*ac�J[�_�N��"���\�����5���p
_�'��q/�Ç�ۓ���q[�L�.��ٰ>y��l�6�E0a�u}�)9�h쒜������'�wu�w���c}o�9���>�L���s��m�4�Nx�3�?��\S\H�~w�>NE�{D�*p`qޚ���4Y�U��N��#J�f:Z��k��Rݷꪪ���������#���(:4�~s�4����!WL�N�z�?>;�0�i�?NOn>tz��<�6f�h�䛐6~ݘ?��#j�$��ȯ�]���^W���j_�s���h�����o�M�|�+tx�4�x�>�?FϿ�MzrGT��EBn�ȟd�co����%ٔ�z���[��~��w���pY�e����سa�F�_�K�;�/���>rǶ�����s°�g���C4�o��@)
��v9�^vWX���W8�r�?��q`������}���Ñ�O���>Z\��h�A�3]4Y�"��,�a��vĊ�*�6b^�؟�/Y��i����V�Che�e��ޓk`�k���=`���odu��?��iُ����}�3Tհ:&��,R�RZ�U˛2:���P����94�BdE��\n��u���d])��y�ʵ���wG
>�����v�qZ	�Ղ�e(��g�ʠ��m�n�-���
*�h��V�ܨ~���_�p�6e��`�6���hp�Ӗ7ɘ6&+C����v��������GZ��=T��Ɯ��!�z΂Ʈ�sm{�sޮu����=�\��fp�<ú/��U���)�nB��.�HU����x�d ��n+S�a�$���8��ky�&8�]N׭���ؠ�0 ��5��afր5�gz6,��7P΍�'�)+���Eoj׺K~q�#E�`�;���T��η��w�I���ߦ���i5��Ȇ`���Sj��S�MKRZ����oZy��@Ɋ�����w7���Kzz���s�>���ч~��zn�ᢆ�+3�G�Hc�M(r	�S�U�;b��X꽯'�,\0�,���:b(�S]��/�-�le�`��L�)����ER�K��B$�a�������j��D��,����D=z�����޽�n��a����ZYi��I��8�&	�:O7���m!�[�'n�C�_�7"��k��9���x=�V�>Ў󽢎7�X�~u����r�Lh�yv��^�Ǎ�/i��_&�]�Dr}X1'���� �Ō����@\������?�����y+Y�N�bHN�����ݯFpQ���;aHrX��f��z��bŋ��"���Lv�Ie�݁<���tXOg�S������lMvb�B�Y�Sj�d��5���{�F�C�QH���������>��紇Ë��aR>��g�9����jF�%˛� ��H!x�9	�f��u�瞖�{���ON-�P}��_�;:2ŝ֌�ɜ��Jf�M(���Ʀ��_�H�<���}`�;6���%9ܕ	�~T];�"��u},��}�����2ogk���58��p=�D�1�Q��̧vg������>��s.�Q%�qH��#}�X�-��N�����r�ɕ�ѹ� \����G�c��|+�w�3Pm�����rJ�VIϒ�j�fӯ��[y6�	e�����mO�Ur��d��y�2�����逡S�jNW�c���[�����,#�1�{O�MQǾ���#�|#2�:��ҋo>�����T~s�eW�P���^�{��h Mϖv%����v�$;�)�y��p���������=���>N���>��O�O�کt8�N���q�A��k�l�8B����e<'ӯ�����E�h���V��4�)�߈���#� ���d�@�U`��G�ۈ,�h��0�"R`&�ɛ;��q'����rĆg:�@��S7�E���!�+�I�I5v͵J�Hn��]�"�&5Gjw.��6�������;�*SI�D��͠�'n8����&�`~��z\��A�Ys�K���S�?���2e1}�6��ښ��o;�t$�ׄ��HC��-F�B�	3%�ނ��	�v8�~�IAJ>��2���b��19f��C�=}ߩ������j_��{��̆Ɍ�g�G�5���':J87�nR��C��Y�O:ͷ��'�:_�ίP��[��CѫeV�;"�M�;JW��
*��Vm�/�k��z�9Tu����Ozϳz0gw����!=��y�t{�˞�&_��eT���bz�ce���C�A��lI,p��xe;K釥���M]��-���r�	��$�KI���آ�i.K��<P��%���c�	��ǳѕ-n1��#�?�ѥ~*�H� W$,����5�H8��~Odk�=�g�u��R�H/yOK됇?����k����z�����������o�h�w�{��SFL���v�K�Q;��3�^}v��o� ^��WY�t��9p(LɅ�>��+�M���\(�t��6��rB��a}ח3���23�i� k��vdAF%m�D�k-e�ki�`W�6/ڕb��t�����K(��ͨ��������[�:��̺��Z9�$�`��a�� �0���+b���������sF��;G���L�Hi�T��ЮR#�;͕7�\��Y��
No�c���f������2^�ҵ����k I1�p0�� ����.��d gP��Sx��|�)����fj=�/�}-�f+��>�KP��H�M�z�J�y>J$�rR�w�F:��Q���ʭ�sĩ��1�����ڡ��3�����ϕ'3>ˁ��'��}�=;������G���7�ӟ�����:���Iu��pj�;w���O�s}�f5n��.bL�[{��L����S��G��b����t\��POm�q|��u�Tb�(��3B>���ʆ����v;
Я�1�;�� l�����u5$���z��p���ѓ�'"���ՙcWC�N���Neđc'y�7{�vBh!R��ϧ��r@��`y�~��cN�@S�&��z��{9k�l�c%��� ���F��9اc��.��W��@�⡃ɇ"��X���K�!�(�%�D]���á�9jH��e�w�G3�Wz<F���jrJ�cǧ�
���1�7��Uz��N��{������HwNw�h�:U'�M��7q��f�,������r*���8�c�ĳ�m-�~�M�4�l���yC�rK_��/��?�O����_?�U��uz�:�xAm�GK��e�5�b`�)[�bК1�S�)�Y��X#���3�e����p/�E��H����ʾIs����d߶�
�wn�J�23y�/?�YB���b$ۡ+m�X4{пٖ�������>w�L�/"֑���p#���/Wu��p�Sۖm�m��5*_����i��lahN<9���{���u_��K��0k0B}-m�>(u�Rk������??�ucG����'��b�!__��B�q��8tb<���d_�e�ą�A�"�]��[�o�`���W�s��M��u�������a�ye�?@��l�f�}��u��.�7h���n�8�����mճFM�9��X7H�zu@u��U){��to��/U$�����Md��a�Cv�#��D�X��~u �r���$���#�0��_�����G�!}���=��Z���A�۴��+z�ˢ!�<Q!��i��b�����"ԡ��8�׏��N��O0�T�Mzy~P)��ev�8�^�!OՉ׏�:#�E[��E,i�>xPm�͎=���'��s����n��d;�u�;ڟp�8W�pe�m��wz�(C֫�jY���鱗��������sx� ���D�	a��s��ƚ��Aj��b#�������*��<�/����������-�gߋ�ć%� ET���'|!4���R�9C��9�t�+������:�W���AF��nq<��S+����3�y�FǙ�ӿ~�	4�S���	�����f8����a��6ݦ|��˘"�7��&U��UOz'�E�^�5|j�5�;�q,j�]�8�3�\�ˑO�Y�����������?�Z=�B�ݍ\�+�d�ÒE� �-�#��>��T(#� !����uj��#{�A���?s �cV������J`sp��h c]�6�q:K[o>�-Ǐ!Fq�y�W�3�sy.���g��K�*g�Ҡ��LXpd�n��pƪ��o�g������(u$5r@m���_��FZ�~�>5���F)��ظ���_H)��Zš����~�|����K����|�˗�ЃiZ���[0����IP�8�ك�9LK�@5&���׌��Mq�,��ך���,PئW���*L�ߋs�7�����)�
��񝺑p�ܔ�B.��,0�\�%�[^�71����u����}z]�<�a���$�K�kV�v�ɗ�ٻ3����F�M�!����(�Z�S������s�񛷭3�n�wd�~vӿ`�G�^�nM�j9-w�a#��>+�p���@Z��a8����<�D oTW�NكUD��L���s����o��q����� @VG�R���drJ[F��=7�p�a�g�1g�c�~oG��I�a�n�m�Iԝ9hȖ�&�`o�8�z��^sr���Հ%�Ұ�	r=9s��E2����K���mN�� ���ղ,{��B������g�S�s������>���wj��j��Q0���VY	0^�����3AFᑫ�`W8�I2r����ɜ�ĉ艹?ەbb�>k'�A�5J]�J�,����t�ƌ4I6���Lf\�Q��:2�r�:gTÑ��L��n���Ll�K���8Mz���Yʍ�Z�2??=�k��#N/���'�e��f��'u�5�3N���5p2M�&\s�Ǉ��p1�aěLz2	�Gf8B[��&OP�J~Y���8�����J����:Y���&w��p<��	��aQ�����LG�5XŁg�2�';��(��
�7��P{O���aYV�,!}�-�cX�{��X7>�ʶZһG�ZK�X�k�P�����q�d��5�v�L���/���o��8�ѳO|����⿢w�
��/�"�}uR����N
�pх��#l}�m��]:]Y��黖����Y�i�c��u)�Z����<g*jc�r5��y�Ȑ��s�����/$SڼZe�/�����,c�2Ʉ�}���Á�_׮��x��~z�~���/E�*㝭08�@sV7SȽ�?�p
ڏ��aF���0�����s�-�z�g͌��ri�~E�Q�sy�ҫ�<׽����r��|�e���:�Y���G�y���n3s�+ٌ��q_K���Q�_����66��&�[�����1�Y�&�^M��F�Vj��{���%�M��W�o�I��}rL�7ZW%x]vp\�Wv��n�����=��=�V�2ż��/���<Ug��"��S8���,�\�ۛ�M'g�4�I�wý/��Q�����b��nR���T������M��������{N/3����w�M�t��2���6���*�v�7��������d)���Ʃ��d�ٞ�0�ƨA�/�� �L�3)MN� ����dku@�ٮ��G��C�d�|�O&�$�u�m�a7� @���A�:.u�x�Ł_;;��p�Oy�t��Ϫ(�R�WC�h�p� �=�(=1V���XWVޔ`�'��`:������U5؅�&YP��m�_0�f�KN1�&�z���H�'�`�;�7��J��w��dNo}�mD�[�NR��0p�'�G�Z�oz�|�c�+�qJȒ��~�٤#�M��W�n�q�?��w���J�!�$�z�%�2q��RpݦpBmy��,U��N���^u��Q�k��ߠ�<����o�Ϫ��߄�q e^k�U+����R�I���#�]��G
,I���.��XԖZ� � �]�'*�U/��H�}p��s�Kￎ��4��l�s����6��:�����p���m�����^i���˫YU�ɲn��������I+]���>�yzʀ�]&��2��}}�K�<��w^�מK��d�}�F�/�o��\�S�%�䌏�c�6Gkt�^ߧOmM��am���MJ���}Z�Y����qm
Z���m\�;�:�}���b���}�h��Ӓ�0�n�Ny0����p읻{�O�~>$�Q:Lq(�Gq�'��i��jh�9��>�y~<7���F����SC�eK�wik���x!����PF<�4�d�n$C��$��ܖ��\3>Wm������0�h����5-og&�y���K�sU`�X8U�ŁC���81�~���	��)����)Pm�.��l嶥�Ӵf����<|w����v![��h'[|x,ȷ�\���s�I�=��=n~�x���s���!�tcTj�,#�y2��Dm����(�mf��զSt��oS���v@g�N�4��T���k�TX��&�w�ڿK?���Ћ��ұ����iwj�#z��#���Wx��֖�V}�m�h?�F��!��I2��q���,Ʒ[�l!zi�v�ܼI�ӏs�Ny�#SJ1�l��ꌡ1iwI�Bfq=��vO��rJm�ũ�I�z*=�	F�Ifq���������qBIY����	wr�X?5ʼ���\O��8��+�0�b�ϛ!�J��N�J���P8\4s�l�T���SC��@�����p�P��zU�D�a���w�P�r�y�Ǣ��6�v�^�q�+	gx� e�xi��(�?R5�v}��A�!�Hg�Y1��:r��]W�ᤃ�;�d���<T��P����Pƻz������ ��������G�B����'z�Qhv�M|,d!תǙ��&� �^Oh>M��e>�m؀�7��j���.1n��4�,����������9��'��o&688�Ǩ��W�m{_G.;l���Z��j槽���4�w��RkǛ[�1=���3Mi�c�Y�y+m���Ej�Eԓ��|�-sz��J�ǖ��Z�/pt>�e��2>_��k߹4ҷ^g�e���{�ƬǪ�}�����J�G�<�>��EX��V�a/� ���C�h >��)�;��+��;�W��f������bM^�6����)F3�;���6v|��>��Z#.���2 ����yM�\r\�����C֧Gr&ǳR�����o4�O�����2 u��mW�_V���=�}C��O7#Z&�C����S9ӟ�����g�/^���^#���k��B�F����2��9�Mv&���gLqE&���\4"�IqI�P�[�nJ�����GEDTp�ʉ��C��Pw��Oq���
Jw��A��q�c��2�K.�9kԈ5:����o)�Pk �i�D�H��5��X��#1��ƾ���*Y�g�UЎF��Ϸ�b��"��`�G����+��v�i#ME_����8^L2ƢȈ�^�=iTB�1��ur�W��;u�$��)�
E�p��v��p���εZ�6��V6Ri�Q��"s���ʪ8p�BƦ�hi@��M80AJ���J;�W�D�n:��s��r���Y�W�o��͓��O|���/��ʯ�:}��,NMs��r2�fʼ��!<%\	����d��� D砢kv��U~�|�j�v9�<��} �{])���	�j� �?�W�[X�k�1���-�v�.|W:ER?��QN��%����6o�-eإGc�eO�Whȟx�F R�=�M��&;�ql���������|���O��O��o+be����� &��en�೼stY�i��@>�vD��S�t�����9����ҳGc�4jC��{��l����6u{�����߈�嶬0�c���2VJk�QY"X޷��ԯQ��u��+,��%��ɮ��@jo�O��:.JsI�t�x\�"���ڸ�K��;v�x'���Lj?)���zd������������L������*	��G{�h\hÀ�Ӿ&�׾ �}��[�2����g:[�����<[�י�u�xh9�
���%ӏGλ�s�`�n;�������aOU�B�Mk�b����h9�E����+�-����xZ�����b�_ֵ(tg���{��4R���V�����g�iUw�#����fse�J�R�h^?�ES���py��q�|�j�?��h�vݩ�f��d"sV�3��z�d������~��{yw����R�LJ�j������$`��F�ma+1�P� ��֕Q�\�4��W`�csBd�l~�S�">�y�0�i���"�W<t�_J:IU4|�r���ac2�H�i��ދ������jk�Z�>إ��Sq���i!'���3}` Y�i����	��E�flIM�.��yļ�<�J"E�W7c���ҹƽ�6��{�~pD)�i25�L[\��r������Y~�cބN,b�������9֌��D�o��k�z�S����E�x�mQ�������2k�c��O_[E�px��N�2i��Y�)�pL~�ʎ�������~�O}����!z�;��;Ω�� ��Sv}��3��8ŪIo�?�g� �y�jJ�w�A��~j�1�M��/J��_Є�|C�Ե��<���g����%�e��#�پ}5��w���{��aI|}/A;M*�����8��x�+����\h5��j<w+����]r�@���yF�^k4��~�k���w��]��h��z/>���+T�>m�hj�����+H�21�9,5X	�z�@d��H�c�˸`�G���\���W��K�\/ی'�l��QIV���~�����?U���S�9[��T����Y��I�l3Yr&6�r-��֍��o^�<�U��W�8l�������=���B��9���8 ����Ix�6v�fF�8���_��́��
��'>F�e�c��5��8#�/���z.1jXw� A��q�ȷ��ή� Ҥ�N���n&�N�oPk�)��c��[u�V������Dٛ�Q��D۔U�_���0�B��1�	p��畔O�6��\�� ���E�b�hD�i��7�o��@����0��["'�!��`����?�S�5A�W�ޔ1K��ٕ�"�9�pДs�9E�κk����8R����!�qѭ��j�mQP|u�G#���9$X�1��a��f���5�A��Oe���\�3���������Su�9�9���?E����ů�i"v�C+�E�ԡ`u��cK���	���gY}�~�<[�%ϟAPl>.X��-��N�_�6L����U��L�0�Vދ����sc0��n�n�n�uLN��C2���4*7{��)����J��j���ѫgꏂ(����~�I7g�U��,���lc,��w�W����6�Ь�(�u�?ڃ��/�k���1��F��N��V{�H�la���3ԝ�V��1#B��xn�{chz��[ p �brǺ ?g����5	��2��oF��H��j$�y!���?Ή7�^gkT����Br�����+o	��a'��4�N��WF^��� �(����q{\�dD] �H�e�)�/sT�C�g�O~��Y�������p�Dk�u�x���a����N=f�D�������Ƹ5��f�6|�)���+�ϸ��R�;Ej�j��{���@ƹ%ԝi��CY	
���\5�8�7�kHs+öhƆ~-�$U��������S��<�R�]�f�l �/�Q�z*PY-�e_�C:%x~ɋ����	צ@^؁�	���M�"# +�[c"Qzc�~�x�^�n��F�c:b�NEl�2�OJޚҤ�w���(*m����ǌP��|�fZ���i)\NH�/ۭ�z���#3��?2E�%m�0h����}�w���+Jˈ�q���3�S������h�q��86ޑ`�C_m�m�EZ�W��ւ���^�`'?�[��>M]��~���Ez�R'�ʙ��L��]�0<:}/(H��>NE�2�_Z�*̖:�qi�����YN`ֻ�g	/��� b}F���~��{B/O�wDr)G#�HXn'���-����7�iEf���b����Y���6M�b�ԾɱO0oM>�xk��:w�%����a�G�����������Ù�%o��f�Fooo��j�ͷ���P�DO�Yփ�e�8��_7����q҇Ӗ��#�k�y��L'�{���J�anN�����#����nH�k�C����q���y^%�zN�m�`	��UXϲ��\�lkݲK��&z�f ��?g��uJ ���lk����#���%��)d:wή�S|
�sdeڟ���ݭb!���'�A�KC�|�1��/�I{�Zb5�B�cP���nw�y�|cת�7������9ͅ���i���X�*đz���p�*S�{�`�o��N���ݻl}�/v�B��R��i�q\���~: آ��d�<!�����I����8{�E� ��W8�LQ���Nc�K?���W����y|����|��i�+��ຖ�b�q��dgp}P���-p���$���Ri�D��Э������K�d�}�!�q,�DK	�D�c����$\_�1O!�~�bK,�)�#h�ȵ�D�&wPh7�1�ڦ��K��$����8���n��Fv�Y�egמ��S}�;���魰��P�dm�+�)�^�Jn�چƩ_i����CL6:��;t��:�����H9!���u���o(n�q����������������7���ДD�ޏ�[�*X�E���B���={7#լ[Y�_���p�q~P�w�Θ�D����O|����?q�U�M�Jf��Z�y�8j���A�M�������>�>�4�qT����K�s�����dQ�|"ى���?؈r�����d�*>�!�3��5[�Aj�,�^��F�	��L��2�k�H�2������\��m޳�s�-%�7�\ه,�e���ys+�#(%+�R� T����Z��A�2��]� ���j�X�g�ӷ����F^�M�ɰG�ڻ$,�Tg%^1m�s��RUvB�<_'^8�5�M�9ى��?/���2���>���z���p%sz ��W���[#�@�lt���p�L��-m���}6�J�JIs���s]�J�A߸�m�"i��ǆ����s(�I�V�X
�+�'���	��O�uC�h���>��_��c5UL��^�!F�z����q�gc��w\���zUK�L��?kXW�i�p����"�SaV`���}��[!7zm��1B�q�(�8� 1�A68�j�˘�R�0��k�f��N��4�]9��B�S0�);g�)+m+N=�$��Y����!��T^xo-oVN1c��1J�:GKb9��h��s����h?�dm�K�]��|B�nF�`�~IXz���l��u�ذ�_S�&�&�C���$��Tg�bs:��j�h�$�	)ɉ����x�Ta�0�H
%+�*f��=Z��H^i^����S�	e8�,vW9�2jN�P���p����;�󍆲4�Fߩ�j�=����|����P�6G!1�9�X�m�:�5�15<ӹv	�S�wF�im��$�8�}G�#���L��ӫ�|�L�W�m����E#��X><�g-@S���q>��R+���n	Hq����8���˗~���������V���z�Ybc`<[�{���%:�a�U�����y��&��
�2���r��逸��>��V��A��^JW�4��&���!Gy,=y\IX6�K:��5j�3���Ln���p0�̙\��,��������,���hxkЇ�=�}4��vP��p��<��AZ��q�?��z�g�ߋG�o}�-��U��K���ɳS?N:��^��(;��p������\�U�;v�&O�$F9��nT��x�^;O僫s���|���<��v n������SQ(�q����D���mp�e�V����M���c��a�r@`��'�ݹ����e�������z�l�ׅ.,���+��Ь1�})� t��6Y�Gg���%t&���u�)���;����AU1%Z���IipL�N�ouz�TP�Z��[�ZE�h'�������1�e|����	��-�O��:=�V�NAl��å��sg6������iLu�`[п+ߨפԱ���l$��2oj��6_�җ���<ݟ��ʏ��c�+�瑵s�=1%��p���V٠jD�e��M�N���n�#�6�674��-ٕ-��WR9��~S�֐7��Z]����ԝ��)��D-]�f>�X����\��M	rU��ƥ�Xt�x����n���ۮ����?�?N���}����b�k�G�.��/Hz��p�b�u��>�5�c[�q�F#2��v��д�^�gоT�v�-�j##~����xի�'�:�#�~.�:K⤝�����a�z�� �Vo�ӥ�G��H�����rS%�c~��-I�J����L��--��:ζ�!��д�W�a��.W�G1�L[}�0F�C��c@��b�l�>��	��t_OQȉ���wK�Qsc*����m8ӧ~�_�ߜ^c��^�����5e��Z~lj���{����I!�J�|�� Ӛ~��#��N�A�?eC��e�0JKf��CR���&���K�¯0|�jAe�;����ᯯă}è�ў�\���<A�uyh'�6���3R�(�{����>ה��mPn�j}����-k����kO��qQ��?���>��?D?���}��TN`�9��݂U	3;N݌�)Nc�<K�&��D}!���轵%<���k~��ZO��W����xT�w1\�r]�pc#�v@���{�3V�	1(���@B3/&�nd��4�El�w'� 0W�椿���?ѐ���|�<�yn�Pʞ��z]��bw��\��Zyfw2W��b��T�������Ptl�t�n�q�]�7�;@ƆNI���/�61�_,�%��da�m>t��G��(�"'��~���8Z{��Q������#ˢ�+4x���zB^"^XG��j��.�X����� ǣ��Y�r��]�i��z)l�ބϸ�	B1�N��02�1ݝ(,��dkRiR���@�u�k�I��s<�u����G������h��ը='Z�;������]�o2�':��o|��Oe�;ߡ����=z��K�{�?����Ix;�>wƘ8��r#���yaJ%���7���\���,�+������7�7.3!q썄�G�Eɕ���q�t��vZK���/5��8j,��M���6�9�Ô���^�xO�f�g�@�QYD4e�m"P�o8Sd�8)I�%p�8mf��#���#�>�9}��G:g�k�
��اo�g~2(��sN�����wU����g
S�>�uX �<�3Z��Uޭ�D1Zֆ��^r��z�|��O��+���%��rt��:��ëR�!�;����-�<OKC�]����;��p�ț�P��� -]h6�Ǟ�~f�c��:����E��{�W���{נے�0l���|߽W3wf$���!�z�4A& )
�a��b�S)�)�*(�r��l
0��Ꮛ���&�\���m$�y���4#�4#�F�����q��^��ݽ�>���̐���9g�~��^�^�z5��{ə e������ͯ�kx�3��=�yp���wr[Z��v4��ytb�x-�]OQ%x�@u�����d(���r���y�E�L����(�ѵ�I��7�abX�$o�l�~'�m'���Tzp4���Ȳ���#���l�z T���,���u �9@�Iҍ�X��_9>��$��
��H�h�h����ɕ��uYv*���0;���`�20Bȵ��0B��߲�1u�+�p���Q�t���?��r���u�co�=KݝD��q'�����R`�n������߶�g��[F���<f����l�;�����M���Pw���E�8?OW�n��ހ�S��Ǆ@��vK������f[ g�҅ƞ]��n�Ƙ������&�DpI�rd]m���"�]��c�����;���8�Y9� k��i�w�ve�wul�wcwz���m'||t׮>#����=o~�[��>�!����*Ёr8阰	��,߃�^~s)4���9Fjv±�~~���cY`��KKSr��������|�_ո&V��s���!�M��T���,l���,�2e�n�SJ��~��d�ڳ?BV�e�|�m�QZ6�n�$ڟl`�<�P��<E�{�s��٠H��N���7-ǝQW+���8�"�|OQ�6m�����,*_����eX�JuY��#^ͳ������'�[7o#�u.�o�����c�Ā��ҷ~��>C�S�BFǄ��]��G��B�,[Q13o�Ҭ"�@̮���u�2-՗�3�>�C�)����T�����Ŭ|u��a���eQ�e�}8@�,	��x ���OB���H�1��W株x{�ݢ`݂�Jv/g;8��:`�0܂><�ya@ۃ�=?O6wy%C��(�|� `�9W��1��l�7�7v��wJF�lI�n�#�IIܲҊ$9!���lP�]��mF3�^eqOȧJ	�Y�R0��� �8L�0��
���l�e&ۜ+�1<S�1��ꕁ��&��0�I�&���w{'t�]z��A����a
�h#A�k�S6�QB˹�jd��i*o�_�|0�	 n��KE�IZƣ+1�g�B��	O�����걈�ob���h)�`���p&̯G���䲁�`����������N�r�
��z�������]��Yr��	-��햼�ш��\�.���y=	;p�Iz;xa=�C��;D���;��`�nsh�b����K�1��_���	�L�f�A�ag��3��`蜱{v���h�Eb<�Y0��%�J�}�b+���Ցơ��Nc�8��v����Dq��$�G����B��Odd�~m�!	y�R�d�x���:�D�f�q o��:o�a`�Ea"�1�&y�ȨM�0�n����6R�Z�>2"�3��׌�b��s����N1(dൡy�yi�l+	�7JϢ//3n����Q2� 4DN�"��f�'y;r�9;��_���oNwr�9C��s��n�N(3���z%Ql���MȦ�4L����*��6��"�je��J�Q�ט:�F�P�%q{&�'���A��q]�x����4�B���������mxy,3U;b�����I.�z9_��d�R��F�t��p�����!!�Z��G����=���q��_N0�n-r����ח�O��;���=o ���)���R���Qۄ�2t(Ap�R�f7|�x;�3iO�ic��]�\F���z��Z�Fk�P6�!p�a;.��Q��l[w���4DƱ�?�%̀e�M^"�����?����9�6Z�b�Dh�6����5:W�������������*�הQ>��7�;r*����Mx�o�����kW᮫W�����n]��.�lУ�zڜ�t�~��t�9u$?�*}�m*8>J B/���B�UD��N�<"щND���N����JB��
Ϸ%�F�z����z�8��('�����A��(+�wc/Ӷ^�Q�gc��#��i�ޗ��Q���ŬK��n
��8}���W{�\,�R~�+
#�E� �HOu��A���M���r(��[u%�e`T�HG�����Y� r���L��S0�H��g��ݷ�(�IŜ���R�0 GZ2�s�����;Շ�#KD��:I.鯗3��uU$�#Y��ZY����%��`��i�.��m�����I�|JG�	w|u{�cw|tNNϰ��(y���?��78G/���`��M��6����Px=�0v x�Ĳr�U-�4YR��8�]����#e�ٚ��M� ��r�]��QK�����A`��6�1�^y?�˓�_K�d;Y��ߥ�$t�nڦ5��φ�J��^x$�K��D��^OG\�58� ��2EbQb<��Bq�6>5)��d"�8�e��9g�"��A��w������~��ț{��h��C�!�}�\��n�QK����&-qy|�֊V9�e�jr��C�ے�ŽhLV���z[O�K�/�vY���v*���Ѭ?��
�ȋ���м���^�G��,��#p�ܴ�Rk����;[�JC��FO��V�w�e��<K��-��r=-�7A���	�m���V��O6��\�4�Ph�Aݵ���bsۚ�]���K~�+ocQR���k,&��P(�F��I�>�	�=�0<�/��ۉ��$�l�%��3o���D�����uFf�e�UMb���גl��֕1�XݞDS���7b�/N��|����2T�IQosߖ	kY^n�2��Zm�b����;�@L�'�|�5�@W����G>�Ǥ�k�Ȥ�]M�w��I)-��͹Q��ډ�陚��8�|�fs,��8d�8U���U��u�Y�A���q���F?�@�ڏ�2y���>���/D Ri��{�t4{N������S`t7�7����c�������~�Wó�aH�D�����o}<��G�j��紱/d�"���G�xO�I�{���� �x��SEQa"CW4Z.�Qq����#�OE��N��� �n5D�1�lq8 %Qu	-K�"���X�����D�)��*���G�:�9,��b��K'{�GkB���cϧڌ&r�Ռ6��3QvrG�0R8�%��"s���廲.o���O�Մqq��(:�@A?N���О�`6)��_��32n��q��b2�b�y4�n��/b��H�0��P�%�ᆎ����J(QC�>��$~g���
��OyڼyZ'[�/�BCxç����d˞O��"�0�%O�� ������~��S_�b���{qC$m ~��?�_���|�{�Z:1�^_�SsQp��8哚^^yǺ��T*��K�+�
]���i���~#2�c�ci�"/M���:����k���Z�*�I�ji��^��Z��V��Y+����L弳�]�&�5�^`�/W�G?��k8%��״�V=|��k������ɑ��xs.�I`��
*3�I;�:%�mǺ���cu�J��5p����x�MT����9��g�ܺ&r�e�1<�ڲ<℈n��/�3}CH��,��n���'��Ԯ�'���e�5�(3����xqaݯ�ߨ<@L���E4��sZ�<��Gd�=�G7O�a)3�n|�"��Ei �R!��;Ƥ�=����价_��pS�,=�u����������-ǎ}����ɰ+���D�byCj��?��f@g��'��S>�~�ʯ�2x��/�h{�I�6Y7�g�������<��M�����Q�ڒ�	&����
t�k����+h �s�A@�G���3�ɘ~��/ā�#��tM%��E[b���~A
��[��h���\�6$B����9џ�z�Q<$�[��;�]/�+E�`[L*��0X��y����_��L�ֲ�ʸU�;���ƨuK�Yty��
�{�c�9D��99X�i��Pc��'�f̢���D�#ف�u{�M8:��*�ⰾ8
!E��H;�{sv��iɉ#Z{�ɴ�#�s�����Ftc������.E,�:>�N!����o$J���8g��e�
�2�¯�^p�#2��{:t�.8�n��y|�W��%/AG���ܺ}~����W��>�(�H����1P$��ց�'#mQqx_�8�̖��gvs4����[�������G���|t���P����E��]E�;,UT�ߗ�J}Qt=P9-s�py"���'��Ȧ�4#v���#Za��~EN������K9�hAMv���R>_4f��S��$��6ˀ���{	}5��^G�6���~�w-��U;|�=���+���y/��P�U��#j���@�{��^
}(��mKX�������o=ݱ=���(K����$�Ò�!�����	�CP�A�$O�����u=�i/���}X,9�&2/F��
�h�+Iw�7
��O�i��҃�)�`>�Q%d|���D.��/Y��h}��FB�MZv���.�Mt5�d�N=�Je�0�#��W���}��-����yx�N�~�s>��� ݉�p�5t�dC=�c.���.*Ț�[v���L.�	7`�F�<�I* `�<����`�2��&�D�3Sz�U��q��. &��F+Vp��7�Ie�Ars>��+����	NAGCt�&ҕ+Ww��9����}�!T�Qa��|IŨfM2P�\���	�B�gB>+�b�����q�����k��0ϧCX���h����t�g�v� �"ёȑ��FlƖ	A��L)������J���Si3
�N7^Wʚ����`�����2!�ч��X�|�����.��/�	�G �%�Og�g��_���#��n�܅�I�alP����:JԸ�aX7[�v�[��B����%�i�=��"2�BV�ļ�я�d�n�mh���́���d��
@O����Kݫ�ܭ�&uB+Y�8ZS�HaV�1�ɵk��(�@�ճ^ө4	M,���
�GGG��h���lL����5"j����1��(�c�q��Y��-8_q�p���r����Ny�;>epy�
�3���w�WF0#��eޡA�\���20��М����r�N�E��%�Hi�,9���4o���_
7���ɱ��&�S������prZ�o�,��-;;�S�,�`�6�J�'c�q�g^�����\~�Ù(7���m�m�r��K��'��;w=�Dc�$�� ���:���?�����x3rd����7�e�����?��������SZ?|��JWU��N�(����6���VB;�t����v\]�:���[�x�����z���'��Vd���"��/�m�"2��q��N�ٮ�W|�9�/ҟe�y�XH�q���AMz@��c3_�@|;pHn|�v����;w�������)�`Z[)D7��k>��8�n����. �z�2$��\L���g(|��Sq0Vو[*�E-!��C�Z�F��竩m��!�]�吪N�s�k�q��y��\���i�<}���ЃLv��(����`U�U]��t:��MAd�������|�q�	Pм��3V
O�C�d�|�?�����l�Q�q2�}W���EV�mH�L+67����/����捪S���\���7�q���E�2co�ᒜ��
|ٗ��_/~��(�'9o�<�<�kd�[/��'�׿y��p������x�NN�FjM��X�d��!t�;�eJ�z�e92�E(��]��E�
F~�"=Ӷ�+"U6�9d��qt>�u��7*{��J��H��+�:���wk�U�w���z�3^E=G�����J����3����"��,�B�@Ef0�(�$҆�d3�x�0��b]��>:�."N���v<�{ua����?H4-v��4��DE̓2���8lUgQ9�/H^B�-� E����'�g�L$�PHWN:|z~vz��N����w�y��d�f�!]'F��%�����5� Y��kd��q��#��/t��0�;p&c��ie�����'��R�C�IOL�J�F�����X��G8�J�w��� ��y�7�3V�
29ټ���W���H'R�����������W�_~��'�'��~����;�2�K����!��9)Ճ}R�ުCy�B���%M��~��e�Km���6���y��H��f3g���d�@��j�������'�~��&��M��퉫�zG3�hʹ#�tt����B։"3���[N��)��M���刕H�}[�f�j��=ږ<o1z=�(�Ɛ�*�M�"EN���+r�L�Ƈ>�A�����xo�k�U�)𷤑-�����2�u�j�)F�KH��ґ�>9�6n𦕧6o9�66�@h�����슗�"�̘F�=#p�_{7��`��RcrsO:�7s�{��c��
�-��hx"߄ ;�Ń�UhUV���}����qN1p��.47�i�B��7���#�H�ȴn�ȍ�y��������������_����W�^��O��2�\T F�g��F`�=�;$��A7�hR�\B���!x�MPk�s0B)��ʳ�q!Oz�t �"du��j��/4 �B'F'�b�>����Jo���֪-jo<�@ǡ:W�#d��y�����.��_�pS�
]?R�G��{?��a4ژ�6${Α��J����&poa�%!ѧr�H���ڬ(�#��1�q SR�ŀ�&�OZ��[in=ί�r��������U���,F(���s��<��o����W���*\�ON��X�L�E�]ϸ/|�*�X��ϏB���6�'m"�l��p���X E�j@�u��0��� Wo �o6K�d<��\����\D�+�b�3á����#�=����@
Gr� c)�=B�:�N�[>�k����gk���int��VQ,�H�g������#���D,%Ա�U����a����<���|���	]�0���9�d�O�l O5��	��N6����޹P�[�5��U��G�LNF��A
]:E��K�Ѱ���'�D4^��͆Y2�uh��[3����\$��yA'�(����]kL/԰������:��Q1آx5��g�B@�AN=�c�8[�r��$`kC�t�`�q���[t���:�(0;8��}ܺ}
�fő��9%~�����뻿~�����O�<��x�1�q�܎r9�MsK�q�¹j5
t�(���X���S=,+/�/����q��å�3�)�Hn(�̔pWfi��D{r�9��J��L�#q�@,�Ѭx ��|'����,�����p���y����UO��t]�6ȗ�3�zey'l�n)��p��m<�����J=T:U����g��JԎ�� ��kj�1��^�ZM�ԡ-���0�@^s��HIT *	��#otp��*���G�|~�_�
�${�	x,P:/s�̏ĸ?��ϔ�m����!�Y�"���bٵ�1ǍKN#����$��Nb��#](o��G���`THR^Qd�OUˏS� ���ۚ�3��v%�<޼*E���A�K^�����{�j�՚����)�vI�+-:8�e>ݜ�3��,�v�ڮ��,���Έ�B�^���]��red���k��k��IT��&�8Ҫ�l0<z-"�,u�vcձ�o�Ud=R�ǙhKG���l���x˛�|�Z���
�⯷L�#�݇���ѫT��4����Y�!�Ķw�Q��0'H�cי^���n��ObhHI�t�t}(�Ȍ[� ���TN�qe݆�Y�b�%�&::o�9����kh��J`�{��g��S�r
�ҁ���"x����9�h�[t��9:�EV!Q5Є"L��m9���o�s�s���uQEg�&?A������N�����:��\���ԟ����"��Q\�����`�������N�!	h��1r�
^��π������w�~�g~9B��U�6��X��}F
e��ᖦ)�;�j<a_��6�4=���}d�HЛ���z��,'��^��[�-be�Wk�=Vl8���WƘ��ѢL�^�:��~���{�c����i�A��`������+įr���~�q�5Tt��<�������ɑyz���ꆤ e/��7QI �`	�EG¯��u/��|��?б�*��'�<-E����%���O<?�}?{�Oa}��U���mF��!�1Ñ�\=껓�����i����YHG�yA~Y�Ӂa�92e�7f�b��}�����W��������2��}t���9�Em'��9����Kf">Y(\|-Ƙ�W�g���4�X:]s
��+�>W�L[ʔ!��)��?SE�<���	�D�;2b1B���y��H����;��g7���~����y��7ۛ�ʵ+���l���u3�\a\܄�B�2�Wa$}�S�[7��A�n�>�9��A)�˱O�pr�QXɝ������*
h:6��6�ԁ� Z��Y��j+,7Ɓ�8�*VSq�N6��h8�6�ة��ywE�I�<;�	����	����w������{��^�
q���NÀ6x�PKxB�y�,#cn�X�����V��NKc�IW
ː�c�w�bg�K�٢-��2ꒌ��/�)��R~Jׅ��C2�+�����Od.�_�yŇ�'�G���>�}�v�Hǀ	�y���޵�=���}~�W}����O����9<��ch�?�zgn
��RG�W̑,��.m��)9����������E��A�
��\�x��l$M3�
*�\Fb��~�=>�#�++�|�U6��X�XI^iXsuN�	
�<!}�`��&������8-l5:���Ѯ,��4Ar�(q�|�R���z�F�5�@J���	uF3�rJ�"-8Z�8�H_�Fd��yHF��^�0m�xO��cng';���	�t
s��%G��!�v�WZƀ�uГ2�\n.��2�h�����!�AW ��4(�EY!Q���K�'�,%q:ɢGT��^�J�(Ɖ,�>�pb6��n�8�}�*\�������L������6v}�'ɍ�z�-��3��W�[B�+7�O�٫>%8�^�3�"bf��&�E�Y�ː�<cr/&R�5Bk�|s��:xA+%�#�Nk9gn�e��	��F�����B�b�.�G�h̉��PDvc夲;�Q7r Á'�x~~��ۿ��ַ����᛿�M�i/�t�CZC�� ]	�"��d@�˝���Ϯ�:|'�$KF����B>�uekc�H5��મf)��J��̨�+�g�|����G=Q1�ܤ��]����*�������o��E�+\9Gz*:7�~��]�韃���p��Mx���Yr�ŗ�Rd���٬������q��R�<�]9F��T ��W�&���f���K���L+�q�5�s�m-�+[�M|����n�������*@yH}G�&�d��hu��$]d�K�HbSxFu��gڊQ(�ڒ���k_�_���Q��v�ƭ��K��N��kPnh��`}�920L��OOD��<�k�FSt5y/t�s�N�#^؟׈�D�!�<*��3Ĉ�� y�3�:�,�@�ס�DQW�W�H"W��p�veW��"`���o�� �8�Ľ�ФV��t�*5s��r���'� �s��Sh& 8J��kǵӿ��G�p�(m��ýH�kuP����;;W`4�a�NE����(6�����/��y�$L�ᩧ�2�Bmlt�ϭ�C�����⼑O����d�M��x�����q��O(�F�zzr~L��On߆ӓ�t}Q|=D��s�{�����~=��S_
��w|��=��33Q7�� ����
X��ё����6�*c|�T�=<����&����q��k�*�Ŗ
�S��rި��?�����J+���?h�_q�`�Эe�Ǽ|l�}�r��z ~��������3����=������\W��m}=Ə�^I���]�T���+XTΌc�$.�\�cF%�-�w
F�Ɖ<Sh� �K*�u��8N�����+�uz�]��: �@��h̩�����aĥ��~�d����?�޿�M���G�&"}�9�lW�ny]��Q�{�dN� ��,��o�EM.+S)�M�a��6��}�c�"�g���kEǲd�'��)�\9A�1���[7?"�:p�F/�5�!Byߍ>�T�j5���'U����Ђ� Q���}��
;RO�_ݠ���%i�����3k	R6A�7ٜ*���`1c�"܊1���$,����n�����y
���9yԐ�!l� Fu�}�mO<�~�)�r2�^yO{����K�]5�lm��L�����Y�쮨��T��9�m>��P�Ϙ������$�rU�U�Ġ��m��E>E'��'>�	x��c�=
IH��^�rL��xR�2�+u6Ip���,��o�Aw*�j���U�KgI�f��}�9T�T��5��M�E������c*)���A��;UI��!� �^
��B�S�4cM1�ЯI����l�}�&�ٛg��歛pr�O!�#?�g�[��Q0t�)yQ7�L1˯�R�]z%�����g3����3��&�:?I�r�`WzȦ��J�'���S>�^v�
��hb:���F1{�Æ|���lJeđ�;�A��b �;�yV�8<�̓N����te;��2�[��\�%u�m�<��*/��/�~���28����F�WB6�}�P�K�K���r�/��_o�ꢫZ:6�)�T6��M��I���*�v���ϟ���������w�oBӘ��y�K�������o�* ����f��>@֡�@NeNNN�֍�1��t�j}W�\��s��>�_�}�s��·s���ɺ�s[5H] �2_�=�5��cl���Y�.tw�Y����3K|�z}��X��i�c�R|��R�pI�]�)����~}�K�Bŉ4��`�>ߨ��2ڈk
i?�
��t�� �n߂Gwrh�39Obt��嫝�	m�N� ������Vަ%2�	N1�r!�ö����3������/7	/��c\��k�|	"1x�%F��~ ��.�1�	B7� <Z��xd�.��?�y�;�O?�'xUD
{e���|y1F
��T�� F&C�:����|���+�:HWo�Ö.JgZi���I���.&&��U��ar��?)��7	'ĉA���h�'p���wע���ޓ�C�䕨�rc��{��3X�{�}�n�܆�-��g��|���W�r�2ql���F:�J��c�>ЉѬ�!��Sv)�#���cV�z�c�6h�⥽��Y�i����i$O�nF��a�`T�d�H�ԃ�t��T��r��K����^�s�E1j�_�!��z(A#�9�ÈЩ����9!ٯ��p�?�'8��A����kM���R��G��TWR���CҼ�(/v85�����9|����~mP�^�m�`+����3��f��5(��c9��7��7[�AaF�6�o�>�骙�3̓����@�	��1��j7f/|����^������m��)}*xh�{7d�b�j���a(��t����E;5���ʯ�DD����`� z5���5e_\����'3�ù��>�����p �-���8_�۸^��QZcg���O�G�������ᕯ�,t[�ӕ*���"�^m�[�\�e����m�C����-��T�2�os���ƅ�H3 ���=/�ߪ�_�k��L�u�h?@���=��79aH�t|�IT�N��v��O�_?o��_��9'�^�"�>��u#�X�(pH��e��ܜk� ��IJ��7�RS�|����x@���Rf��&9U��-Ӓ��7�s��&�&��������8oh����s�����g^A4'�Ƙ3�1�ZF�����#�g��|��۪k	1��3J�\�����jw�VE|��>��"⽂��!��'�f�t��I��׾��7��߄��y�č�1<l��1yTS�?�g`%^8< �l����MA;]7�O�>3��<~N$t��鴉R��2���l,�ge�m%�<� �[�,ޓ1�`����Q=�O�̵�e2P�ݬ�@=ߓ�r}t�z�'��}۷�'ҳ�_��-��G?�Sji�3ݥ��=j{�~W�~�����<�����Ҭ��9��5�����3��Ro(P���Z��"�ȝ���@�]#�=�޵��|�6�q�;�~�V<.*�fE�!����=���:�0y:�0������7a\t�H�KA����r<m�Q�bh���/����[ {_k'�$8r��Ν��[u�ٸ�FJg�">F�z�ޜ	�9�!|�k�"sP�Sxg2�����Џ ��ň,t1�������I��А�r�h�SPx��@�A�Y�x����L4%�X4�ZƁ��x-�@�7 ����6O�B'9��<S4
˼q"�L���!���}��X��g��-�u�M�'u�ǧ?i�9��`�FM��V�E����;���t^�2����kV*��;9����)��񎾤;r�w2���(IV�ii,+�N(����lts��)Gy2*'k���ϧR�R��tj���`-�;�ʵd�CRM�)��^o4�C�E0;�#��u�t�i��y-֕�p��3��3�t�nM�����{�W|�g���w�{x�^7v�M
���7Ё�����پ�Ml���Aa}�)��SȪ�����i�..[�wNǩ���/��������e\~��V3&�P.R!��������P^Hn�;~��g?^����>?���_����70���*]{�B��� �R��~�e�2HO�ǠB������ӳձ�Su��eљ�t�ͦ�+�<L�Vu�q�Y�܆�L[�Ӵ�&���4x>ۭ�8d����P� s����A�:�~w~~�z�8�<���x}�&������b���#��$:��U���Z��v�ΗԏΕ��F^��Uk�X-6�N֣��������{�,q3�ω�.6`���t�Ha��[
��װ�~�W^W(u7N�P�8�uj���y�mL��v��wӓT�#:N�Ҍ a��q�[ۃ���?h�L�������T�i���Ic���0_JWF�+η�+|8�4�"��!? ����TPr�6��.h�22�~\r�Uv���];��C�n*�8YFҖ�믆e�klX?d9���bE>��aI__#ON��j�vE�$�DL�Z�No�La�B��4���q���j|��n.U����Q@\���I�>�R��A^.o�C��|R���Q�>�)p�(ZR��1���e巏\1��*�s58��k|9Qm�=�7$�	��6�sx��N�g����=p��w�&KZ#7����fǋ��1���Z���.��+t��җr��֜6����V�ۓ�8���)��딈^����u39-0�N��=>K��S��5E�ڢ-�C�m�;�g�����V�w�Z0<����uj��$�n��E�B�=Ӵ2�{��
}CQ;��̟��L|�R����|��ӡ��+|"���lj�i���~c�����y����_ 9�h6W����Rմ���q1
�S���>�=�u�$
�����@P�̀���䵁Xt*�ԉFe�!�\�ʫ<��|*r�تJ/@���E�#�O�=����CU��Nb@T�{t޸z�*��[����7�rW�]C�`˛)��qQ�z�S���dj��J"�����!�Z��|�\ZrOYI�/��Q�_�8~�{NHx��0�;V��&�hC��I�po�;ql�6cB�S��\��'���Y����߇��u~��~�7�F�[�d���t�s
���#�#4t5��O�I1O�J�/b�*�x<3\����� ���9P��K���9��\�l',�3N�������Z���)tp���?|�{�+��둼�W\��Y��pޯ;`�#�I�qo+�BԓE�&�BQ4���j0��C�|�'%O����I�����r2 �<�(m�&Y�w|J�*�8�A�F���K=�0&�'�E�A�����o�Od�'���t��'��ÿ1~� ����`%�0�J�P���y�=J�F��%���� �pO�ad7^�F���-��l�nn�}�":NV`c��!8!}�q�}*Zʳ��>�	1��#�Y\��d(�l$jGm���d��'{��j���!�wQ3��6?�*��Tw�Jyh2�;ӏ����}���?}�N��X'���_W�_��u��"n.NS�>_(�*��ŜdAG�x����&#��R��<sF�}��su5�4myFynm�㡿B%�r]}G��mJ�L�(e��2q�(�s�뮻�{�7��}���s���D�`�N�%��+[=̰�k�Fzq�,T?�q'\>o����8�s2�!��:KR�ɦ��o&˸̞��x�9FG��|���7��@�0�Bȯ�m�6�t\b�(`9��z|�
<����%�y��u_
=�Q������7�Bv�t�;ܜ�y��ϲ�����ӏ��T<�����.���Z�y˶��>j*�G�B���S�}��9x�vs���U�Q��;���&�c�~�_��`���dڐ��y��ɒk�c��*�@7:*:�8gl[:0��<җ�Ym�u,��'W}�"_��Σ��_ �������{��;����v{w"iOG�8B�V�\��h��v}$�B�W��G���z��o��z�_E��s)��M �̷+K�c�D뷇-�ڹ��3�q�������Sp�t��n�.������f��ggu9�{�a�����������o�����������r�FlE/P�K��C�M�(� Wҳ>Zʮ8^�+��*�=�suP�ޘx���
SG�/�NHQ3�IW�<����o�����_ɚ��BM[ٟ���0�W:�R͞;���Ŏ[�ϸ:��pP�������Vn�:�j�P�C����8��O5��.�<��
z��yFM8;���杣:bd�M��Z)v<��%xOv��h��_�����+��q�3P�IoS��ĩ,��o�xx�����ѕ���5E���h��i�,_�c>=Kx��˝�K�����p*��Y�P���������5f_�������FDr�P���*������� �[899ú�~>��?���sv6�nsv~�������	��C��㏢�P�=ur�4���ؔ�~7O+���mZY8v*�v�2�5j���h�I��`J����#݅L��k��P��ik�z��א�%
|�������6k}������`#�> !+i/�#�Y+0�{8��;)22�L�e����G��"�6���t��E�B[���lܖ�ͽ��ʗ�J�3ؽ!���rG����_������_��tJv��t8��)$l���0v��v�����]VJDa!�6zU��8�Ԙ��l1a!��AԻh��2�����	�Y��PF�@��L1t�!@�.ҭ�7�����Nʰ�z�9=��H�k'm��#��1t��#�s��9e�pCsPˍ'R;
��\��^DJ���2p������x�����?���O�Ǩ�.Ϫ[cy��0�^�F��Zݷ�Y�͵1U�e�Z_jF�;iX�c}�><�v c&��ƈ���7��2]^NjO_���hk����/��+G��׽^��OGeE`��*��� |Ŵ���nݾM�oKOd䣼H��5��� |�� D!3B�kx�<-ruf���m9��ѥ�m��#�)���`�
���0��ї�iZ�p�����ø�.���m�Tv��N�PF�:�G<���9��{:'<�3��dk�C��(��˔-72E�[���2A�.d'j���{]ԡ������%�~������d	��r�i��4��mu�1�
j$�2����JH��5�\0����RF~�4E�鰎�e�B!N$2��&����`���eD�9Ԥ�v���L��3j�tD��6Y����_�	��>*H�7���kh���M��^��w����w�������˿�hP�W=���Ou��`�Aoc����I>t�<`z�4kr�Eu�R>���FM������E3�v���J�^�3g��(ќ�Ӧar`����&��o�F<�y~�Ά͎V���&t㐝7$��n�ິmj`LFN� ���N��N�F���(���mة�.�ad���N��t���e��-�V�ɍ����^�����"�����}t|Mt�T��A�IC�2�:ܴ�jzHʻ�|b*�ƽy6ob�}�J2�o%ʪ�uJ3W>8�쬤S�is�y�.|�w}'|ŗ���;��;s(�`��ΰ��Z�w���>��(0d9���akz*R��7B�y"��7빤�����xNh<���O5;aN����m������N����_~����g�������{P�I���i7ٍ���UA��#x�N7x%�ȳr���������eZ���*ʳ�p�Gp�[h��Y����^n�+�`m݋���`:��!s��J:>h����<���6E{�{Ҹ���y�ܑ��t�Da���J�K����h�	��-�x����zקr3pߥ	���M^�,lEhN�@ӯ����[x� �M��t�w�WB�/#{�C�X4&���|Л>D6-�g�D�he�y�w�n�v��e�Yc8�^u�yW�"[�N�:��%�C^lL�"-%=zй�1�$7���n-���m'�B�(X�^i#�z�8�H��DiM��ktU��=��;B���ӓ3x����[��k�s?�����yW!$����(���rF�#�Gj�����Ɲ����Vm�C�J����O�K�/�H��r�|I�S��/�O�������js=)����f٘��7)e��l��9���em��S�Z>����.���������u�}-�w�`�㥷n���X���F��������zܸq�	�:,����m9��E�����S��9�5���t� ,[��dʣ�-g�W��_���7�O"�
�]�,������l��'c{��y�G�No�Sy���Wr�h� :�s��<����E"r�z���st��զ��u�5:z�k�P7��w�=����lq�����w�=w���9_ ����	n=~o��_����?��?�kTx���qN�,Q�E���Z�.�`$g��D�e\Bc�SJ���@�YM��>Pꝵ�5��Eq���8v����ʠ�%>do9O1�M0ǂ��*#pd���K��z�K���B{���#&�~�[kr/+]�8x'�Ms�٩1�2�.�k����G�j�LF�m��k��y�����R�}�1��/�?��Na�
99A����P9�F"Lw�J���]}�}����tw{z������f��90o�d���;�is3�C�=�BS��� �F3G1���0qt 3R8�u�N����(9�,��7J���`y�̑1i12�(��irv�H��=*7�W ��%�'�9X�0Gݪ�PGɀ����`�B�dz�~`�4�N��Q՟vT%�#��l�OaH'tV)������g|ڧ�y���N��kv���T˒�d�j�th?��q��y�C�qo�dcCd��ݪ㌬����,�3�6�҉�d�x���O~�G���'�˾�u�W�
���ϼ�x:>�,Y����&�v�vn���~��|?^k� ��Sx*��Kt1�j'���B��F'��ޑk`Ci)�|n�����'#����%�fNJrbM7q��*]!aYC
x���S��1��i^:y ��Iy��:i��=���#w m�t=�%�hܚ>V~�+M�LS Ul��"Cg�%��y���*��q�det,<���y$�Hdޙ�J�3���I�j�"? �N|���[��ec���'��<��"�O�y��H�贴%�t�+��<p����o�����S%�n8o����嚠��}�N{Z���c|�^i/��#�����q}�X�K_���wxw�|>����m<]��?�xǻ����V��G���1��:m@>��S�_��~�To�ͥg���P�~���t��:-�{�{�3�F��Q��n��	�Jtm�"�_x?|ѫ�n<�t�^a�ٞ��Oz��j�����ρ��h�&��(YI_��%#f�{�s��H���ɑmآ�s�׶l���hh��[A�:�ُ�2}1ãQ��*%�hF6c�.J��_�Q�CBp�Y��x�G��8�6� ��.�;2������������韞y5�8��� �׬�`9�N�0��F!֟�ɣ��� �F?#��PԖ�A�*�i�n݀O����/x<��p�d��J!�A5�Lϧւ�g���R�ʃ�+]�.��ҝ�_�u�O���JQH7��5[��f)-ەb��J�>8���� |�~�d'�|��}����
�z����}��I�$��uIx����ǟx��G�C�ۃ6 zK»;~��ۣ�C��y0��n��m��c�Y!�w��n(-�3<6�� �X�0Z��Nd?���`�9$r ���CR�ҦKǛJ�m�p��w�̕c�u����=��&M�w�c�.��P���w��pŵ��\��/ =
����D�@u�ל8d�kR׆ו|yէ
YC�Cut��l��kk�H���A]����w����G��l��$�Fd ��d>c5�%�����kK�-u�'��v��~�2�>��h}�@~k��;K^��E��ѓE��%�Ǥ��������hË?��ݏџ�>٭p���W�"��� ���wû��n�IW�v�]��i ���ƴ����Z�X���T�NQ导�����E�KՄ��,�3�M�đ*�i0�
���6z`���w.��ut���Y'��K��q���#;Q�0���.�O=˩W�^�ox�7�+?�p��	�!��Z�R�#�+�E�&[�
��ʌ4�����)h#��Q���ga���J��x�H��h�����$mMw�E�(�V��wz5��w�>ԩA�A��ī@��E��$rGY��2:?e��� )����x��D�Ň�%��̡\�'� �Ai��'��yC"%�}/%����P��H�[�=�O�ON�>z��}p�������
����v���>���<JY-��I��>A�jk.+��q���$���^KaLd�|R�Gy���_���A/+�R�,]���t"�:��*�@�KT�vֺ�UX��t�X�j�qa*�9c����h-_ZǮC�OW���IL�z�9���m-�k�OY��=�����[�m�ۿ����]�ҵ0�b"ʗDQ�P�RRk,}��/1�� x�t�`��!�j��H^�iE�&A/(c��$9d�/�����?�{����z��l,U�q�"������G�j��LN��Wk�q=���M"�6y�뽥��wO��l���@�I
��S���Z����!�"}g���=2<;��I�tb-9���o߆��Pp���'�)_W �5|-B�����ҝ��M�v�)dw����2����[�0�wd�"dtei5�����v9=�'z5O�6�����7�"�D��>��5:[�w�UZ?�3�~�~n��]C%���t,m��%'��8���Jt��;�����D�j�jQo|�k��ׄ�1e�G�Tnl�"��1�wRJB�X�`' ��-�ë��1%���T%�X��x2n���4i��P]{Nճ���|�D�5����V���Ť2��&^�`9�0��>�?�ܧ��q_��vڂ6=��̀�]�7��햍�8��jg1lƐ�jp��z���l25�*� ���]��G�-k�ލ�(�2�[(y�m�	M����_#Aq~�+�W�x�xk��y'�'���GG�^wp|�h'?��`'�y/��G��QX@�K��tt8)�P�Eߗ�VOCZrĜl�Ƴv���j:�\�K�cZ�k4�u�Z�j:UKo�|r�� ��Mo�{��P��Oxw�(���+tBGw9B�����ۭۘA���9�D�h�:Srԡ�Y���R�>d���|�}���w�ޖ�����G�Y�2>�L�����A����@��v������������6)��>��+L� ��ӈ�"e$ܬ�IoI�xs4�W��!N�L�W���̇��!-9�����9::�<��;9mG�����G��GW��07{�?��^��T���6H���9���$�xƓ�.��ˠ_��2I`�^t�pYG��1VV��\�B���<���V��!I�H��������Gv����j� 6�5�:mJ�}o޺�g�p��_�z0ZA�r��!��c����ֳB�����o\��L���O�OĈ���m7L�{��x�$%ۄ�穝��9��>)���$��k䨭�Kg �*!�(����@2��;B��G~Ǒ�ͬ��)-U�E3^�ϻ\W2G�8�q��_k�82F� "p�����6($�m�$�>�J�ޕ���j�ss���8�<m�V�\,�g���s5>�7�˵��r�J�K�L�k�����k��������JI\�Q)P����t��+��!:N��F`��9��~��b?gb�ӗ���}SN�V;�����_���Ȳ�����l	~,�ۖ�Pʃ�O0��Y����.��[���BH��9�|�1rhbgv��!�۷O����/D��-"�D�JI�k��1RD��z��ˢc��fP<4҄p�Tw����"��J�ɾ�A�@xEqa6AWTo�	"�}�=%����Jy�n���煎�;����u�qP�D;���-�20�kkR^���N��>�w=��W��l��k�U=0�U\�]j�s@c%cD��
�&��t5]�Qw���]���{��3poh�:B��g<�.��{v�9�?x�;Б1E="z+N��}m��;���~	�g�g�r�pIk��4�@Z1P]�(v^�����z��.��y���2oE��8�����Lvr�+T��v�~��7������,�3.Sa}a`�؈Y���Ԩ�6�y����MȮ�+S9)eQ*c4e�,a�1����b}���7���c���^R�%<�0�ᑌgI1�3�dI{�(O4e�{��3>�%��p����!�����Ղ���@8�ea�b�(�Ɋn`�%d��ܸ�=�UR�\�it#��ۉ���)�VQ4��G�qY7�q�R믚	� �7҆b���l�=�؉�h��`c�7�@�s�T�(є#}���?�rN�7)�7I���縦���RZQ��R�R�,�+sY�Uw˹�%<��z�Y#7"\\�P�*� \\@i�<�41�����8��A�Yf�)�3�/��3���QR���p����9��nI�m�6��A���������b0K
���jl�����WY�b��󘲼.[U���	�y�P��?3�kt��GE))Mr�joY��u�h"�E����g־�)�[���aK�������/D��J3�ڦ��[&�2��	��4�h3�D7�2�!�
^��n��x	G�HqJs���	��1�%
SP�[�5@:���Cg��b �X�z�R���ph�r�������!��5�T�\�C���qy��4���Je2"F'�S�۷�wo�j�Ls���UZ|�)E�
+<�n�{�O`�9��o_P�K�ƒ|��d͸��3Fy!��ֳ2'���ޚuN���a)�_�Ѱ��8p�r֒M�)���\�M�T����|2J�h��EEx��O�Q�0����bȕ�L !��:�Ǘ�P]ǝ�e>�ǂ�(bPz��;�șJ�V�h�8�$E@���H�pm�|������O�m�x7�p���h�}�R��;gJ�2&����7�G|��֤@�7iL6[����:�N�|x�=᧝�z�I��s�<��5�y8:��z,�o<�A$��w2�cY	?ڠ��uך��<�k�����VWi�{2m-��բ�-���݉y��֖�?eǡLU�'�^���2�S�{���ohw�z|��>0���y���Ovr>F�Fk>E�v�
��ҵFk��QY{���V��j<\���ȁ�kn�#c�}�hLf��bL�;�` W���6��dR�7�BШ)mՉ�df�eQ�t���(���(/����y��Q��:�E�^�Rf�G4���d�c]J�Z�6iĞe��a7[̓y�p�|*lsjpu_�ȲRpt.��c�-m�*^�Ζf ��K�[�0�8?΁گK�A�n2$ÒEt�(ϓ���դ+:��^ �%/�<r�2��&��m$�:%;eVpz�����'rp���a�N�$��q_�8�,��>������}����f ����nR_��!�(��t*�BGl�_폫oQ
(Ag����x��^�]��a��A�|�`�i��VG?����)�7:^��͛�-� ���V6O����N�;��������y~v6��t�,�?x���$�T]��Q��|:�u�L��*�Q7��������i�&�3���I�%��ȩ����u3i_?��A�k�ȳC֓��|�q��<��z��QXrx� �/�G�E~<}"G��&��yW괂s��=�e��t�/��G0�M�-����G����}��U�I�K𜟝�nr��'sAWYۘ��z���r�JL5�@���J���9��^��]��{�1���	����]K�Ј���������/F|��m��m_$�9&��
i �f6y5&$�F�M-�ѿk�T3ԍ�!�����u'Ҕ�+�k�g˨�:��%��)۽(EJ���Oޏ)�VJ�A����U���x�1T�9�@LHI���S�>i�s�]s(��0$��2Ȋ�)�]�4bX��&�9I�ޝ�qIć(�P�'4O��Y����߀!�DYFR��B�>Q�9Oa 5���x&?F& ��O�Q ��(�z�����( �ot�	���FN�A����l��R�	���˺>^���h'|�Rܑb�"k��sȚ�P���uZ+���2���"z�G��9ZP�S�hG�s'�
��~!����
S9^�U���d)�fm,�d'{i�s$x)��]̡��L��{}�Yi��nZ.����Ewh�)%�Ok���E��^S�;����iM)�����φ�ceK�a@Z�w[	�e9JdJ�\�I��>��lP>A�S��%osU�5�$s�҉���N33���Z���� 2��hLj0�2��`���L�r1���[��$����� �N�CN�����?�"s9ld��i�5u"d��|����u�����l-*��sS?���J��/�u�0�۫*�2���{��.��;������ �JQ�ư�ׯ��Ѻ���z멄oJ�喤%���}�0։j�嵵�$-��ke��9�v��t�Ɯ��t��>)S�_|}����su��tUc2�'�t||�0��w�m�y��(�CGQ�����ǧ�E��BO;���lAO�9D��Ic�tP9 %t�fg9Z���
�:d�qd����r�*gX-��qM4�m#���:��~3���L5I ����.�C��!�����!���o �s*�:��7:��X����>�R�ez����g�?�Smi�SG�q�ǚ��t�8�����<�d�%4���fJ1��i��|{K��)}�"i�3U�"�\4��.i	߹����V�����Е�<��k�D/��-��Ȫ�M#��Hn�m%n4
���W	�8x�C��4�c�;�/�+?���U.g�֥�M]��&�'�t�E"����x���,3���^�����@��7�J�k#�s4?�u��O��>�aJ���� /�FP��S����ۏ��I�A��y�h���۔G��z�2?K�^/�w������6�JG~�9���W�~?��LuǱsN��Ȝ���:_>.^��i0ߴ�dt���k�ad��o�I�i��ގd0,�6��Z�S�	 z}v�u�}U'��p�#L��Ϫ> k@��CT�7��.�7�!�7����0��Q���p��Ш\��T��ed�fW<X�"��mU����{���(� �l�y���\��X6��a"��xM��9:�%��&]��=�o��Y��`�6�^��	 �Â��N7�sg�E�k��RV��Q�sf�ˣIEצE���R~����@%}�0�+�גq$*�Qxl����J�j|\݄��)�G�O�<�O�F����x%�ɑ��#>s������wl���K�"�D�)��&}8��_rFGgЄC�����  ��IDAT���+���7J�Uli�s�y�F[���VG���U����C�{��P�ʌ$O�!����W6&��,%f{~��<�E0&��9y��~�Ju�^r��3=��^�vL�#.A	\`�%P&��F� �6a�����0�
����H�m�������'R���εU�q�Of�R������p�$�j��(S�_�Gk��!go?1#Q(R|��n�b*��B�̙-E���fH�JS��gz������={l�L��>�ۯW�.�y�O��`�8F��]T� V�yӪU�S�<��Ǽϕ����o.���ʎ6���`'P�L=c���c��nS�����-.�^9�J���R��l��h�>m.Mc�kC�^�������ɢ�w��%u��l�E�Q(}��y�ϗ�ʳ��Լy��B�&VGl��	�k<lan�u(��YO0w�h����Į������ysi)��x��c���7�^q���^��WHA����{<��>����e˶s�,�����Y���t퍳�@.�v�ϩ�*�څ�4���2!�#��fւ����2�U���F=!��W�7W FU�K^���)ڏlsʉ��,_;e=���$󄠊���Tj˕0z^�--]�(=��EM����WKʴ��T�a˸8�Z�ҘFۜx� f�?�o�k�%9�]d }�D����œj9PP��xo���x��Ht&���AX9^�x�������;B͢�nI6�썴����"�1��4���\�|)}�\�SsI"��`��ab1�k)�1�C�����5c������Ƀ��`u�M'���r��1�Ӣ?K�uu�(E���Y�e����j�E��o�4EC/Zϓ����ڼ�i����ߌw]�����Ж5��Aj��й�9c��ue�L"�<��\_�X��n����L\�+G�)�{���U^W*�JT~C�߬������D`-�x�'׃�3+_�@�2�����B�P�Ǒ!��f�3��$W���Q�@X�q["��-�b?���"�hĽ�žt��+L�=�Ü^ ��h����퇎K���ar������ X�,[�kR��aQ|$Q�Q8*udk��\J;c�CӎYp?�������6����Vln�m^
LA`l��"�1Ne��J�^���>DƗ�&0�j�0����
����U�4��������]]��H���tfPz��8u۔y8�08:FyrZ�Y���b݋m�ܟ:hť?�_�-�O͍/4�a�r�'��7�o�Ӷג�%v|�7��Լ}F�K�1 ��^�+������R���k/�q�WA`^�!KB	m�7��ҋn��w�.#$�\�jo��[PW����c�F4����^�V��J�m'S"=VJU�s�I�ߎr��k>L_a^P,4`o����X�6N�:p���Y�����-�>J�X��,A�mZ�� �T*߭���c�)P-��^F�`�E*to�I@%	?g��d���b��w�.8vѴT?$�E��.�5'.1̥�Cd���I�
m���A��1����)$u�mA�3�˦=-er�ᮜ�R0���9���;�����y��PX,𦡤zv���+�ˢ�P�/s�D�vY_��0�Ҝ�fi޹��z�4�[-#�ʱ��)�y�h��)r��;�/�wਥˤe-�Tiԗg��-ܝ�Sy=���o�H��Y_k�L�5�?�Ұ���ó�R��?j�Y*�F���Fƿ�����4g�k:�B�.IOG=GR�%�n
��X&7�\Q�*g���E\��ճ���y���u
o��e�'ϕm�Z�q;��0|-ӡ��t�/Rwk<j4�t6}��`vN�4]��!�X�)ԧx�>��/.�\�Oj��S��Pk���T����T�Z[�LW�]��ҹ�s�9%�Q-������t��쓦��'������ev1����ԥ1=���6���hI�Fʲu��-��R�>\�V�dZ[K��D!�q�G^�5�:�+��j]�Y�� @���{$�h�?�%e��ӾQ��H1�q���b9���_[})�@����[�ia~�&��D
�&��:~|1�˳eJ@��@����A�`�<�z���������T����r{��	�W�'�%]1t=�;(�Hn����8b/��$�Ef�(탛"Bv�)K�Eu�o�F����$*OjKgj���ZW��ʚ/�t�3j̂r�Y��tlL�y�S�΢h, y�t��(т�+c�HW��`<9o�m����d�`��t �:LP�n	H��r}�ǻ.����,�c��;)ܿ:��h�����JP��~Bѵ�H۳}u�vJ6)S��9����
=Hc �����8���nE
]���b��&l��ڄM�k�k��]v:d�.�������zfa���s��R�K�H����.�C��]�,h¥7��#�_n��LR�N9M��A����Z>�V��xg�Hh��r���EDI ��`M�o��g�\�E�VZjǼ �zk�0��bPІZ�Z�6Zt{�q��l>m7����h�0�͂q\��%�G���JW�)��fZF��y�O��'�	�V���hMK�ˌ����)��?�2�����rNp�Z�� [�:���/'��Q��i��4���fyV�r��Jdu���i���������$rGe�rL��ޔ|t�LOj�Ec�T��:N���q��3G���4Ϛ��n�5o��d��e�Ga��g jp�z%�Ԓ���E�<���0��.ǁc��i�#�|YZ�U�b�b��;������S�X�]���=�ܗ�q3�������V�������Ξ�:����d�<��/�;ɗ�s& q��m��a��u��Y�e����F_j���:^
K;	#<���>8���O��/�Y�ɳZ4륶�<�zǝLKmt-���Ӌ3��)�/���� |�F[𹍌ϲT���e_46�`��q(7<������6���*+<b��x�����qo�$*�T�GqYSC4煹��>J	� #v>�/�=Gy_���(����X��3mL�]��y�[{~�h�Z�v6����Z�2AB��ʖ[◼�{�����P=y�<�Z=e��g߷�u�TA���y�r����+��c&7���tZ���@����Y�ך|2��H����#d:����A�O�-מ�!��t�(��1e[���NȞ��i����1/C��j�^���� $3u�|�Q��5ք�R	�	55���-�mNT��{��2R��L�߃��zu��pB��1�%J~+���
�)��z�ܿ�-�k �AX`���EE �u��퍲^�A(�P��b|jSS��$��V3-�Vs��:��9�"x6a)��c����n�B�(	�<�Kw�����Љ3����nk�9/���h�Vh	:	�)�1�|m�=�?-�s�_�ZBt�l9~��K��5�閚����4�^Z8[㷊�`4�E�1�;�].p�?��$m�N��Nj�	�K�[Q(D���O��J��q��/�j���s���ǡ5�^M������Dj������CA��� \p�<�%�{���;���!�U���h=�ҙ$R0/��sk���A�V�S9>�Se{r՜ǘ���Osy�.�{٧��L�*jx�Y+we7�u�bGzN��^��9�M)'�pO�67?���:���sa�:�'�I����Y��T���������^�Q6,y�J���|��{ЄW����Ɓ�n�]����Z���ZRyԁP~s��Zլ��ɘ�b�:p�t�9�~�F���T��2|���ֳ�<�hLM��ut]��_[5�:ʺ��>���*_/�1���H��/,�����=�>4t�:K^?����_��^�T[�-Y�~
�vM�KK���_��,�7)�,�GiP��>�����l��ڸN��F�$���T��	�4�w��j���4�E�/{�gk�lk6)[�ԚC?�^�w5�|<�x�8��F��	�V?�+t:��;X�f��LW�J����Ro����D���6P��b.M�q���P�3�v���:���՞Wa*�YM]��M��>���+�K��Wd������}�QL7��0
_�����pb�eyC �g�`,�pTeFD��*�5�p������d�z���o���%����߼�*2�t=	�;��t=�]!f���k�7��e���:KxL��]m<�6�8X�5���G!M�;��e\�@��z�����]q�rH�o�q/���ۋ���N�/�Y��*z�������\8K�e̋ǥ^�O۾�)��,�?�k.=�{�J�s�l �����U�3Wc�,�ȕ�YSu f9�o��#e���>�5d�]�D�\�Z�+kh�����J�dC��׈�R�$��|�Q��<����h��M���#a3�0%e�'S�ƪ�x�B�eY�an��k?�{������*�+�oʼ{&ֻ���	�2�X��8EST`��6��V3d�8��;~V��Z�7|P�����#4
�$�sܪc�б]lrZBnu>.h0�J��f|��}J0��S�Ƿ�R�d�$O�K�,���7��1���u�q#�t}c��+K�g��sE��ぺ-��4�����;���H'���
�	�������T$Հ�g��&Ts���s���ɏ|>��0(�ZL;��NG-<%���ԭuC`I�� �BX*�AU��bI�c��~�赜�	]���㎖�V�����N|Қ��ł�N�R~�T�^��(\ӆ�
{)��T �bi�b�j��6#G��IU��t�%�b/ku���V;��N�s��$tk��}q�-k
��M�^�s����GX���&���q0%m���e]��b���aي�$R
��R{Fk��hA�D��rV��挕�*gZkbRf�
�7}+O��G"ɝ��kr�Eu��*�d��O���Ǧ���䪩��2����U��5Ψ@#�G��S������C�Mͩ��+����N�Sc[��Y��x`���qwۼԲ`24j%�0�o�\�&��.���K�i��1��5�G#�.�fX���K�}`��J�\���y�tӲ�4a"�ȿ��]��R��U�0/�c�\9i�O�]���1t�+�<ޥq(�8�Z�G�'�Q�s�g���o�Ncѥ�N5YO� 3'q���C�i��ze�Ui�˳����VP�l�`q� �&��~J��'�xiu{�qLc٦���;��m��V���o]��wF� Y�Oo�0k4�>fu:Q[��q�r�YO�ǿ��;�|-[�=��'u�0���Z���틃�1l��;�ͪ��Be�M�=k�`т�Ȋ���&}�
��s�l5�(��;`�:(Ue��1��N�ٜN}(\�z���O�l�N�)�I���j��
�\��=p������1p��gq�)�uT��`�X*.�"�'� ��I��ӹ�,�椘�*U6B�X��-��)e��x��3��FP��<�T�9�s� �%��b=����)\B�F���F6	�Hc�x<�s�)&\֬�AS�ʤ��ҧ�3Q��LȠFD#6��3''i�MK��0�x/-QP[�S�|-�쓙�h�x}�)���)���9�aJ@�)���R .Kh��gI���"��x�0zV�a9��!����J� ���1[���`W^�_2_� [�0bm6�r�&E7���2f(N�x�ȣ&�r��g����M�Z���(̔O���pI�Ie=���+��28��[�L�����!fw�2���p �X\��v�R�����{)������M�g�ץ'N�����1j�������H^�s��X���~9�gk�VT� 4���v*2��A��#1`�t��<��sY�~y=�oB���0��L�^Z��R'��1i�[�k|����s�ꦥ<��u_[��%�<��L?��'/�C��T3_&<�Q>Th�b9��#k������ws���!���t�"�sN�-a��ЦSYǔ,]���n��W������X�Y�)(|E����%���k�5�r�=�}�>W_�K��QHN�1	ߌ��U�l����,�����!�ħ�Y����Qpb��v��䜳���i�twuW�TuW�e�Y�3�����f�R�]���I�fT�&�1�&]ss0/�)I�̟���S��$_)%~R�����s�zڕ��erے�P������ʭ��7�[�3�h&Z���y'�W���5V�h��MCO�1wͼAL���$@�V�b�Gk��� �~���a®�����A�ywx*}�1��(4f�I�j�ۦ@����bDۊ.���>\��$��d�K�麞��1��*(��I�7��,'�6.�81s�A}t��Okd'w�����Z;C+�[�j6�q��=r���x�%�K篭��Nܯ�:&�1�"�/h���u"�t��Q�ӟ��r�2�x�� �i���0�ߛ�C���g�È�����C)7�1�9�.������^���^t��9��O�Ӟ����8P2�#/�%_IA�q��Q�̢:������P�۰+�KzAe�68�R(4���Y�AMp�.�h�� �����X�3�$X0m�_�1�kf�%���Ћ3L76��Sr*$�X�t�ϟ4�$J�.UE�H��Y�#��r�@���.q��{���Z|j�+�����M<-p<�cܯ�Ӛ���1��o�y-Ȼ��#��q�s'"�����h�n��7ꭍN7������PaYEq�J���\�H����2NX9���k�Pͯ 3�VY����8�E �WF�xC�w@8�lK�� �˦Wt��8�����X(�\*����s?;�S�[+ 1���V�-�*)�����v��uʈ�v[�Ĉ�m�;��a�kI&�I��}�~�7�k�'�1h���Y�����ڄf8��lƕP�j_�� 蘈%�P���Σ&�B*C*��Q^�|m��Z[K�O���e��1+�o�e�ڹ'h��[ڶ�>� ����3o�dKm/ZV�c���ֶS�;R_=�`��i��O6��妢c� ��w�7�N����B�7�^k6���QW�όs}M8{�g��v�`�lCݯ���<��o�z�q5����{�$e��c �<�_�R�.;OiS\�ח@j_iy��'�p��d����Cp�2k��j��6'v1�ך�n�o^���l,a��is��yi�����"�.���.�G�8���� ��ڦ
�زGh;[ƅ[s�-��/�רA��+u�?���25Zh�a���k���qu�"�O��X��e���G�~l�A��rH��+���Ze�6��d��u\�E!�����mD��������&�0��!��Z�K��Kp�6wz���,B(�*�Qf��E0D�w�И,8A�����e�O��-j���1�S
����4����9�r9�
ę�x~$E^][�y�u)=����`m5�ȷ����m�`'l�p�U�u�P��4���[ژ�6S�^���N��%����LM}��n���r�Ai=$�~�ǽǽ�^{�M�C����~�M`�� ���^DI}BYΩd^�p���*'S�P)�7㲱^����\#xC�80�	7������iL���)�)-WkS\��Z�c����S 3�n�+y���W~Z�iַ3�c�m����5�cZs�D�e诅WO��k�܋ގ
��*ի�Ӗ����.H�xi#y3�%υ��Ɯ�z@mFK��פ�3�KIl	k�]��9d�"3�9��i���5�_��O'tQ ;8�0�l��8�@Z:�W�!;$G�����\���[�/Rj}M�Xﵭ�ߔ^���.�{5} ��=�g����ڥ�X+�kMO��/\W�����������;�e}��oXΫ���~�qձK@e�3r��4��-�^p��p}��i����^���<���|�b>��ϒ���8\9�l삷��);���p��cxZ+��:��4���#�V$����W঺�.���`W�՗٣6�<c7��F
!�<]/h%�A�'#�|E[\�)R���A|hxze�D|C�S��r:�k/���r�=�������k���}s�h�h�k��맑͒���k��d;Һ59'�?��O��^o�/��0ߏ&�%+p~%����`iakK�^�O�.j{nU̡���Tѣ�Jk��aa�O!�pO����u*L|<���=h�27��)�j�NIN�F�j�r��Sa��?� /�.����P�Ȩ�Uc�PG��X�� ��h	��8G[*�����>�	
�XQ�8©�q�F��8#�Ew��ܑ5�U�A��z���*m����&�Ȓn{1��-��Əƀ��T�Is� _�)��Ǻ��!�2C����NkM��L0��5�[�%?n�-�m/�si̴�y[����|Djt)~I���QO���`]�@VU�^
2�<��e�k>^�Z�|A�2�ц��ߨ,ؘ`U����)]���r�(WF�疾j]ɡ�@
7���8�o�L�������X�;��m����E��6��8���
z�[���D��tP�W��@|�66�v32:�8�sC��X@�f&[�����3I��\�-�z�P~�G��)EAnk�K�7�<�W"�Q��:��m��8Ô%x/���I@,a[�P�A����̏�Me+�W��Om�:��2�n���8���B��B�2��MF(c�˽���j6eo��{���F_J���z��|����q������x��Klٺ���O�D�͵��[��XOcr�̖�~C�%��B�#|9�#��>	�.���O��&E"	ޠ�:�n���/���W�}Φ����
�R_KxTjc�z��Y�c������~�%#؍��Y��}n�nn�lD�`Tש%�8��������������
��pM=nj��<�+4�e�6��l��W��\�_�rQ�W5� 骞v�:-�����zд�U_R[�ޖ�f_H�5���pj��2�Q�,�4-�Nvtg�����'��Ey���@n[�����ñJ��e���;����j)&�ܨ�W+��?�2�����cHNr~���10f�l!@>�v�N�q���:j|�a|s:�r�)��{����{x�Ԩ0ƌ%������>��k�0�; �}��6���s��0��v�j0hFT�i��E���LC�W�u�^0ǲ�ʴ�)��D.�H�;��Y���V�7��5���Oi0��e�k-X�P$�<���LI��̍M�UXGi]����t���O*S`�[r�#�G��8N
'���~�}H�㞦�2���X.s���@qA�H|^s�ع>��YJ��)�.m�c�9��.����Me"ΠS�)�e/;�I�?���E�o.�5��u!�æv���2���e(�%C[Cܕq����2��l�)2��q쟢sI�����1%�9�4��,�jr������ў$O�����:V�'ݤ/��/*[kz%�?�[�5(0nq�G.�.�o����M �k�V���h��΢O���e�w�L�[6=\�7n�г�QV���`���$�Z�>��x�\�[��gǁ�M\g�����<O�k=�K x�����p��O0�������F�	g����58��;�~ !�8(Ò���|7�Ʌ�W�a<�b�ι�fpm҉A��p�g͎�mS���qje����Y��>�[�w'7�?_��]�k����$�J�5�G+sj��MY���N\[��By��_T_jׯ%��1H��DS�3�u	/IOa�P��i8�ǭc���h���r���r��F��N�7�� ��!��h#�l8��B<�ڹ��dCʄn�藌�^c�|�X��[��d�͜t�K^
�k_;=��(�H����w�M%��5~�q6u���:��C^뢍�;1��$�l_��%8pv#� x���8��#I~}��n��C�0���Aw��B��Ӷp���`�)�Q�(i���}�!q@2�j�0��q��DCC��,��]���v�8y��>j�D��zl_m�V��L�t^��^���l2�H��$�$ɍU�M���o]�f�;��6�0C}��ɇ�N$��8��BL� ܙ�	�X�6��	�8f���HHz�-�KK�N��.Փ�P�>��	�P�S�xՎ�[	(�y��b`�(�D:F�©��M��22��;�׌���~��pJ;L[ �ܸv�4>�}8#;�$?u��L
d ��$-Y���_����5Ɖj�
�����x�1�K�[��Z����\�p�O;ۭvT2w*3᧝6�l��ˁ&Ҏ�;���;�@w�_W^Ie\ѿ��L����K���->�[)@��I�\F�&�ߪ'�8�K�}o��`�֣XE�ްh-�5S����Qzb�թ����䗴���V�M�Kui����Jwma�,�qB�*.���{�G@��[�T����䀙��P�X/�u�t��I.�d�5����gk��O"��~����f����:'��6�˚�UC@F�7���]i������5�����.��Z���mj�m�?�d,�K�����m	�>�仄C�lf/�1�=Y��,��t~%���Z�L�#&�����������l�:V��ޚ�I��c4�T�$���c�q�eR�>³7i�F����Z���on��S��ub�O&����-�'*$9�����Q��h�=�w8�3�f:�I<�����jbR�V��l��L��d��o象(p���0H�g-��a�QJ���s�������U¿V����	h�Z y�%[��f:W�\�l�WM�K��ho�<p �#]�鵬W���[�|Ox�Hs�8�|�~���2$�e{.�����ɏ��$�KZ(���.�U�+��y)�hu��8��0����8ۈ����3d_�9� �����'54�K﫢@e���	0�1�R�x-賕r聩/n}h��<��-V�3�)�86w�#�}���X҇���ø��x�i��b�z�:�Z'_��K;��%���UONm��k�k���~jc�ʁ��g �נ-���1-�MI�.�{񐦟~>�A����=}��YRf�/�|4M;�e.8{p���f3pu7_�(Rl(��&'�o
{�+'�������Y]pͷkJ�8�3��k�^�cM �v��I6S��{�C��by�mj�X[��>ŧf�Q{�����Ǝ�lF�F"S�܏.�B�� �g8c_�Ӱ�q́�6�tr;=Ym����Ht�#�h�\-���͉.���G��i����5�q�x���V�ku�V'j�9ɶ�x��'�ץ��i�V̈�]��z��x��%ǸrZ=/�[���P�Y|Ϟ���ȓ�B�8��M�p�=�:�9��M�n�	\��R�:��'�cֆ��j��4ɞ�"6�?Ԯ�1��֩ىP��k��������;�6k�}�c��4{�z��Lh�7v�d!�~Kt`����և�NIzc�>���'�g8��8���Zh��эh|r���˷`M�]M�����k�z�Ƽ����.�s�)cӟL�>ҖЊ	jqm]�NŠ�X+�x���w� �W�+�E�:O��:��y��Ѐ�<�Sx�&Ķλ��A�5f=:֪_����y	����͇V��0��GDNǛ۹1K۪95��+dS��m����/g�7�h4�>_7r�o���@W���ߵ9^ھ�fm�5޺�-5�$ђ	e[9S�k�:T-×���:�c�_�8�I�8�I�.��}�sJ�ǥ���Z����G�|��0�1�OW|}G{���^���_�TlA_����[mo�㑠$���^~�������^}�����	״���֨��l[����S'<G�u�֋=�B���_�S�A|��Ex�WF��T������.1�o��dOj���L���^��I�r��}T��K��ru+}��gm��+Ŧ8���i��Z:���Yo�K���~�f^��g��,���Z��v��;M��^���_��[���m���j�W�����>ZF�k�X]�aҳ��v����I��.;[�T����%S��Ҙz�K���Z��m%Y�p��_�p�>�Gs�c�1�^�ǐ��t+�n\ۜ�ks��
x�{����977�y_�{[�Im;���զf,���V��^?A�SHt��-���V_K�s@�G�5e��v�q\�?(H����{xg	l㿕��MĻ8&S`�^z����{����0�{�Q���zZ��s$(k�FcLRTc��Ӭ�=�=���[2L0��*�"{.>��a�ol+t�p���4���Y�8�֝h��`�Q�]<>ǯ��/е����kկ�|k���b���N�	�R��{�7�#�������/���7�B����Z�L�_K��/N��6�Ǡ���ZG����L`q�nn,w�����ߜ�e_K�ك�����ˆ1���C��Ơ�ה��ȷ-d�$���G*��� �7���8�u p,A-� �r~(���U��ײ���=�D�_R.�1U',�%��lh>�!��0
�n��g��C�*�6�9�l��9G�-���.ь��:�}�����Nn�G��4����զ��ۂRkA�(~��hIp�T�kN˨�Ou��Y�Z�%s�KW����me��h�$��E�Ж�o.R��do�/\��c��;���<�%�j�&��x�N��0ux{N�K-�s��:�%�n��x�Q����R&��/Q�F�KyY[��������y���dg��l���Vo�����1��G�p홋G��9��_��Φ���	�i���������Բ�Q0��p���K���o�@=Bm���Q����R �ko%��1)�Õ�ϫ�S��q�kV38���#��fo����ڜU��m8��VtO�)Z���ƛ\ǟ�\�t�4}Q���8�^%�'ptG��jkY���U�1.�աr�S���[@�S=���tqsFq�r��s����n�٭`)-J|�A�pׂDk��J���y��k�{��){i�sD��'H��
6��f�x�.�B������#[���\,���H�0�]�^h�-�=��`��x���$�WlE+R;�4	���H��o�:�$Q�����?ඵ�~�B��=��V�u�����	:���^;I�ɗ����%�D������H�g�\�Z̄ù�_n��=I'I״ ɾ�ګ�Oˬ��j�x��8�{��mmA�kleZ7����{��I�:W�;����D[-��c)h��Q�V�5ͼn��9���P�O[`�h²_5��j_�,����􄳋I�����O���7�Q�X�ӌ����A���ѣan�|�����}�-�&�X��G�~���}t-�M�K��&�j>�F�Kk+�Z��&O���2>��[�m4�#�`�%���2���:hhr	d�ui��Z�u1e����FmK����qk�:��86R�+���;x5Gޱ(1���py���<uN��Q����SITwn�8I�� ��l�f�t�[J�ޘ9��8�a}�VFˈ���7��N3w�R�J���׋�fG�5���1-�ߣ�!���S~),�E�>X�V��V}�9�Z>����������F�z|`�iZ�Kw��+{�=y���k�fAk����?J�J2ZcS���M�]�&@�Eݲ�JRe+�����m��rGc�ln����]Rg���?�JW��ʽc�k��=��Z;k�-qފ��r���b���$ĕ�m����n�����Zڔ����m��>�<پϷ[+�j�Gs���G��u��C�I�#�0��N�i%2�q�B-Q��!]�R�/��[������ui~��5��\�D�P�K<���6hZ��&��&Ӆ�Z���q�/-M��/�S�
�9�2�s�F76�����ק8;�9W�����W�N��)͗�������?�g��l:�\�N^=�N8aP;%�Ⱦ?�	Z������͵u�.'<�<�w��	'�p�	'�A�ô�V?�I=�)�2�����9�-����^�v��$"��ٕY;t�o��|0���t~4	'�́���|i���g�D.�K����t�:#GP���|+�ҏO+y�w��l;/)���ߠc�	�'pD�:'�Yy��Ƕn�L]K@pe9�<�� ��i�3M�|ԭ6�Rs����쐭1Z����ɟ'�`{��X �1MF��2���Ŷ~ݴ�i�z�c���=���O�L�}��4 %��p�)�a_h���	'�B���qN��k']�����V���<���H��������~�1��Y��^~���լ�T�- �F�[z��{��^8��_�їsF���Ҷ��XF��lH���/9�A�s�����O���.���,�=qo��^)=�͟��ݜo�����������ó�vs�O�I�����
t�Bet�ޙ��4��!MG�0��m#��.�u`���8��9N���O���:�v0�A��	�ȣ�s����I6G���ѿ$#�� 0��)eޑ{n�ƃ�r�d�%	[�#�Z�k��~���O���OmN4s%�m��z�償p�(�<m{��K��	'j��8�{i=�w�	G�Sxآ��~ �L��C͖���[�2
�%< h=�:�<fA����7�mh�cM�'P�y:ߗ�����K���|ٽ�[S��ם���nsi��Ƅ�Ͳ%_�mH��l�Vb%��	��!��kIk�r�3���k�!���5	��>�ڄuM�p?p2d�S�}hd��I+���I�y��2�C�4�����9��BeǗ!,�u. ��ݷ�k@k� ��=��z<[BH�咓9N8�@3B�� Z%}�@?Ǖǐ'%,�I�Σ6�����l%>৶�d�Z;�Nx��ii�Fo?[��?p�RJ�	h�pO����n�o�(c)N[��=eH)�  �d����z�k�o��n��C�x�[��!��lҞ�Mި����ӆ,����������-<jml��4�����q�r���p�M�g��������o}��0�
���>��b�W4�}�G�K�A��'�,50[�pݟ�o����o齦��nGךzo�g��Ş����'\������~z_�2����q��+q]�q���w���X������&���R�L�Si�nX���J�I� �S��>���+�t-���
�52�G��Q���9����=��4�v<1<�\�PΞ.{q[}˷!�����s�?R�m��L;�y�5��f�;�~`�m�p���:5�u��s����j#GcwH8Hmj�?A-߽Q��~�s�%X��=aI�\�G��Hrg���&�<z=N�@ڛ8<��=�*����}؎�r�g�E��v^?A	�'rp��=P�������4�q,_�kk�k�i��W��a|7^}���7t�ϔmҷ�4�pB����	ԭ��[���p�k~�8c��O��/zL�}e�8w�k�y_�:��R���(��5���u�	 �q4��k���im�.�W�]�ZA۵�����w�2'��h����*�O��N	ӵ��z[W��gO=��&�'t�i�Ʊ��9���=P�Zƹ�j>��95FGY���c�Șާ�_�����'|�^�Z�uK\�m�VAڨk�8��^��r4|ƽ�=�-�\۽�Ѣ��V�����V�~��A���N8�5���J �ʪ���i�� �j~���%p�n������z�E�Tq���Q�;�` k^+�z�}B�l`����	�p�@;�`��;���T�b��ǆ�2�s*j�۠��,���iܲ�g͓Β�P����_����1�ih��&�>��%�d���*�����A�=�p��8!�	�En��Pӷ�f[B��z����`�V���m%cZ:n��W�`�H�7s��iߊ/��1����������~���Sx��8�	c�/H'�f�lo��֠�7j|%��-ݮ��[���mw�=�i�C���]���߷����k���=�G%K�I'�p��O��N��r게��6�5�b�K��6����_�W׮�4,$p�?�6-��-���R�D��[m�K�8��g���x<vl\2��]x���'}�zG�i��k勥��c>^���^[:_{:�v���.��1�5}���Z��^Ox,�8���7��3�ޚ�JE,i�ȶ5�F_�&��68�O�
����樰O@u=H��o��5	k��G�0�u�[%��Y���k�>�(�%�׾æ"��֞� �δ'`|��!�N �%S�f?s�ȭ�C  ���l�O�� ���L�]	��-��	<��Gu�/�(P��:_�b|�n3�%L�N���n�%�k``���C�{M�-f����9
��5h�X����:��ex�l�ΰ��1�9�� m���Ǳ���_�7>jN�L��mḝ2~_X�Fkև^{�9�hO�4�8�ج=�������(�<��j�m���5m�i��R�.>������k��;�@_QK?9���-��Ƣ�尽���a�ľ�6�^K����y����V�z��	� �����e���1y.κ��m�=G��8FB�	'�6��0ч*����O(�Miޓ�1%o/�uF�]Jc��%)˒���ާԃ���|�P|n83Kh��N��@e�=3ǥQ��NM[������f,�����z�&�O=p�ۆ�o�D�j������~d|��A�G�}����u8�9����\�ț^;����^�/�d�@��:Z:e�>���=��\׷�=vl>M��p���q�z���eq�=}l�������	'�o3~����־Q�ʇe[��w�qvt��_�b�kK�D��L;}��u�Zc]�T>R;���{�~���~�ݧ�l��V�=a��B~�k����6�3X�GB!=�:��1��'`~����m�G��6�j�i �B�I��=�0��i(p!��c�}�Zж� hOC[e�p�X,�w��`��H��kޞ�t�~��v*;��_I��v�e5�jV�d�s:�`�8����vR�G�Xx��.��lc�����֑���a��s�>ZA3��.���7���o�񔿗��D��vά���ܤ��ߛ�C�:����9�Z���C'��!vZ�|�֖PK�h�5�ӛA}��A�ϒ�G]�Nx.�����ƽ�wQ�4�$�}�E�d�	��0n`4HI֖�Կx]��I�OF�f�p��R �S�K��i�B*C7@{�ފ�s����6z���� G�y�$�'h�,�έǣ/~u�2�*���]*�j��V��@���'wk8��.M��IL�%�i�W'���?1��(��׫=>x��='�4I@ �O8aX�W@�h�<��O�s:''q�yGko�~�}I�9��^�B���xL�t���}����x�0�����ײ�k6,ז��!l-�Z>���ka�Ds�c߼�W�n���5#��~��DG��x�G���Y��IS'l�cp=מ���i�)���ϸ8�֊��p�	K��>m�cC�Xk���
	��^�n�}�JU�;���9S���?a�Fs���Y6#c�t�)��t@[��)o�AԴ׫ܹ��je[eZ}q�g-�C�d}8np������G��9��iX�`�`I���.%:pma����o%QH�p}��,��p=�փq�@�����3����K��*��p�	'���H��/�&�w.�p�ｬ%�d�:nP�ۣck~.3�?����CH�>�?�S�a x,��H�kk�ʦ�2�7�}	<�,Ё�_yYR[�5񮚟T���I(w�^N��K��&}u�#����^���(H��� [�7^�N8�1`;��pB@F�r���g4��Sm�+�ct��]C�{zj��A�y�����1���&��4����Z��HM?= %L�ع ��N�%{
����q-S�N،��C�k�U��&3ڭ%S���k�U���]��G0^�yl%^hA���Z��%�r���B���I�'l���M���z�7�k�$�Z�מ6)��ף4z��A�^���������V��Ɔu���y�/�� �̷5��eZ�w\�Y/,�ϼЎ�G�Ҥ����d�/��V�����
�c����e9��m@�����8��h@e��2\��=���� ���O'�p�	��i�߽��mە�q�h�ˇ���O�c�[�A���D����p�@�S�J��j�g2��5����V��z��4��M�����	��;�,��M�7߈���\Π��5��(oZd��gn�m��穟[8�2�54'��n�h�d\_�ce �%�������G>���Vk>�󊟤�@�No
�|h�v�rMrI/-.I�i�摠5��x 8����Ǐ�5�{�C�Q��$�MǄ�K6g�}<��IZ������{z*T�7�,����n��2���֘�[�'-��F�=z�-`�Z������s;�5��;��I�1�+��'ؗ����kڐ��s{|m�S���In.�{�L�ZyZ����CQ��Z�vީ/��]����ŭ��ڽ5��(v���<Ak�P�f��7ċ[��g��h]�'�]�/���#A�sz���e���>8��2��Q�wp�s�	'�p�	����� 7�e���&U�ۗ�q��cx�e�ݾ��F�=��c��!�6Щ	�K8p��G����2D9g���r�7-#�]+S�-����E��4jG#&�&Z.��c���d	\���q� (.�?�Xu�Gc�{�_ ���y�E�PF��9r�輷LK�M׵�A�?t�����E��:��B�7׷���B�Z��8��kA��i���@1��33%Z�~���Z�#�Z��8j|���C;� h�G5Q�֑�\)�I�wI�b����@|�&�k|Ǖ��o�(�Q[;�������K���Փ�~	5;F�c@y��^=9]�����%c�B�^��6�ۑO�̱��d���=�^&>l���~#���L� 髚���s�5e8��µ��(�x������;G����e4�8��+Ásx=���˷�_Gs��g�ܦ�2ŗP�j���vt;��--8���Z@Z��p�C��ke��i���re�I-Ň�VwJ�9|[c}+�v�N8�N8a�7�A���1쩆�
z8��� xS�S滏���J�	XIs�5��)>���Ɓ��i������F���t�j���O3'�}O�፸mnˀYᚭ�q��εE� )�*��o����pZ���𘹯V��X6p����v\���M5����\N���`�0�2�&�Zr�セt��IH�Sܹ1H�A
$SY*Ak�y�r9G��3�:����=-��?�9�կ�.Ƨ�omޖ@+x�E{CMOe�L��H<FaI�]j��o�fkx�����@�ԯ��� ���Y�]�o)��ڞ�M��'�[��C��߭���.=�Z�+柣@k��=<ǰfj�G�t����8%����ƾ��l��^.����G�? �����|�^���5;	��%#��z�Ɏ�cÿ5�~��e?Z�ںW�7$ڧ�S݆q���S�u4�ןt�]kC�������[�.��I�7a/��W��k�Wn��]h����M��]qmJ6l����8�xp)����Q���[;7K�B��$�]�q���g'��%}�L��Ҏ�N8�Y@���A&{�oG�|�	��0�W��M��V�t�up!�Qt�WX�Zθ�g��=��c�1����-O7A�25]k�O�$gTr�blΩ.�ş����EfI�r�wR���Z��y08Lu~�K|Z|׃&�G��J��-��y����c	7�L���7X�
ʵFmY)��j����1����2f�|���~����j��V���4�,g����4~i��y��rc�e9�L3w����)���c��Z{�G
TQ�[F5wC�G0�S<z�K���Z��~%~��Lj���vj�O����{�\hٰ�vjx��Z�p�%]����4�5}��K��;G��5���[�[���+[�|Mk���=�]�-A���|�>|���}��{'�3�f�D�5��婚LY�S 5[�Zu�"� �O!�Y:��!��\{�S��ku)Osxq�Wk[p�j�G�k�	.'�u5<k4�音9�n����~�kn���kl�}�, ��Z��Շ���w���������c5?�&�����u�ַ�Z�ңӎ ��<�^H6�����oE��ݚ}4����*���
���7�1�:]ta�8X�Ղ��c8�qIY�t��I�qe��Z���O�6�Ys����C�J��C�Yc�	'�s�<鹘.��㾨S�jg����ѵTO�a����C�95C��r�ʆ��_)�����9�@�n�d�<�s���9ے��@^�N%y ���L�_  ��k�6�'���T�����K�^�Y�x�[�A�Ӻ�)�&���r�Z�4:D
�I6OOqz��g�8k<�K��^��Q�T�J���C�K��d�$k�5'Bh ֎�\˳G��-+ի��V����v[�y+;�f7��������E�̢�.�ts��\{?p�t2�1����5��с�m�c�J��d�VϾ&�5����9��B(���������ڶj�� �c��S��5z�hZ�19�fI�R�)ΰ����s�p�8ۑ�ks�(���~YB�k���{�+K�F�r6���S����p�/������ύ�+���]+���q<�X�}ݶ�	'��va���<�� ��N9S���8��f	.��t�&ӎ�;��faj�Ulk��^�ϲ^O�5�V2h%#�����q�x玅�˽ArVt�7n��� |j�4�i�-��{R�ו�6�]�ɡu8���&pAy�Ə[��͚<�8����V�-U���1QѬ�$�;�8�'�sx��o��-�:I�εרps����׺L�T�9��x����\.�"���)��_sA�Z�VY�����űV���m�v�k��E	?�ǫOI�I;U��T��{�շT�pmK���If��k�-��s��X���
��59���]F}�{�[�]�ߥ��IF��#��P�W�W�������vZ�Ji��y$��i9]вj�ƍ��h��/���$%u���i�ïE_[�_=��.�$�����kuh�-R���<	���s�5Ζh�aRے��&��J�)��?������j�K���v�k5zʷ��)ߢ/\�J���R���1>�25����&�'�c��ՌS�Ai�����[���a��ANXZ�w�	'��`K�'�>R�E�Z�2#,\q8�a~��\�/o�nѴ�:8r�U��8!� i�?�qj�g-���q�9.�Mm���=Έ�]��� ��u�E�!�l���6�Gn�kA��5
�i��~sG�FAv���5�
8�n�C?���|s�jx[3�6�!�!��@-p,��~[t����!�z�kZ���m��^���s^�=�I��ƌ��������;�{��ũG.�	�z�{=��(=���:�轧���(O͝��,WFcj�LP�Y�M�V��X%\�����Z?�2����ւ�5~�ַ�#�FOM��z�	j�@k�׷Z�	]��r���qi]�,[���Hr��������~M�h�m�p��6�z��9�C˵��ؼ����뵳q� �>�؛�f��Hx��%�������^����EcKׇ���wM���{O�����Z��*+}��J\�^�i�{�m���q�h�a�/�=Q�Y�ť��[�3����X<�NxM�����-�ЀZ֕���f�S�ϗ*��W|���q+7�?�Q���P�x��`'��`����{���7
t�$aX�@�1B��6��� iy�����*���)3� ��bn\�������i�Ñ~�P��-�GS�n�P~��$0*�j2b����
\I���).@S���y�Z+��e���@���Q:�}�plɚ��d�jr��|MCC����'�5���o�8�>$]��o$[����X��? nK섭��?����qlM5~�ϥ����y��j�=-���]*��dY�����w������(Ku��[�}��i���bmS�
7���> �|�%�Ҷ��Z���m��5�A�Z����r�O���M�_��R=<�۶���js���%:����*�"���\�k�mN�n�'�Z�K2_�����ԗ���ܜ�do�N������ ���q�v[�ˮ���Z�֚i���y�Gm	N�q�I�Z���K�]Oitb�\?�q��>�Nx6�R�m��h�o�~�I��cp��o��lg��"�M��V��í1���;=���$}O�la�k�3(9��wb���ɨ���񽇁@qYT�9�'l� ��:��ۃ[;��8��G5��Xzv�\�\J�'͚pץ��TVz��[�{�N)�X���f��A����ϰ�&�&��^�-�ֆ�}nG��r�n�r:`�|p��=A̖�H����X��г���)8M�e=�3=��>�A�F������ْ��%}��ڽ�F��4."�$�[��'$ZS��#���x�:�^l����f�s1�G����v���5��J	 �/��S+��^�Z������U.领G�7k:��.�wƠN8�N8�q�Ԇ��>H�sſ	;��.��x+{�5�M���@�́���l7��fd|a�M�A�Fx)�hMX����q�W�H���S-"�?"�y�X0��Q�]k����<˺�8:����Z0���VN���6�h���S���:�G͆�$�[��m�S9_kG[�-�=��5�lɃ{:�>� ���z��̒`�xK�ε�y�Y7t��	���[ٗ��)۱��P�T�o!�8;�YV�~CoUO�ؼKd~�����c-<z��lt�Z2�g�G��U�HpO{�?z�q@���I������0�rI[Ak�C�f��{���B�ǯ�H���R̗;�+����x�r����{�t{��F��x�%4�Bk��p�	'�p�	����-�.p��������:��9�6�'pL���\>}��G��!}��w���]&$��	�&L�����E�ʬu�7nm�&�WfTqF�#��3}��a��)_�ѣ���֭]{��&(A����o�u�@�	ǅ��w$ݺ�N8a�s�=p:�(��fK:��A���r���s�GZɾ�̖������ti�{�kO�|U �i�����ŧN+AJ�:�<q�9WK��\����)i��eG�9���c@�4Hu^'�/�%��zkpޚV�|l���_k���\K���,���ecp��C�ͼ���qI;K�?M_5�[ ٪oZ�����x����E����ۃ�&�u�߿�}~Zk_������|����������:B���1 �2)��~@��������F���E\���PKk�sK���oXP�$�U����7,$F2�� �B�\�
�Y�%��ne�r��K�o	�����]?�k9��.\�����>�c���p��'�F�K^��Ѹ����^��}4��|/�Ђ6��Tx}��
K����q�ܣ�SG��kX�������e�1��6|z��6�'�����8�\�����aߠ�Xj��6�4�׀��%��N��T��:���?H�����i}�.�i����^��v�zM�[���M�}<g��O�/�~�zH�i;�_�:���x�:m�^�c��Btl�������矛��8�ڑʴ�P3.\N����������P�5_K奄������'ƙ�m?]�y�(3]�'ԝh7��0���~_?{�g?��'��>��ԕ���|���G���F{�g�^�Q�덉�ѧh�i��a�@�4P�?5͓�w�$���>+�˽u����ѡ�7j�mo�����_z�~O�g����:,{�i���
�O�l�Fo�����]?�k9�����'h�s}]ZR�gp�&(S��[�9E��90�׉�X&�_3�lWm�F���"�O_�g��w_XX��i>=��^��-ǝ^P��_����r�x��T7��J�sޖƄ��s�����Q �U��	��l\��ߵ�k6#i}.	aM���V������iN1�R"m�����HZ�V{�\�nh�-��%N�6�9z�h�Bh9J��8(I���L����$��UW�y���G/�6��yR����hӄ\�����Ң��9n͏W�>������ί�|�OR�8>����ޟ�җ~s���7?|�}�r�8n����u4��7l�,���j�����r���pD��~���C�	{z���Z�p�d��mf�2����ܬ�	'� ���N:�G@���½S'�����Ј�	���	���[�>�	��ZܓnE�t��+O8�- �'�p�|��U�6��%�����k6��&���h�[�j�@��w)1��<����p	=�n,K}a��c�i�4Vn\�R;��f���=%D��}q��5�$���d�#��Q��S�������=���enc����t��������|�_������V��5�8޿�{?��?�k������;��;�|����M1}����1���妬nH��sҺ�Θڙ1t��i��G3��{fo=z>����S+�J���d-�~hM7.�i�J�Mr|k&��^Y%���'�9��6�nZ�ڼ/���25���ԁ�f�G��^���)���ӧX
����H�U�=?Zȉ��oj�Y�L� ��W�������c�{D_���S�ϵ~No;m8׵��5�?�kV�������mm,�A>~�e�e����x�����p4��j~�����3����h�x,�����pD��6	�\㞶�';��n�-'���m<�'+�8���2鳖����v�,}�M+� ʄk����4�iO�h�9�����7šLd�s�m��G������������O�Ю�=_�������C�n�(Oi۹�l��b�p2������$.�c���㏮����{?��/��		�`�8n��+?����~������?��������)�x���].�ϫ�7\���*)� lk/��8N_h7H��z�1�ӈ������ ��  ���$��c)A��v2���hj9��"��_Kh���\�=X�zW��8W3��'mt��r����?oiίs�:vZU^���帠[�pJWb=e>6 ���Rfe���F$��p�W���9O�2�+�!��IGYa��c[/�m�{,����)�,��]���N@.ߒ����SP�ف�qq	��v��/��O'F�%��)V\f�����ˤma=���'y�N_q�?m��w�X�g�^�O���L>2�e�0�T�O��nl-[�G�ruk����qˍ�zg��S�����6��z�!5�Zǹj��Qߵ�)[�V<ޜ��h�����W�պ����ٕ�v$9�H�S�a��yp�݆}Ϡ��M9ɿ����W�4�p`�2~V��_���l�bB����vNhC���	�}@����'q�㧬�^�<ҟ�Fbؽ�׭���68������s��X���d�	���k�M��.����5��s�D�S�����6�7�m�9�lَk�.������]2߷��Ԯ�S҇��5�d��e��9�jJT�|0]�8Eޫ�d4^������@n�G�(����:y�.�'%Hii/�\
�N"�dh/>s�����������3$�̾Jޗ*�`�Oe@��)�F���h�c�G�o��/���~��|�?4acT�����߿�'?��?���������O?����?��}�>fgLL0��[8�+U�������a���VD��$(U3|��Ȕy$P���3m%�l���1��M[te������r�y~��^��u�QKWt�}�nq�FE���Y���q �<�6�4uӧ���_ԉC�4�� �(3`�aOw����2�j$ܽ��8[�)���dQ���7P/r��g��+R�͸_���i�4���� �d�����|�:��90+��\�������33�ވ�g:�i�-d���oɆ�ẫ�,���]��������mK�\�����6���-��r�+m&��,�g�Gӥ�`�8g�Xc��4l�Dw��іC� To�F���t���Mq�;��T+�{���דdU���BJrx+`�'BìmQ�mY�e�F7c�5�d��N��^A�a٭�B�iy���,T�̱��5�UV�iL��3Hvuya|�}���g�k�l�+%:u��[�C}��4���K��'�<���zY�8a��:l%vZO3�m;lй��ʛv���?�{��=1�0N=�����M�sm�u�2%��M{\��su�䀲��\H'��18Fs�R`���㱆qpc��`ge(�x��'���u��j�	'���?�qyl
|r2�e�$�@;�$�y�O�7��7i�yO���R��р�&s-ˍ�X��f4��������z�h'�L����]J>�߯��{y���k����/|��_��?���G�ok��	����w��+����������}�~��q}��駷�޹a�]��OԈ����46gey�sh�;nu���F�*Z�����.X� )�RQ��i�݄���PV��y���q�r2��p�B?-�N��5[�C���ƭ��91g��z�un0l���Ycŀ�\qjnρ�-f�,�g�s8�՛����1?Ѡ:��?�/�����m�W�pu;�]�涹�Mt:�����g5�,���|>G7�cy��sֹ�eވ^�N�iey��m6F4�1R.��<gvmw��[%�<����iR�N��S8���2�Q&#jN?�s�o��G��Ò�Zf�YE���W�B6��pA�E]1}6�r[c�8Y"c�BƍGH�Z ��X3.��/ÒP��O�L�i��9���[@�*�RU��Д�F��5"=�t�@�~f�Y��dls��'���j�|,�e-7�������S���&����̏79�m��.�4�;��P�(� 6�ӓ&���2V���r��O�S��wǶ��4�Ě��*~�'���Bz��{`Yߪ�6Z�meνt���4_^RO��ř�1��W�2�Kb!a�ج+@|�G'���=r�Ac#g��Y"�|�?X��ħG��dFJw�'O��:.�u�$oɜ-IZK2��;fq�8�њ�<d�J��F�N�5����^h*�Ľ����Ie��EaӺ�hx$N��{M[��gZ�5]M�x�\�r��aφ����$�18�cJ�xyy�O����t:�?�o��_�s?���έ��F�$����������������������?9�>�����$(ܤ���\|��u#r�@��0	����B���X)�;"c��1�	x'c��읡���஛�eχ�1-���֮��H�䨵�2�	�2h�8i�l�\�礪HC�[=��A0+%��G���)�-u��<0�e�3o�f����%-�=�"5Wr~�`�b�39���ĭ`)~�zG�[m��xF!��u_̤��8-��l�6P_Q�v�_>�*$�O0"=	� ijo���1G7�%�So�m،0�[%*� ���@+��-���ZOX�?�u��m\{��<8]*ش���eY8�pDefͺ̣6_�u��"�i�myۻ
�a��fp�;�R�W#yyũP�M!��	A{�=��6�᥶cq%Zvi��1hp-�焉�@mx(H#��!%��!.�8;���ʠ�ޜQl[��k���o�Ξf�#��M��lL:2�lv|��A�b]�xM}�č�t�6^�>���O_ܔ`u��b������+��O~��~�o}����3!�
K8��r�ݟ��?�?���\���������/����O?|�xB�!������$����ܴ�t4G�ԙ�hH���8�,���M1����6 k���%C�,����b��qQ!_n3a�Ȩ�c;� �p��>BZ�c�ZT���2��1>�X��<����z;[A��s#�>��b�8������I@���E����q4�A���b`�4M���C�^�:E�c��ر�@9��YZ)5�R۵'��=�5tB	��êu��3*�\���z,�^�概\�����X���U���1G��TgVO2��)��*?֭t
����W��k}re�?�&O���ڃ"Uu����8
t�qog/�F�-]��sM��n�\�b�0�s�O��e�6���S�]�a�၄��S��5r#z-���ӡJLW��$g�>_�(T��|_��b��w�NI�<-Z���s�k�;��>4�i��(W�Rv;�t��	݆,��E*c�3�6|�I���t�L~ȥ�7cC�k/��`�487q�t���w6Ln^��2-��/D3B;>L+*�%=���1�j�3-3Ӊ��j|2G�q%hh�?��~)����%�f;�>�žt7A��U�����@�c�n᧕yG�7���ʚqI�}E�-�`��J}'6�ߠ�����K��8��dL�����LE�����F����0m�ݥ��;����/!V�}$�����u�[G�B!z��w�o�K�&��l�QsB���'��U"�����i8��?�qP3�=���{��%��4cy��UfH4<�� �I�p���s� W��7��I�'�2���y�>M89�&bS�_�՝�Nn�:�����ş��n�ˇ�?}�v��_���~����_��?����[�f�˒��0���?����W����������������o~�o���O>��ˇw7��A=���W�2����8>�ez�J\��u���1(�>�E10t�	$~��IqSo��x��`&F�1'�9]\�aHZ�ߙ��ތԏ,~3B?y�����&��B򕳙��O6�w�����CDǁ�i~����.:߹(_��-Ɣ_���Ku �i�>�`�q�!/%��uE�#v!;�&#��0���/3���x|p��A��!̐��4�pN���y�0H���� ��>/h���Mxxa2`��J_�ż�Zg�\�D�3���0�/��q~Q��%�A�t�*�+�k<�(�	�G�6΃���@i�Z�N����0ħ{`�&;a����`7����a[����<=$޷i��5 ��I?��1ř}q��v�r��qK�n�.�8O���yq���~�L�DE�/�v@�:«�\���]"P�v"م:����s�Ot��9�KoњM|��� "0��Qpi��'���q|yM�R^�ژ�(MeM+�Lj�7�$�ϛ�H4��5�'\K�
��c���'y�d��@�(�*,��l^�r@>���B��8��>���3����]�G�M�H�/	�D�X�A��,�La�dY	��겈=����s������6-1_Pa<���G�]�"�G<��/,�[���s����2��uH���3+멒�`�ʱb>��D�c�-���K/b����>
�Y��13�E��!4V\�G�4_{�i��2f�L2�ź��Bg��O��]6{��<�6x��R{���sz���Dx"F�A���*�hIweYI�[)h')�p/���`�N�3����DyM��%ie�/Hf��1Y��ӮP��V.[JY�d]��,�ݙ��$���1��G���v�i����o��-�I�g��o3{��%&Ð�^/*�dg�gL�uIAf����lk{ATʼX&�m�k�`�@���h܋�Pn�*}�_@'��j�e����l��@}�(׋� Xʨ�.�f3���2,lj������C��r=b=;0���#�%��ք���׈h� L,ȣ�ȡ�&�*C�&e���dY��l�+�Qq=��-�%��
�^���8`�㕄��:��b:��u�1:d�&_�
�mR�~��N���_��1m# �����B?�}D:�G�":�dC�΀�\Ksh2�Pyfl��h����+�b)3�2�n������I���a�<�@�	�~��e�d}�es�*�}�ۙO�m����3��d��\Z���-�<�$��ۨۑl�A
�� �R��:5�?&Ȫ��r�n�6۰`O}���� ���}�0�i�
c4�Ҍ��5<Or��!�� ����e��f:9�E�6�Tǌ��i��tӱf�)�P�h�l9�H�/�:˿l+�$�퐥e�3}[�d?���-�uB�S��%�h�E�s|=΁M(�5s�NR�y�
���_���m���t�2$^(b��ظ8,�_ҢEv�=��p\�ל�w,�V���v~�X~��ƺR~bM����ċ �C\������3�.� �6n��k�H�p�;�A�@>��F�੨��L���uż��v~���Э�T)1_��|�W�ܬ�q�>%?�bPE}�r*Xi���0���5�%�f�[�0�"%�Oװ��]�z���6��n^��3���ئ��+oY�\c��2>X�O�]�>]:��ە^[�����G�8Ze!V�l��q�����WN��-۳Ky��E���Q�ټi}��@ijc �_g�v�-t�M}F�@8Ov�t�:��^���~�`����˷۷�������_����7?��_���:�ni�׻w�~�G��~�O|�K�������S���������k��^��8��ٯ�����:�Le��=���{>�x�e|I,Hi��2�|�U�(*m�[��	�H^�#��^c�l��8�Ș����8&/2Q>��/Z�?a	46(���!����`��C��0�⮱%h��)'ݜL�m�%9[r���=�(���9�{�$��H��ysrL�����i���@��%*m�0���|�5���&�|MT�?�����$㲃?����f"�t�
s3-c�#^H�~���/�0I��q ���oƔ�	�-)8尌���'���	6��k c;���%ȇ��W.��:}����L�>J�0Ƥ�}Ҧ�`P>���=2��&����t6&��
�ߗ��eB6�_\
6�?��̙H�6��%;}%��~�����f-G����\5��r5�눑v�$e��)����uŚy����c��6��d�:%�
�e�y���3b�,�&��u����e���\\��l~Jx1��,S �<�b��T&�)l(߮}��WC0)B�C� ��f�2C��<���,������Я������M���U�7�Q�=��5<�.ѥ%2t�л9 ��˓��Y/ ��q� ���Q~��-"f���IW6q~�+l��@Ol���Ŝ�5md��]�����uP�W�vh�Q�]�h��1E���v9.<ԑ��͉ �y�{�h�]�����	��Ф�Fh;H�+�\�w�B���McthC�S��M:	p��7�ە�k�f�ڃݐ�K�,�|k_���t�'#!E��!�[hK:=*�ڸFt��SAwPecad����З��/hb���A�7�b?��j͙	!�ڇ�I�FY;��m�v�M ���/��~��5cӄ�u:�0�$��w���xM� р�����!�6(H�̛֤�c[�yISWX����N���k6�kz7��0bQb 8|E�1�_�ǡԘ�E��ű%��^g����;S�
�L��Řlo�둇p��N68���j+���1�$4t�ȟ�F��m�#�r����Dd]�"��WBs�U�3��I���H���3�z}�m1��2�&|��΀5P؎�����"�>ݿ����z�$�K��ؿ��?�0��9V�]q��Fh�ܘ�:��KT4�w��i�N���_�7�K:�:���eA�gk�m|��7���B2Q�#�=�U�K� 	�\d����'��^�IT�aeE��5����n�tT��I��yk��\�B;d 7�>��J�h[y�u�hƹ����j/1�!�ʱl�e
��E��D*�L���Z�+��:ˀ�f���L;�ˢ�§���1���^�9s���(/�������!o���� ̛��R,)���crI��� 7�It�Z�⤪P'���~zH�=�/C��>`��_Mq/vP{�f�ˡlZ$�lJ=�dT"�R�k�H�ht�R_�Pj(�����L�j37b�8�*�k3�c�F6��q�(�	yQ�X����| �E�?4ZG���gD���]��" �ќ���os2u+������S�$m|�<(�m��#�Q��&�E|>F���-���҇���$��e����5�!��\��)���C2�Q��m�;ʱ!f4�+q��a�z����{�6]�7�a.e�k٘G�(b�ڗA`*�L�`G��:4�ȱ��בC����+�%e�Kp�^�Q&�8���n.��۞�}0x�����g#pe˖f�{�-�n�G��7
�p�\���vZ�H���h̒_m|ֽ�Ljߒ�Vy�~O�v�+񙫴Z�I����쮱��JyV��;��J�#`k�;��i���-����gM"�ް�|ͫ���3�k.��]L���l����{�MB�Xהj/�>)��8����z���޾ç}�3��3?�3��������}����⭯a�$�&�c��0������������O��O����w����_��/������������������������}1^=�����+�i�C�6� ����{P������6M�	js�v��t58ڷ	����������8ɸ��+���Aj�ϫ�Z�1�+���$&�9.`�y�o��"om�oc���͝=����D(�����:�V_h��q�`�6(r� 1#�w�9��M���.S9<�3k!���	vIV[�8#�C����U.q���=�?�+���M'���tm�װ[lpH2e-��`P����9�'}���0#�3p���*S[�9<7�ΐ��4���S%c\;x��b/�lX_<W0G�������y�b����~v��!p
����ʌ�q��E���3��x����^��8�r�#>6����	z
|�+�\tz�im��N&D�C�C?��7C4�'�����̓#���6�\!ԧqO��r�s�A�(�0q��-K�f`҅���|���C?�Y^tQ�e�d��?/���h�����_�%B]�|��ߔG
*q6>�#�������2�G?�ա���B�pV�����o��t�����W�l���`�G�l�����)щ̓E�Ԓ-y\�#�%��Rզ�J�#j�ŶF�#`�%�� �8:�0�]9�,�̜N���'z�?Յ1������Ah9\ߢy������͘�P�L:�+ǊP�3�I����5�.�'�3Ź���aS;�:^'B��	�w�\Kl�ҹ�h�9�kh��5�e�w�+̃���8QD�����=�),P4E|�q���8:���ɸ|���p4,�U�!\�tnҜ��:��� �D���Y�7�)2��~��]G�N�PC�)*z�}�Ⱥ��Fc�v`.��t��2Zx�3�MoY�t��<i���x��f��P��OĽX�o�FI���)���Tf��ºL��6:Y.$�N(�z�^ڨq�!|�Zr�|\�S_4IN��^�����&�/̭�Ȟ�4w ���%;�%�ˤ5�
q^�qZ;l����,<͟��d;}�U�ok
S���m��"i~Op�&�G|�*�Q�CO���k���S�^�F���u�����N)��iv*?�Q�� �����qUm0��h'�9)
?����>����y��\�Mz�k�qH��@��%6[)�x�Os<���$Cd4iw5V�2o�������Ql�`���)6���x��O��τ	���%��}�KN��r,Y˴Q���T&U��P	�0������ӯx�K]���_��L�~F�QO(1�B�q��Y�ڸǖ�q��9m�&�@ײ��C��(�o�r�.�Τ.�±)�.ˍR�ey�i����%Ρly���ۺpa\g��l���{��~>���_NFFB5�J��i)A�L�`�B�IF�i%ӥ��c����	-#��D.Q撓î��6��D�����_CFA�_��dr4��������N��|,O��X[���A�0Z������]c��9�4��i<�t�Q��N8���$<L�U�@�E�bFnE��招�8f�~����Q��zy
뉗#ň\�!:���D��m��
4^W�1Y�3�?Z��ksׂ�A��tZ��G ����xo*C� f���eʔMv�%J��"����L���8\�5Q�&�z�:yV�S^~b�!ħ!u9��a�S�6���d۩�+_ҚB�Ks~�1�9>��Ok\#��s�f4��{���X��%CN$O�����s>U!ŚS@<�z���Bi� ��2a�c����>���1>���'��=c���B`�4�q�6&��h���f�^~�7~�aZ�myE�+ဨӐ{�5��~X�>�[�_�<��}CYg�rUZ��<��<�n�Ʃ6����#�Osp�Wo�`����yh�����Iq�6��ܬ�شn�>fE��ΌA�{�Y�lm�E"�I�1�J|Z��m�����Oh�;3�S�I�m��5�����u9To_ɾ��|d��v+�}.��0��t����m���q����)/���
-�"�a�%R����jn�����������>��?�/��?�?����/��?���˷~��ҭ��M�M��O#_���+_��o��������}�~��_���������̇�|���0�����͚���8�1�/������V�W7�E�<�b�Lr�Ќ����L��� �HK4䀃����x$���At��G';@.)}����åD��ɖ�IAo]��D� ���Fc�
8x&��qD��8��bR���j2�eg��d2"����S}'��E\6�� 0���9�Ƥ�)�̃(�V�)�Y� �l��y��;da��kF�
O?�N�z��M�EE��3�
8�9�5�]�3�갹_8	xy�"ʡ��Dc>\�$x���S)@D�#n��� <O�it0�8�<� � PD�fۨ!l�I��<�9�Ĉt�H���W��j�ŀ|�Isl�)A�@;R�x)8baN�l�U4+�\V{9fCd;)"~����V��$��U���X<-}%���qr⦋��q���,h���G�oH����Sao��<���Tn�e��8$�Y�AݍEr:�<�8�� ؑ�	��3���FEJ2	4���a��!uƞ'į=�S��\�G.>[�<�ش��F;>���kS�0�#��4籆�l�N6hͰ��#m��y��C֌��ڂ�������`lb��J�����-��=�x�Hf`F���(�`�M�i)�U��1(��N��K1��:�[���,��ÆMAkA�Y;�N�y5�jQ�Y���7դe=,9��q�����y탬�aJ�\#�+�{C�јt[�!^��D{*_�d�ϯ���4�״�Y��=���љ�6�1iw2�I�N�и�T��l��0�v�B��	S�]�O��(;��`�B�6�'1F1�xrFc����Hi4�Ե�_�G�D�4yZ���
q�z�MF<��e�X��ܤA$�����g��I��y��N�E����Y�X��yM5�,����aq0�M�)	x���	�u�E���d]�7
���I����5��D{���k�uJȉ�7ԓ�	�}��6��:H_�D�mX�l�yZ��	gm�m���A�0�� .&�&���=YV�b�B�i].�f�Dr�L�+�$7�×�>�>��U��2�C�^�v*s��ı���'�иAq��7�^�2$�p��I>{B
�>[��1���qF����y�>��$@I�,-�FL�CH��;��'�zdY��I	5I��$��k�����7N���ˈ@���H�Z#���_:Ĥ�D�C��I�, 	h��� �cQJ����Bv�W���Y9�qvK���&#)�.^��Cv������(�G�#�}	̄�}�6䧇>
Zq>�:%\� � �#
�2��trHX���_�)H���T #\��LJ@|���hJ��g���_��/	/���Pv�O��:dl��6ʸh��V�N�N �0���b���-"��6l�_R)��d_��6c�F�+�;����@4m���F]!㠸�>諤,���r��� �� ��ӺR���=&Z�z�j�~3��㘓'C��"|�H�å�;�=�A��ɶ��,
˘��h$V�Ϳ0 +�1��ID�~��ɞ��8�y�$=�[�� 렲>�]��#�nL�c���a��m���{�4V�B�� ��R�k�̢�����2��+�@��bI眝�����|^3��,{m&�o@e��ݦ�F=>(W���/>���_��	�dI���L97��&'3�ȟ�Xz�vT��z�>�[2���d���p�.%��G�T�����Dw���ͭs�y@����y����sD��C�9��Q���X���8����Y7l���j۾
�/7k�e�f>���i��9k�f�������sh$�r��.�z�Z����?�Dn�	���E 
[� ��E.ɇ���E��y���J��T/��彋k�-���M����Q��*���Ɛt0܉�ɪ��-��޹y3�[�ea��#�0�Sh���&����3_��7��[��k?���o������O�{��������͞��[�O�����)1��t�    IEND�B`�PK
     C"BY���    /   images/86ae6a4b-562d-4e93-9595-3c4b0d09f42e.png�PNG

   IHDR   d   M   PA��   gAMA  ���a   	pHYs  �  ��+  �IDATx��]y�Wy���cOiu���D�-�l����l1�JL���
T�T�����G��P!��J8�ml,�2Vd�n��eku�jo�ݝ=fgz^���1�=�=3{8*�����y����{����6p���>��=�!�k5x��ï�/Å��r��'�����p�1��^����}��k�vbS>߲6�jΛ�;��K_������Ʒ��_��fA�G�K@�%����G����?�]Yl�W��Ka��v?=�T/�׶@ݓ?�-��#�[�\��&-G��>\��3�Om���_|�#�Q����O���3Y�p�5Z�YW��5M�qX��'�F"�t:�
̙3MM3Q(J�,J:�.ZS[�_��dǳ�c�����"V�RȘo�ݖ���	�Tkn�O{�W���[�����}X�y�}�\K$i9��? !C>�WMڤw{Aʋ�"1�o�c�v$1���$)�����i���m��}V
!=�	�͐��;D�ve�d)vF���ƥ�u�,�h>7w��0L�X�u����l&��|>��T2�M8��4L�U	�2��^�By�ri���k�J��n�^4B�	�#�BM>���HC��;��4g�Y�CzГ�m�|g�SNR��J�^�fGB����b�4H�1��i���P54M����|������m�޷�B���*����0�:�էDD���qn1��*i��
|�`��SW[�d*I��j�mH)S�[Kd�c�c�k�8C<Ӈ�_:�"B&`�*]f���{ރ������A�3
�����4g�6X]���"U�ËUI��W6;���KX��E���$�ˤO5��C���%���Slw�4�[ǎ�^,���Q弿���ڥ�B�*��i�`��Ǻz�:�߶�k�ɶ�+ĘX��`�����U��R)����8z�(�|2���OȢEg�|�S���w߭�`�q��	8t��cf�5����7 tB�����C֤0w�|4�1�������[��[a�M[�Hb���J����ؿ?t��$�&�(����ࡇ��X���$�DK��o�J5l���$�Ih4�<ِ��p��wa�D�K�y,�̶�"�n�^:�]�������+]S��,U�=]G��{� ��JG{���.�������2�_���Ka���y3�y/�E�T���!I��y3��6�L���۱]����=/���_�я�������W�������C?�l9�,1>�`�'j��ě~� ��-%��0���
C�=�34�~'�W�Z8�fך��՚z���Yʯ�݀9򈫎Y����1��[oAz�j���>����L�}��$�SJ���w�~�#�³D����X�[gq�l
.�m
�3��F �$��=�#!1o�%�v��D�K�x�V_4+?�9��56΀I3��d�����MC5�#i*l��M[Ƞ'�c��:�GH<���b	�:��@���9�ָJ6����`X�i�\��Ї��S�&i������%<ɽ��!T�krW��L����n���)�����dդԃ� �u/�"6�S�҈��[[�tB<����nh(%D��*����e�n9n"����q�3�u�+
�r.D�3P�#��7�ꊨi�6V��;IeL!�X{o���\xŲҢb��k�`��B��S~S'��q�������q�����!�L�|�@�U�,�ʪR�˃��2!𙜛��Щ SΑ��bJ��7��@����ҝSSݶ��ɥ���zA��xR��&���%�m��!�䛺�h���+��lmPֆ��K
ɩ�|r:�0l�IF?D��ǜ��rd`��:�Hϧ,��YT��qK$�{��@DV.���"	2	F۩��8dꂬ�������olDl���Ɩ�����C��L���z��y+�x[�<�E�|^����S2 B:�뙉�3�rI��z�<R�69�4A���i���7���k��Ճ�=��!��#�2x�俋�?E����b7�+\j�H������
�,�<��	\��mx�����x��%���H�&k�#]S��9��W[5����h��S_��~f�c�ǲjwD»T���f�M[��Nظ`.�©�^��z]"JD�O�9s�^����\%a��M�J�������^�yR����ݫW����.w���y�����Lf{�]?��)�@��~s���u�e<� �͂��Iy<Xk�"R�}]�7m@C:MB҃]ݸ>2+�nr1�w(�$t�_jå������x����w{��H{�����ɂ���g�����(�+�Q�/�ް���<�6(�0�l/nݹz�̙�k##x��1�)�F�{��9��zV2��7��
��PyS#�~p�(v,]�?&5����7�|I9B�YEF=Gܱrn_�Ghv<y��2�̌R�`)���n��AʪU�R+4ZspHN�1��ˑ��J׫.���x�]�� �0e)���hot���xٟRC�M$�t�v��w���׮�٬Ud[�P��o�87�OS�ۯ��%�k��3g�)$%aHq-�U��^:-]��U��W��y�%�%
�[���5���IK����o�S�pm�7�!,�n��� N�������0�lBx��b�R���̪�����P{ߢ>�1�e՞%g�Ӿ� ې;V���װ~�<���w����	��K �Sq-"����UG㦉�m�����z����e���F?趆�T2Do��� �'���y59@c��m+��"Ѭ/�q�(�v�GӼBm(b�\��;���4��k�/���Go$ۨU���N�H�R~z�+�������Z��Ԝ�\�謃���ŧ�"L�ٗ��d�^z�ڝ���5��P�OtM�sY6F:U�OGn�.ޟb�VYI���԰Rd@�̜A��v�&�GBQ�Z6$ih�m�
�w�)�@�[��i�;Tg�s߯xo����2�)t�ڱ84�4�9��sY�ọ�큸�,\̮�JTWh��2�qgOmb��O�7AG�{e7����eF���_�P6�
ۖ�pM�M҄�@�!��̂���sB�ӏ��mF�/���������C� ��۶ۗ,A/��Ko��k`0�s�N�J����Q���U�����6i�Q��^���l�7���x���ރ��^�Ze[�_do}��	���o1��Hc0b;��'뷓wdp��2j����i��1�Ѱu�R��u(�����VN�b���s�J� o��o�(�����[9����	�k.Q ݥf�R]v��'��[R�h/���C��	��U��ה���sj�����]���t8�d�xϭ��c��#o�w�K|���@��m[8���C6נO�1l?X���xk��RY1~�{��Zoུ�n�;GIA�� i��D��U����~e���oQ�u�Bl]���e���������]|��e�kmL���^���Ǌ����xt�uvdI��eKhЋHG�����nHG��Ѧ"q6��.����mKa��ŊQ�Y�>��=���V���y�l!a���B;��^)kayY�S<�6.����m�Y1��}}*�U��xq�����S�L�\��n\�U�gc���$(G��MSD�ӹ�7����=��n�Dz�����)��[6�VB�TK{��W[/����ظpn[�Lq��]*o9BOk�a�hH�0��A�<�9*�`�&�!|�SY$�\����U����H4�*�Ⱥys���U	a����Ͷ������U��[�N�\�ё�ɍ��gR�����)Q�H���mi*�Y�uf��}�U����8��E��@HN�3H��%��c��/^���$$KqϚ�x�䩪\V>n�tf#>w�H�u�Dw7���*��6,<��t�hjJ�-+���`T�l9_t��f|򝷠� o�]Q�RYa���h�ߐ����[���X<����rŵHT"�
[����+��9q�:ZlB��VyCN^y|��fl�?�V,�_=�"��l)�j���U֗�w/f��*�����0��Fz�^��C�wR+otu�	�v;�p�#]�rV��*��i����.w�\�_��*C|�"mK�:^z|Q?*ƨh�<�r�u��eNw��jnÅ�֑�J�55;�5
'�l�o[��G��Y�P��&P����r���̛��%f�R��ܓ�U�,6�]���s�΀��� .��w���E,D�6���gs����sL���*]I^E}��O-)?s�4֐���kN�T�����=�u�eɤ��s��:�1�D���S��� �vt�۶�wl�h��~𐚅�)� va���d�-��x�T�_�^�"��c/�� �,���\�	k�Ơj��~���
ˇ=��CJ~��tᓬ8�m1!�i�
&^;ߎ��;#��e��T���b��[���-E4�'���(�Pw<��e9a;����F8$�fj�D�+��jk�<�V-#�IBTVX�A�r�V���xI�o_x}Cu/�6�yD3A���i%��~6��zW���=���:I�*��m��,N�q���s�=������QÙ�*V�l�k��cæ�?��_�5@d����\����W�q'פ�"�����YȾ9�eMMX�XOn�%ˆD��g2&��d7�^��^i=�Ng)b
R^E`��H�ܾ���y똷�����I�2aW�+�vC;/�nߜ�Z|t�;���K�h��bHi�:6TF��t���XNB��xV̙�Z�*r��_)�J8e�&�S�.d���h"d1n��̱�&����O��ޡ!U�U���l��ՏlE�_*�t��G-U��Uт�kҫ�C%�Ŀ.��Q�f^=zDw�˳d���N;G�[M:�SI\��S�'!]	3��8&���[h��U.=3���l���q���vYZ�k��������;�����ՏS��LS?k���'n�A�����4'0^�݉���U�#���rSM�J(~�ݷ�aO����w0c��B��y*�ˬ,C���&�V�lk�t�A����Vh��<��*YDp���{�͞�2fSm�,Y��Yn��깳�Awv�@���m[aP�@�·W��Qt��f�ّ03��|�i�"�b���>6�1
�z2��� &)�j6�G�m���B��2ֳ����`dX�7���S)�����}a��Г	D��,}pqf�=�=g�b����Т��%�0�B�J���r<3k#۶[�.�O��@�$x<kېR��7��Jז0�RP��a;��kx{r��Yj*LV���J0����9��v�����b���7�åΙ�(ĬYĎř�>���k�*,hl��G��i�AM ܙ��Q���)�e�VYs������C����J�%l/�1�q2I�8��_������ ��O9���<���Zy�09D�%q�t����|\��/��m4�ݤ��ϛ�gO�vwAN+x10n|�`ӂ�c�B�k~t�Z=Ԅ��Ɂ��4=ZC�߲w��pޢ_Cz�w�;OD<�vz���e�T����E�p	���0�˹������~����f3��;'9�u%3���6&��J��.g�X0R�.�k�C�n�����寋`xŲ(�eM� ���+�%݊@59	�8�R�"�w3BH��ג��JT�Ϩ�x�W�,�E�*YN��ߤ�n%D(20f`a\�$���i�v�n��b��:�S*���{����ҍ�bӫմ�
u{'�!D�#���NL��Ԝ*F��������J����^:{'�b��7�����T��|{"�^9��4�y�C�x�����T�K�8�f����|"��"��]��󲦞J�d�!��N]'�&��דSnأ�����u���I�E���?�l�}�}H��`�����Q����A��tk�,�hA5D�������J5x9A�6�jp
��n/.��}��
c����5V�F/u���ff�0v�<���o��$S)�8)�A�]2��pT{��񋗬����}�A-�BQ�$Jv7�ٽhj��㶲m!y������z�� ^��x6�A�Dጓ����FG\����s�R�����~O���N�V��^cC2�@MM:��|A��`�����awS�:O����ϡ��^���Aa|<����صk������^���^��?�43��\�Y�������X߼K�.A���z�Lmm�jD��&���}��J._���Μ�64��,t�{�U�%q������c�����֣�L���c��?}S]��C�y�o�F��+�/��ի0n��e/����d��Ex]黂��-�r���3W��)�g~�
����z��#�~�O/X����;�կ~�z%��	I�x�uu�SC	;!Q�g��,�H���\j=kw`�ƒ�hkkCC:eI�cz�����K��`�� 
}�$����_���`�:�\�}7i�zO��s��6$j��I6Ƌ�l9z׮)"x�D��C��R�"^�")�3�݉��6��P���T���Mku��c�&1Ĵ�5������N��,�X��V�|,���O?�	`ާ��0�����-�U*�.e�O�E�_���D�0[ύ�(i��%ї::q�����Q1#T|�����z�AgW�i&����������w	�|�7~@O��K��7(}�z�:^��J�Q~�2�fE�ĺewH�jF�4�R�tI��El5͈���,�2=.f���m2��R�?`��k���ūb���%�iD���I ƨx���#�Nl��_C���$ko�    IEND�B`�PK
     C"BY"-�' ' /   images/43e4be74-284e-4582-91bd-e4a77387caa5.png�PNG

   IHDR  "  H   �9�   sRGB ���    IDATx^�|\Ź>|��Y�*6�P�%���*��JH	�:�7�Ʀ�B����/!7��MqB5�&Y��Er�w���m��{fϻo���ju����9S�y��-3G%(/E�	��T}\�R�"�% ���\�R�7	(@�MB���J@7�"�r�D�JP���K�n��T*�B��p$ �C��M����7rWj�$��P$�H��%� Q��� E� Rt@��"�>��D}>J	(P�Hс~!���/�)�F*@��	(� 
�$�r	(X
,:�FE�B%�B%�]�������+@!*ED���}7�
��앚	(%6@d�ۣA��T*�2:���V��N�<�ԩ��O�Ԫˢcbs,fK��fkR��G5j�9AΩU7�Ѧ�� N*��[�,j��j�Zl�M�V��V�Z�Ѩ�Uf�
���&�Z�͹�ߩ�v�-j��T���iQ�,j�����QNj���	��\M(�B߫�V�c`�i�m�����v��n�8�d�k٧�f�۴�I׹�Ԯڇ����d �7��K��O��C}A?��}t�¸�{�?|?\����6�� ��Nנ��o��Q�\��i�Q�=�(��f�٣lQʈ�9�L�͎�1����~�;�_�[O����
W>��h4�W���9o޼�*���39^^'A(q�ԩ!�ϟ[���k���?S�՘�Q�E�Zm�j��6J{N�V�
*U7�qHC�S�@'U�8U���RE���(�E��JPi���j
v[�>���ޡ��7V��>UvT�Z6n��g9�+�[�c*D��{;�Ņ	!����~��H_���J.�����?�P9�ߣ�������i�B=�.�m��>��clXl��S|�������~�Inv��D�dQ���e�s��(�Y�	b��5j�Jk���QZ������j��5��o��oj��(uuu�9���N��m۶�z�>fРAB||�`�� u�R�Z���0L�"� \���$L�RԢP�o~ep.�'�l�x���J -�q�oo��Mi�?��`fg���jm��-]f���ĜɯN�{g�ԩ-��߽u$u8���ﮭ?q�xk���u�q����H�рb:=n1 �<� �@:���N*�1	D HD��a�gcc����q6;'����ϖ���������u����c�&o�Vq�N�/<x����$DEE�7^<�Z@�F�]7W���(��ʍ~H����M��¿�H�ɓ'������������k���_*+��ب���������t���RRRz �ׇC0Ĕ�+�Q@(Pi*�E� D !�3̋���̙3��9Y�̚=���#��ԏ8x��C��z��,99YHOOg�� ��J� �'E
eّ������;19`ޙ�f66���'��ZǍ�����OM�DF�����'N�U��<R[[;---M�y�X�g���^�B�F{3ᤀ#�����n�(V$����V��IΜ9#4�hhϚ��bv��"ȧ������p��v��<�L�~"���b{vm�~�8��3��~"����@an� �*��ƀ���#++kyqi�����k�����#
����_�����]WW�}�А!Cz h"٭޺%5��]����׾ܬ\�H �$�
����;���^/*)z&l�(�r_�f}Y�Aw]m�	�bbb�i IY�!fϊ�P�C)O�@_J �X��b�j�*̿ӧO �����=�@�n]y����cm-QLFF���VMt�
�ؽv���zid�/�ߺC�@U� ��C<x�4����H
D��g=��jt~�ƍź�oj���OKK��ÚgD
1"w��` �[�d(7�����"��}}1."#r��DFԕ����YE���d *�U�����!@H"Yt��*QU/	V�b��9���뻳���(.-�SĚf7n,����o]m�<����2"�iͳ �4j�5r֟�Wj�l�K��W	`.�
�f�������3J�8{��z_�
�:�Q�`
wu�[
5U�kkg��GG5AB၂��<���@D���Z��]�"���a�t��GY�R�>�/	r��!;�ߤ���{�-@�6w�H��/̟P�!_��Ĉ0�0�if���~s���'#��5�/���|"��G&y�6�(�'�e��ib���g��=&6/_𛙥��-e���B�|!_�sD����wfΚ����츯es��h��M��55���-��F�11"�H�}��?�'ـ`D.���@�<"�JOC���+�J̓ʐ2Pb�<���wT�,:���@���s��ߝ1{�cD�k��j��������@D{ͤQ-�"�����ʴ�'���G*�ZXxYb��Dえ�%�#��M9�SH��4pg~�ut����h�; �����f<�@�aÆ)�j��w���<ruM)uD]Q��N ����%���c�7�Þ���.����j���f�Ձt��T���<�N%jv��;M�ƹSJ�8c��7H~)����1�(����0�5AC3L}P���ĈJ�J�XQ���I�z��D #��h*��!��ț�&?1�
�۱��b���=w�Q�NYm�S�����֭Q�Mv���X,"��@�4��֨�v��e�	�QњA�Q1i��]7X��hF����h���t�<Kƙ�t�K� ���������Ҳ�%DkזO2�k�رc�D���x ��O(}9�x���
��f������a6�;�c������V�71*�Q��bbb,v��:h� ��lf��E�G�:�;Tq�8uWT�*��nW�5Z�I�����ܑ���V���ym[k똮ή�*�*&***��"`�L_+���'��XJ}R>ͼ^���� �!jV\Z�4b�֭[7٠3.߱c�$ 1"�b�r��?�� �;�i������hjkk;��ܼ�j����a>�����g�����`���?N�W0�ԩ�	-M��,�pm��r��v�F��HHHp>�9�T��; �F݂i�@��Ys����*����ͬ^�~}�Ag|c�Ν� ����:���G�SY|������J�յ/���[��n��&����s���jjj�����%&&����ߒ���fjF����_��m*WO�R`���ږ�����������::Z����������4M*�0�?����)/V�_�> ��)&�sB���a���:��#���~cFٌ'#��j86ׯ�Th��^߹s�)���P�e�	���T/���b8�'n�����d���`>|G�=�L��ӧNllj�?t萯���rӈ��.\�8�O��[o}�v���+������uztL̨������8�xS0�@���Q���I5<���1�W[��j��z��qsNN��%�K�0gΜS~�Ų�a54��u��;v� �y�GrBm�Q�� �OJJ�p��͕����V<� ���l>�Q�������_�ќ����>z�\�2����cϟm\l�Zg�0�d2�`��&Dfa�49C��H�j1A���Y|R�3�D@��p��)�����	Y/�^����矖C�ў={�
����v��^3��qD�{�i<��Nb����b�C5�|[�"G2%ڍ����.�Ju����AI)�͝;c_YYYW��l9+W��>y���Gn1����h4c���c� ��Eġ3�q�O�+s��$�P�u�{Ͱ������9Y�W:���9s���˽����ه�=���Tc]�ݻw_ ����Wz����<����'��V�p $j��h3�.~�D�`�Y,��ݾ;9)񍄤�5��{�,G�2�o��VڹS�r[������ё�����(+�S�����Az��vx�'�X+�1�D�8ţb۲sr^�=�������P��[�ѱc������Ԩ׿�k׮�D��Y����1�wީKO!�(�����v��)@R��=O�)K� ��Ν;�1))iyjzj���[��V�Z5����?���g�j���aÆ10�1����M�;Q��/_�/m����0�q�v��ǉr�gV�8q�e��I�w͜"�I��v��7͠�ysǎÑC�'4�b/����\>Q�����4�#���`���y0�2;ڊA{� L`A����J�:�Ui֥MyĈ;,X��k�}}�ʕ+5g�^�������� --mHbb���S��P;}\$z��w!0w@D�K��'���ж��������&0�3K_,++kb:/��[���eeD�4;p8O_S���h����C�:�h���+)�����!$�mP�F�H�mC��K��������7L��={�>o�Z׌�j�K))u}�D�����kW����*A�9G \��A(�&��w���x�-~�;B0䏊�����������;u���?�@��n�k���'lذ�Պ��������T�fvudD�
FyD���C<��f2��j�Z��d:L`Rp�j����~�TN�2S��Ld|�=b�[Z[�$�%��59K�m���S:����;W8����D:C�ni񐚩�2jOm�e�䯡K#^X8��7JW�SX���H��3ϰ�&��|(�ljl��;�a��1/_w�u�������k�deDhTyyy��͛o*//�yLL����X<A **ʮV�m*�ʎc�l�����n�DdSl*�'�C��#IH|a?�F���l6�J�2ww�L�~vuu%X������a"��״)����9Xp�upp�7#�A3�[3��pI�~����V�e�Z���Ǐ��|�������"����#��33&&&���j��d_��9n���y��ill��慶���f��I�VY�����F�R�4�9�d5iD �J�B�����\�Oz;��E�ټ��J̭�<���涶�V�ٲ� �`���?m�%�5��� �+V��tWk�ڴ(uT�C�Z�϶k�Uj�
�U� X�*A���@6�.�1��]m��K�ڦF�ŪRag�M�� _�,��j�kܬ�j���N�`�N�93��S?MLJ*��Ȉ!��N$s���D<%'?VI��`r`z�&���m2u���:�|����z"���+V�644Lk<����<-!!A��4�D��%��m�^|������1�'O�9�֨�����s4!>������Kww��n�V�TH��@  A�U���J�
6�V%ZAeS�U�+.꟝M���[��6v�J����m�Y�LV{�Vko�r���n�練P���r���QpF^y�d���TG�D����.�w111=����m�����L{kk�}�̙@w��b�{���/����E&�������g�y�[��4#:�;7�o�C��$��9�c�o �Z���¥#.]�x�bYB�ޔ,���[�.��������'�����y�,�O��4����.DdR�>�/�I�]]]�F~߈+F�LNNn\�`��-�v��믿�jnnf6XSS�-..�ܔ�����p�*[�+�����h�GK.���4;>1��
̩={�X,X�8J�W���}�Q��ի����E���$$$�"{��DP��#i;�U�`�I����΢�p����������I��^q��g�����
F����^���}�����U��f��G�О4�R}.	B����I'|"��j�ʙ�{ｷ��E5Xy�����}�ា����A��*p8 �� QSS��СC;/1�����eee�T�d^z�����ojj�������Ə��$Y)�N� �U�<�f`�`D��0%o���� E�/o�@T^^��f��Οo�/)))�!���Hұ��̳ Q��+RG'��i�ooo?Y�p��˯���SO-9�/�яF�駉Cݏ8������l�74K#LRV�����N\}��Y�U�-������-ZT�"��D�������߶��ޕ���D�jZI�P�`��f�&g��fA���6u.MOO�~��'#��L^x��F������RRR���#�A��1�`�E������Ƕ
�ټ#�`���a�t�#��lْ��'�<���~{BBB���B�:���ذK)��Cy`D`mȞnmm9�����a+�y�Y6)�ۏ޸~Ŋ)��n�6�^��2)�/����0�؏+���t�y��S*����)!�.Ғ)�� ��jݕ[���E���½�D�ׯ�z����Z�oMHH`���Y� �@Ҝ"��ܹs��'O�F_5j���〣��>��榖�7�KMME���v�S£; b��Y��;���l���j�3%��λﾳ2�A�7�7`����|������햄���p">j�
�Μ9�~���/r�'?�蓏�%	�2W�\�����ݿ�����L�"ړE�_ِ�:l�LOF�]b������w-^�x���#�D[�l���O?}���������h�����nmm���I��z�=�����/���d}M��K.����6Dҩ���·2 �4;���Y�L3�պ7?7ﮅw/ܪ��#h�������O>�䉖�V ѠpeDl��N�(|C��h5��ݟ�������0�����뗕o���̌�9Q i �I�8��4W���C�X�]��\��Y��}�Sr�u�][T*U�mJa<,#ڰað/��ri�)!�e���Gs����ϟ�����9t�C<��`�(l(��ӗ��~;s��-O%&&,HNNN��F�A�ۥ����C���i� �7	G�� "8�[��ngF�;�	����;wN8s�t�UW^�������`��3:T^��r�ʄʊ�;���J�I�\��.J{ ��Y�b�������tF������5�xg5m�@t���cƌz8� ��뮻�Û*��T��'T�?��jA�������ٙ3;))ə�@@D�|dL��8�!ȭ!�͊�(T��ʩ�P9��=��܊�}��%��߱CΏ�3%�=K�.��DޫM|��#���̱cG:t�P���\+_�;�h�D�I��2�`����6GQx����A'�9r�P2�d�#�<2 ��x����Sv�����;w��!C2��~��:�M�w+@�]F���@\��� ���8:�ĉ�C�o�;o��zhG�������4��P��b�߇:fĈ��D�p� �ܼ�ŋ߹I1͂�� G1�z�����������z���Κs��K��#힗_~9{��W�dfN:t(;���fV�������w�uW�D���� ����mmi��ܦY0�ѡ���̚[v�#�<�w �ۮ._��ʍ�7�---}�����hUYD,#�ڬ��O�[��� ���#�E��i��Ə?���� �`f9�O�8a>|�H�̲������ui9�_���ek�\�rJr����G#���0"������޽pC��/j� Q0"_Fz�u��iӑ�GזN�}���{(�2#�.����~�rZz�5���1�����ޓ6$m}_�ڗ�0`�{�>���ZZZa��m�����^3|w�������W��(�����?ڗJ.u/_�|�گֿ|�С�$''� ������ΠM3��`n~�=�ƍZ�k����|�,aD�Ξ=�U���yqɴz�c�9��K��s�~�W222榧�G����e��"��PnA���k����T��{���	q�,��/V}�$��+!�g�v��ׯ�Q6�����x���BqR��%��o����U�7my5mp����t<��?�����ߗW���ρ�W���:�ZZ����Q����#:{�LW���ϧ��=��Cw+�H�W_zu��m[����6-33O�rn��m�uЌ�j=�����Ҳ�/'L��%��+�_�1`�h���!_��pikK�x�-�H��̙3��ǏUV<���*�j��khh�CB��̜K.��m�!����z�5��;�^}�4.}=��^�������?cF�ꀀ�{�a}ŀ�5_�牖f��5l��_աI=;s����c�g̜������&��L���ر#~ݚu߫�_�/1    IDAT�=?dH�eÆc��c��	v��+���Ǘ�������M�B"_$!׀�Y���[ZZp0Z�8���v�����J������{eX��_��<}Ϯ��;w�z sHf
G㣎<P�Y���=� Q�hr��_�H��V���F<3�ज������_;WQ^�V�m����r�رk��҄!C�0 �眹c0���}D��ك�i���+-۶m[��~�d�3"i�����8
���+��K����p��j�U����Ҧ��W���<XHOOgǀ�<se�p�Y��s�̛��Z���ʔ�B�\��>Y���������fҍ���G�677�332�9l��Ů������x�z���WT/�Fi���/��F�!w��g���<�Y����Oy����K�|��!�O?{�����X$�G0�:::���6aP|������s&�|��)���.��k����y��e�)�?IM�HO��g�����=8f��/���~��>.[\�����?_����֖_$�'�GN��y�7���-��]Mɛ���E����������mX���C�-��̌���ʵ��w����tq�̲?7������5.�����AHT�[p��:m���hiiF�>��=��̙3��'N���������禿���y�˷��������v��������MѠM3���ܼ��-��+e���@�g5VVV���?��ڂ��p"�iF;�i}�رc�&L�Cq��̟?��τ������Ӫ�W�����6====55�mt�l�#�Y�͛�{�]�ܵ֯���@潡_�mݺ5��O>[���r{����' ���ܹs#G�����qK,X0 �3�/.{qҙ���r������ A�0!0�h~�,�Y-���l�� ��:��X *//O�b��%---�
w ��4��c�_�����A�v%�z }h������m_4/׼��[iF}��QQQw�Lݗ Z���D�?@d=��_p_zz�Z�<�(G)�" ���QZ�A�J��C2��-�abD�lx~z[[[���s��4f�|�A��(�����_r����%==�$666*11��@r�U�����_�7�+%j���O�X�n]��5kkjj��¾��bLt���|��Rn�?$Ͱ�J�?������ӧN�7n��cƏ)��U�����ݕ�|�ͷ���KII��xi�^N6)��{�����N���j}Q�Co,"xF��n�.���׹����<"_:�k�iVUU��������yqBBB*�ՠ���I�J�rE�x�ǿD�Ir��Y8�ύ5��k�������OD�ӥʿ��;c����_�������'�R��?:E:V���P�)�T�KY<!@d�Z��zl��
#�E�rMEEE�G�����������A��]�}D�vߓYFY�hs{{���gq�����t성�������x��O�>�綖��{Lݦa;����$T�8<�� "�B����"b��vOΝx��ŋ��i�Y���O_}�U�����=s��oҰ% o:ȝ,�dD�$╝���U'7���7z��7�{s7G���f{͜#G�>���C�IR@��h�^Pr��ڊy ��f�ɝ<��E�.����"�i���2n�>��������DD�	A��
g "E� x�L�O�A;u������/�'f��w��m�k��,//�=��G��߶������7�a�����^��dF�|D'O��Y��M��E�.Z���{|�/�DU����������M%''����(��Ii}dDXx9�J��q򹺌o&]BB��!����;���f���+G\�⃏>x ����V<RzOݞ���K����h��$4��)���P�#
8�
D��
uc�N�<i5��ks��p��w��LF�[�zuLRRRtll��d2i,��d2�5��j�2����7�F�qqq�Z�M�A�ٻ��m�Ş��hǧ�l��L&{tt����8K���.��rCZZZB���,�?�h���I�!Rl��nmm=��:�_��^��-��ү9�W�1���#K�[�����:z��+^NR[�U�ߨ�+ �o����f���]6�2}rBrc��d��f�Dۢ5�E�V�������v���m��lv�ZmU�T��l2�L���ϗ5C�k�B=p(綾^��7�\��hF���ƙ��D��k��Tj�B���vr�9ۈ����x�i�m�όO�Je�����ʲ�>�Zk����Q777���o�?�ꌌ5� |O>"o��ސ��eR(�9�a����X�J�:b�2�L���<p��:�麗��t��G���L&S& � !����L�S#6���m @D�$>���d����b����,m��V���V��*A��U6�#0�ǝ}B�ſ�Z��E]�� 6�5�U�ј�VkSBB���Oo��f��);akŦ�[~UY������A�%�b���]P�?�
B&A� y���w)��MP	(�Y�P��20���iooR!�<Ld�/�>WJ�yJ���,������i?s���h������#�o6��<x���S�N��F��[8�7�W�[���|!W@����B� �[u����C�bQ�Ӄ��>4�?�%�����fp\4o��ÿ�r5Zj�0�Lǧ�8��O�0�M��D�֭Y�m�_k�kf���':������|��!0��3����J��)X ���N����������뉤���a�{������eW�X�����L�2�n�j�3�Z�%L��d>�4T�9&���~����ҵ�J���F�\����-(�}���/��坕C>�/^o_�~����+�_7��E����K/��9y������voƠz�') VV(3_?�(��y�k��N
D��<�<]��t:))�"J�3c������됣]�ֱ���#�8|��nRم�̌d0V�hW=m�gf���]r)�C����|�x��:������i[��UgΜi�<e�;3�f�����d���T�O@ʆlٲe��mU�<O��1�RhPB��I��I�(�W���N�U�q��}~�QPeI�F�Sx?&&��b�GE��{���/n�ō'.��or��x��'Ύ����yww�5j��
�V��mm�qp�+�%(������#W ��[z�I�u�h1��֩S�����>�9{�o���d9�Av ����PY����P �iF�;�R�F\��30RZy�01#w9�v�ֽ��NRR�S�Nu��w3f�W^v��#3F+���|o�ɗr?����j;~�����F���hҐR�4��E�	}'��ҿC���ҏ@�qBT�+�	%�� +��#:q�uBք/�������^��}�D��m��VS��h0�^2t�p�a��c��.�H<��i�DQ{Pj��H���a�ti?��x��a�0�0�ES�F��g�������&e�������ݡ�����7��ɳ��Zj�Xf�L�K�Z��䳦i�����>BW4X�	�g���
��w���5���������ƍ��dz�ݳf����<�#;�_�>����ͺ����� <
��+��������j�b#_<10�Iwm{�lu9�SR "��|ɴAHC���둉m��6��Z-'O����y�?KKK;URR�k�������w�m8֐w��ៜ9}zbll�Ȍ���m'���q!�p|�-u���.���I��MЛ��[�uSS�0n�X}Q��;�ΝQۛ�SٲQyy���m��k�j�GD�o��!���:��Y-uB�*CL����=�����l���J�6  �ŉy#,�!cL���vӠA�N����ل��	�v���Ԅ���Զ����k����_�\�jՠ��V����Jjk뺤��k��f�j��s�}��l����h;�G�If�X�`��$��o�}�^�:��˛~�R��k�A>"DYǍ�szI����-˖فh��͓�o�����|���j��wwB�2!o�����Bv�r�>b��_q��nmm�������h��Z�jucbR�����\ziUzr�����sZmbWtt�Y��#F$�:;;�ŮU�TQ���1V�5���o�l�h8}jL����gN���Җ��ݙd1[����R223c�!May޿���]+��_������)����
�No}�  ���`DYYY{�K��={v�?�z��@�e˖)��z�\@$��:��f��蠄�>w@�j�%s�ۧ��M��Ę�u�JP���Y�R7k4�f�J}VP��FG���m�Z���6k��f˴ۄ4A�%[�D�Œb�X����c�f3���u�M�&1�_�$�@
��[�K�����E����@4!koIq񢲹e[�:�?���-7�����bD#�g�y�vI#=����o$k\�����M���f��l6@Ĥ���U��Q�FC����G�Q��m4<��v���#���6�@��b�M����dq�ܲM�.�����nܚ[QU��h0��D~�/�[ �]1B5஀HZ6]0�2�M��/� ���|v��ߔ�̳>��	��z2�-��T�(T�����⢢{�'����>�mU�+C�/@���7�9T��U9�@�g�4�)>"r���;�F;��Ned��)L)���
���+_�'��������&�����x ��J���r�r9��D���Mw@$=�*TQ��eD�+F��$���M�M\�NJi��7�Y踏�Lῧ���#��/���!�w�D�&w���}��{�Q����i��9r�Q�����+�p"vZ�D����@D !�����)��Op���Y���F�B�z)'�<|����v��lh��ۡZ�B3�KQ�Ȼ�BzŶ�m��n�x[aD!�E�y���RS���R��=���w.	�3��� �=_���[��� Q���4;y�0!+�`QI�ݗ\��1"M���N���|���C���_Qݭ⁈}��f����=�9�y��<��r�;w���b>"��lCY�
��^}�n�m޼9�r[ջހ(Խ@�@��A?@�H>��2�<9��J�-�={�ƈߗ�o˪�^�.�I��%�`40�(�S�pD��J�͞=@���Y��Ul��PQ�@�2���'_@ 
� Q R��x����0�1�yDӊ�=�F��zف�UVl�y��Q�(�P�t	��	�N+.]8wn�&9d ;m޼y��mU "��Uʈ�p�T |t�_�3E����xD���i<=0�o���9{��-r���@T^^9�z���]��\�4�~@6>G9t�W��#e���^iX�VJ��+*)�sΜ9[{OJ�+ #�"��A�I���\�Q�pfDrt��1 �(���-9v��1kެmr4Xv ��X1FtV�sV�ڰɃ�Dr��R�@��F�uqi�{�֭[Goۺ�]�A�� �@Pu���,>�=��%�*�[V%G�egD�7o�}[��
�1ĽXG�����s��(;+kwQi��gG�Q���WWWm}Ǡ7L�3 ��QdxDJVP��C�hg��_Κ?� �$dgD�6l�������0�π�����RGJ�2D@TWRTr[ټ�:9FJv ںu��**��� �c��:	��� 2N+�vۜ9sv�!��Da��!ǀ+u(�%�!|�+�Q|[�>`QaD�DP$>pD�������r��{�hm�0�ʭ����#��[�#H��R�"��I���O����d��s���6d}�P��@$��:0 �+����C��s�;.�6;����1r}D[k*ޕ+|���{iu��V+�G�< ���i��?�!9��'@$g�>,����*�$����:z��y���e��ϟqL��Dr;���1�J}$�0^e<0�Ϧ.�7o^�R�����/���y�`4L�#�H"9�H���J�#�t�ԙ��_3��}���m�v���m����	D�K��P�?$�l��Ĉ�K�Ϟ=�ޏ�|i� QM��z��&<Vʍ�B.�k�}��W�T�ߪ5�������D�� e������W��~����.d���K|ƅ?���bò�HE4<���=����C3fle~a����Lh|�W�UUּ[SS=�6�XL
����F�z�c ���'�Y��~���8!�6�L��1c��Oͻ穧�� GBj����*���/��ʸ���VW�Lt����7#
@J=��	��ȸ%��q�O���U�
��� �ƌs87wʯ�^��gޥ�!"_����/��������z�t,�x �m>�f�T*�F� �6@np��Q3� �s���G&N����~n�C/;���_G��>�����xt��A�i�� =��_B�� |L�50J<��$��H7��I�L3�0Gƌshʤɿz��g"����+W�u��Y]U�'eD����*��ț��������D�����}l4�/2��9?f̘�s'����V�XTP��Έ^|��+�+kޯ��.t��'#8�B�I�4*�]pU�_5�}DAiN��W0���"��R� d�X���ѣG�4e��˖-��1�}D��T�߫��^�w�#��y o�Z"o�ؿ{z�9$�M���� D���D���Q�G�4a�MϾ��.9�(;=���骫������~(j�|Cx�/��\�c�m��C���.
�G���^9���?�D���C2�������2`?~��pZ�MO>�dd�G��g�2��P�v�N7�B��OI R "Ӎ� ����q^��
�/l���	�x Ri������+
��߼t���<�^QSU��N�+sD=3�/0"bBNP��@���@ĭ�
#�	<T��ϖg�+Fv4iҤ��Ң�~���Sl]�qP�noUWU����f�c����M�fy	Bo �=�B� �TZ/aU/�V�b	l�G���8i����
n���~wT���D�;ћ���Y,ze���!!3����1������5 y29�A���$� �w�bb2M�pVgO�p b�h{՛:��'�3��uG� G��.^� ���o�����,j�
h4� D��Ql�eM�ٌ�!�O/V��b*��gE{u>���b�W�B���Q�[C�����i5ьdO���`j~�f��m�o{K��ͤp=ψ���r$@�}��ޜ�5���ҫp���Hd��"�� �gFV�o�t�H�R��>"�'ęf  �|V��D�NaH��ҫ0V�@$�����L3���'�/�Z|����?B���?YuU�;z��T�0�����0�Q����SK~�@���/^��P��N�+qDv�$�Z��H|F�W&�M�0S`�9=%�_�(�H[<ا&���&N�p z�箨��yW��)@
5R��*�	�Db�ƒ�%�E,#�k���t��yD6��U_�GD>!�'G��0n|F^�W-W|L^E�.X�Bܷ����Y��4�(�͙4i�Ԓ��If���q�����t5���Y-. 
��+�y�@� ���D@D�{��'��N��-� S
U�s��UtAa��D^05Č�	�*��u߭�ڥ�� rdV�D>�?FAvF�lٲ�t5���:]��j���x8�
s � �5�z����h]Z]W�	�cD9'n*�Zr��>p8����>"cM�{555�6��5����g�I���r��J�ž o�	�-��9���$�U�"T|ػ�#�Z+nz���\<��ֈ��~��j��}]MU����)�  ���Д����@"��dW�M�R;L3��Ȏ�8qKA��[~��?��7T��Q����z*��U���O��hxQ�X�ހ��a��c�e7��7�T� �'K��4@�H��:zg����� :��-��h�ĉ[�o��o��E}��@��s�]��z�{z]�#��d!�)@�R��A2ݬ QO�lbNNL���w��j�YQ@�׳���	4z��.��i%�=��zC��2��E(���    IDAT(�1bJ�"��"o�ky�l0;�����;L��������*k����TE#
ň(e� �0��9ۧ���cE�ㄞ{�W�k�3�{����O`�J����iG��M� ��Ɍ��J�"����]އ�8��s���`E*�_��pW>�t��V��'B���Uyyy�>���o�m�/��`DRGCh<��xpg�+@�ː)ׄF*A%؝�s"Z(i��A��f��$�'��xzR�����@dW�LH
D99ՅSo��c��L�|�Wvӌ�zǦW0"�h����)�|눽.Ke�@�� ^��mIz�(���`�r��Q��Ѥ���o���e�
����Cqd"�53�T�o4��� ��� ꡱ�9���(	j�"���Շ� Fx!q���
0��K
�P�辠�� �:<��Mp��R�,;;[�������9�Pv ���O_]cԿ_k��#��e�D=$� �
�_���a�[��lL&�6@C����R 
�|�������X���ƌ�@�8�1''�X�?����<�;m�V��@�l�Gk�ޯ5�� �Tl��s�� ���U1ͼ�����x�qww�����X�4�-��{XhOϔ������g��:�	���f ��������[~���v�؄�.��^x��`DuFC�; b[>��Ί�(��Vnv#��H�)�E���# BmmmNV�L5�#����U���o�=�L�j�`�Y���Dh�0_L3�����"�Cid�g�}vL����Z�q
������8��W� .��z�t!9�9ԩ���3I�ӌ��ZZZ3"��9 �3�&�� L��F�r[\l�  ���s��~�ՂU�_��>;;{g~^�Ϳ{�w�	D�?��XCm��Fc�d<ߞ�2�E�{I�{�b���3@�
4T�}�c|j��	�0*�O���Uhjjr8�E&���/;�eڙ�;&&FHLLd�T�3B�x�#G:>�G4>+kW^A��K�,��I�A^$;#z��g������I�H��QH��*���I��X*�,�`�b# jji���))b�3�ą�DL@d���b1�˰�<8�����@���6:�v�h���ф�����7?�ģ����5}D�4������r��@0@�@G�1F����oj�4�WPޢ^�n���I�Kj���=�������4ks �W-��{K��� D�-�.�Hj�1&���gX�]w3��'�jY�~|v�����_D�i��g���3��� �i�冹o*P "4�/'I�IR�`F�+T@30&:FHqc��eF���#�t z�O�e�t �,��0�+zUX� "���>"��q2�$"o���BDĈ&�dG<#��0�&(@�M���@�@�-��җ@9�2�|�!���d�.�ͽ��'��Lg��<3Qo0"j6^"���R�7	
D��SO@D�!i��W������YY{����"b�hٲe�juz �8"���A��b-	w�	�����'�#�|]�!�@��gD���.D�b�D*��A����#���1"��U�@����'��P ���˖-�R�3�g4�*@$�+u�"�P ��V���qVD��� �7	q�?��ӹc�{F�q��ll�`��(R3��أB��p�F:.�h���������R�*��'F�cxո"� ��#�� ��ˈ���|���]��8z��-��e* jisD�(�O�oV9�.��nTDo Qn~��O<���f}��ٟ�}�@�7�3�(��
��^��Pd@]�M�"v`�f��}0�y%�1KNt���3�Ĉd"9�깧�+4���1�#
�Q�
��Q��Rh�h�����q}�E�8��sO=7�P�{��h�Z"��X�E�����;��(j�y���=#��77?��'�xB'Ǩ�D˞ZV\[��h4^1��y�xpB�'��O��Xww������?���i���^o D=#
e��/,�����	N���-?-[VZ�3�i4�䁈��$w�G�w�.X���7q���6���_�7Vq��\��UQ5ju���gf9eʝ H�S���n�N�Y\|���dr5i�.vԋ���H;�]Ɏ��ox�>���G��,��.�	�h����):���b�Qc"�94��5N,BG�|���j�Z��x!|�C�������F� ��c@����?@Dmf��ǀh��M��������U�?+��Cv ��e3t:��`���I��o��HBs�3_DhLF��jgD�D���ȁԌ��P��E�D�XzX��~L*��R0B|yt/MW�0��A�C@�zxy�o��1�:���zp&��z�@�u�~�����t��ֳn)�K�C@��Q�q�����p/;���]<�����ư��o��n}��ǫ�K���{��c��Z��@Q�?AyE&6@�f�E��?���t��&!��$!6Au�󓋁L�ҧ��mC�|���0�z�����ɑo7~��Q�`A f:��Q��Žahk?Q$7�D���q$I�\
D-�-n��え����3F���ma^���=��vo�
˿/�h��X���h�<�����v43�.>��X�@D�u!��2o^�Nz��%������@B
,lŇ!�3�{�,C�]
R�_�	v���|��J
dd��R��m��^ %vp=�Ç��Ύf������L�S[y�i�Y�iF�b����� �
Bi�M���_�_p�cO<����wY��n������F��u��pY$ ?	h�%��}"R���m3�<�'�� ���D����+�����������'�KLb9�<$�飦�^f���
���P*��)��	1� D< I���J$@b��fc�Q�������NS]����s�܍_1" Q^a�/��`t��{��'���b��Sk4�=ҀH�� ��/EJ��L� %8w&1�/D̆g%�SL%|OozH]��R�Z<���zx3�o#Mrb/Ĭ��-�š� (2���G�ƳbehC��������b��vX�cC����rǈ�n����M�Fy�����]hll���<�d@-c���gg�/̻�����+�s��@�B�s���F��HcD�z� �I�$E4h{��=ހ���T>�e��9�<+ B�cR�o\COMII�������hoog�wuu�ɍ7�� ��"b��!-��F��@<��C`���&��p����sb�T;"jh�PGi����L�i��X�dV�T"6'�LĴhL�.<�mB���]Ns@
 �ܭv�I؃}�� /�peD㳳�+�/���'��d
G����V�\�9z��<�����h	@�˖��1|�Ť���+���l���/�����u 88 �رC��o���o�LRSS�!C�cƌ�.\z��'����;�<�Cu��	����#G�s��9'%����F�C� BÆc�9r��������' �P����ӌa<x���ԩS�p6�Ů�j��g���tU3�I�&	ӧOgL��� �Z�6[{2�H�(�̙3��``o�!g�h�\P� r����L�q�Y�ro_�t�`�����D��_[[�*��&+���/yDl�I��<�ՍD��1��W����ʇ���@�o�`"���	���~�#a	.��v�$�'�%��B�|�ꮩ��{�=����E"�
l@0j�(֖�����p"�JLl,*���B^ {^�`�����o��/bN<$g=���wNN�0e��+�`��Iِɪ�s��v���Mhhh`�={�:�N8t��@1>Ƞ���L' ���	7�t��af�Ƒ>��G$5����{ ���w��|�M���d1;�h[G�	�+��3����w��=5	��@T����%�_R�|�{|%R�Qyy�V_]=�h0����9W12)�0���^)h�����Jgdd���ؤ��^�`L^L6#�
�� ����	�l۶M����.��z��b`���  'O���  N�H���+L8�@�GgϞe�`v �p Ӊ�H��v��|�`��a�E�B�.�/F��)��&�?w��1Թ~�za߾}��DB#Ƀ�gVc^(������[o���AQ48��E�|D�	��B��˗+V�`j��Qs�8�Dۅ�Ryd
Ң�>�"��J ��u(� �WK�.���⮬�"DF���N����������w��$'2�I�.��b]� b0�J��M��&�ĉ�����1�Cl�]����&�'h���dr�M���J���_***���=Z�?>3Y�*$&;vk�`����i ��h��@�7ڤR	�.��ɓ��Ͽ`i׮]�o���5 �=x�`��k��͛��+Ԃq���9�EV8L.�/�-� A02qңM0���
�7oΞ>#t��9}D��*�!��n�M���v�:V����I��%��q�x��*twu1F���C ��M���a��G��s�Dgu=_ :\�`D������������&���'�2�B���U�RfC+,Vt
Wce�_���X����!k�$��,�_��Dȅ!�&	P�uL(�t�f�n�*��oc�m�Y���̙3CH$$'�IONY�>�=�=G��K.a[}AWl6���E8z��`4�/����Od��p�W\.�y�0{�l~ '��T �U���,�Vf�� �����9�۷o��ꄯw�b�R8��`}h3L�������N|��D�7#�1�	 �6�2����^}�UDh3sXGG���4`��ZZ�w��]-�}�#��u8� ���K���us]�3"�u���\����h4����9n���>%W�
�*�7��;� ��L30"61��^�iI��聵���A�,�̜2��#�i_�� XTTĘL$�_���hnl�;&|����l�^Ə��0w��	v��5�V�e@�ɖ-[��4��uM�:���`2s@ 2��� ���'��t� ,ȋ]G�Q�L�D��㏅�_�cm�,r���1b����_���L5`c�u�]45��jJ�) e&�������7���}柢,r೽����聋|�g����7�������߱��K�0��++�������5���
��)L�M2"���J(��f��� �;�j�ɉ�&	"V�·|����#�x�\z酮��~fҨ�¹ӧ� �֭[��7`0�~��06�&��.l��ڶ�1���zH������@����H; &�����1 ڸq#��>�B���]w�E`�pf��0?Ҩ��رcY���bq��"(uwv2_��kV}ጰ��@t�p�UW1�E_����1ߗ�צ�0����P<�'D��%���>*�;ZȈ�� z5-�N`�DR}�C :�WPx�ҥ���L��Nv ڴv���F=��RZ-���@D&Ej('�A z����e�qx�IFNk����\����2��S�&&�'R��`'���h���X�Z-�߻W�ꫯa�bG�0�`�̚5���&02�g�ffr ��	��Θ1�E�`�P DmmL�%$
�G���׿���r�'�3����ŋ�n���6&��C/\�~���?d)���$�� $��}76��P_����'�16��6���� c�Q��	fj��o�a�D�@�3>��Rh'?�	�ě@yVO������9���WJ���G���\��%_0��++�Y�2���~�7�_�)����d=�����-I;
��u�T.Es��Q.��p��;����=&�+�v���� �$�އ9���7� �>��`3?��9s�r�V�MCLT8��~�m���dB?P7L+8���� �b�N�C
����iV�zq��;X�0�PMb7� �{��BX}�p>�W�L:�Z*l� ��f��3gX�kV)�j8��d/���$����<����� ��Pg0_|�c� "b?h��d��>A$r�;$+�MQD��j4VNF$��=�;׬4�/-Ý�����޹t�k����/;}���Ɨkkk/alB<��`xj�
(\1�_E<�`�Ì@����"�.��}�'��%]xF)(������l�o�3)&�) L&Vz�0�|�V�f�Hb�#����0"�K�0��NIKY���6��+�0V@ ˀc���d�7���{�_�}����G	6l`yE`]`ow޵P��uױ���cD�O����W00 �$����%\��B~a�7fР�	
��|���~�R�sD��ʘO��GJI�}�~�&E���� 6����ӱ����� 0�yDx��������"���B�4��"5�\�4(�_���yf4S�m��e+��_���K�tn�s��@�z��F����sD�yC��*%� ϊ(�������"D�0�\��|�ɼ����H��J�D���;��0UJKK��L����ZZٶ�Y�ػw� ` c�������L)))alf�#"��C=׬Y#lڴ�E�`ցI�0v��ZP/�cx+��H Ą^�r%"~08�s�Ϳ�]s;�$Z����̮���2F�5�E�; f䔼\ff����O�b��ϳ����[�������LF��k�a�_v�e=���
�+�R1�(�8ŀ�rk�t,` t��sg�2_�aǍ�-��X-� �|&�(�z���t�%�9��tR6 ��:��_�p���V�(�^+;��^_��u;�J/d~��+��U�7��� !L�X��!ILC��T�t�+�̛��N�7����ʝ1$��C0o0���ҳC�LB���xjt:aSy93�0xp���D���i���!�ZY9��AD����Mj L��s�
i��=B�&�1��?���Ph	  ������P6gc@ ]�ӣV�O�`>�U�~&|��'���b�e#G2�lr�� N�+r������y������� ��� � `���c���4#�g2��w0.�����S�P���x�ӱ�b�m�űg���} "�����>�FrQAn�]K~��`�/��D����k�j���w#�?E
:���K�h��<���(�xfNo�L�o�3]�bL����`�wᴩ�I6�?u*��Z�=e���:� H,������e�YL{�


a��q!��l2����y��!�ȑ���bb�?�rj��Ľ`Ǐg&��H0Ė2]�F`����	���X�1���p���k�	�V�b�D�'ў48�s���c,������4��,��2��n�Ȉ������g1[ �\$���D'�}��y��<cB0��z��S��2f�	�#�@!X�7F��ؼp��+eg����4�L �a4�`���E���/�#.�]`�#��1��8�d��S��k])���Q��	ť��L���4��'7�8�-�32�@�r���o>��S6I`F`2Ä�p?9]Q.1# "a`,&MttK�Kb��:;�It*����'';�y�� ;w�V�^̀���R��9���k���P:s�����z�6�[��϶E��-"�_��B��t�p� ��je}G�]���k�20�LP7���$�C>.!�B� ��$��Y}�qC���4����@w�7�c!����9����lu��!k'#OǤ�t�#�gR��A�����d�7q�������y�w-]�����>��ʈ���c+�n��h0�PW��Ɉx �S4q� ��` ��/bD�{3��C"0$�������l~��x�p�7
�II�Ahnjb��+7�A���L�BY����?�&�/l�븱�?Z�Yd

+:�/���� A��$c� � �f͙-���	    IDAT:6��#�	�/j�Wk�@D�
l�E�o��aÜ���� �& -� ���K�G2"m�3���XX{ɔ�l {��b���c� ;��7D$��W���;��!=$ ��Z	; �L0O@�������?���9���QՖm7��j��8Vb�1�R����!�3M"F�5��偈�' �h�'��k|��&]˃/�Bab�
L(�p�-�=�9_�Y"2�/�o�0M�o�`JP�
)	e���G&��ѣY�6ks�*����S�#�� 2��`#p�X�2����v ]qi��_X�ܷ�<�E��W_�>��3f��X�2��a��-&<��κ,��|�����X6��X��I�x�#x�GW��U�E� 0�r�,߉�������4�߾X�9s�#2���{�(E����bD
	pf�-0�����f2��hu�e��DǽPXL�"(89B)�M4����R�?׸�����y�c{�F���az��'M�,da+�hV�y����M��;Grttw9|�	v�`�����1��20�P
��r#	v�7�r�h*�&�V0QL+����*�1]�������M+ ��5_1&5��
�	 �8y�� ���=��r 8��j��YM����u� &�	]��}��1���H4%-�!p`a+?�_ �L��@�2M��=0��"�yKM3Z�y��#|ߐ��wWD2���ʸk���Xkxf�Ν�,�GP�eCR!e/������<#�����i����"�Zwm��ҵ��� �FF�|��,� C5p|���,�����������H�#b*��E��Ʌ��y�,4����  o�&)��  
��ǁs;���%R�k��72 �i�M�p�B�pTô�Q6S�-(p�nV�X$� 	�`D�b� H�Q!|OY�� ������5�v���C� � ��~�#Nr�9 L/vTm\,3'`�W���Ob�	m���)�m0 @��� �M�"f���9�bNYo��\�T�?0�SH�(��`�ҥ�}���s���Y��ʸu���O]m�S� "WuDP~��\&�����O�6&NL���~����'&�qq�HUw7�< � $�i8كI ��li�}`�q�=_�%�V����DL&L,�B�&�,LLL8�Ѯ�$���q����A &(������3|�2�r�jĝ�d�����Ey�>"DY^Lx�,�<X"��{�@D@���	�O0%�o���Ľ(���q�l��|�0m�T!c��WQ, �#���h�I���#�����;'.�=t!D��D���x�D7����i�ΝL�_�v�; !vC@�	�7l{���DD�)|�vS�!�C88m���6���-𫰰����:�[���ر"c£nP&Xr��r�����پ/���q�&�C ��#���s�`C)&8��f� �nh`���`hX�t=3��,#�9r�0DͰ���X��|��@�L3J�Db��	F�ͽ �xʘ��eM����� �J2I�.J����\q�U���t&�����O��bK�DԌ�u:5$fV31I�D.q9 X���U�V2V�~^���O�v��`Y���`|5�<ZDImD !L*�1s��n����
��iN�; ��� d�?m����`�	�ո�r�����#�~�� "|�Dńʞ���na�Q�Y�v��Z�@�pƛ�=���p��Rf���ÎƠM���x�<�m0��,��X��tK�d�pѴ;:%&4�`5de���6<����޴�"�O��tZL ���Z�#�	f!�K[3���m.A�� �uO�Z�s�|)8��cǏ�5�q�	��ng&� �xP�d�r���8*np �<Od5� D����w����]��Y�xx99x}�ut"!�u'5&<�!0#�V���������g�<�۪��/�N�,dC�x�S�I��0���*������e���ז�E���2
Z�-e��_J��ĉ�vBH����#	�����Gz��]�j�R�;ֽ��{��~����=������-|�Ӕ�Vvl�'3�$�>'8���ʒ�����p@i5��|0]�� ��ô?3�*�.�����=�����"�i����ɺ���k��c��5�?�� d(!�� �E�Q��XYG{������H�VG@'����������A�w�;@ƶI��u,s��A���0��b)���L�����R�ѣL}�ڔ��b�p��@=
"�^Ѓ����DL���y�$,?&L����Y=T�f4@1x�;~!�D�H��p{43��1H�O��0Z�[d}�=2,|��)P.�9�V����9D3rs� � c�&ƹ�I����L\�> T@�7�$(��.��� ��
jςgX���L,�����V�������Y���o��� �8$\������G�M�6l�g��0��\�o�B��"`���"�3vl�#�
v��׳K�7!1ў|����;���P������x���.ݳgeyE妪�*"L;�1�K�牯b>"�4��zɦY��`��1PaB!;������4[����Tf����OYn�.ǿ�� C K������8�Yd=�NYgw��Hhu
�3`��"�B�>vs���*|��y ��V��(�F�ô��C��������c�4�
��k�p=�2߱�.v�pY۩S�Z��,a�F} X�M��E������; ���,�uh��>7�r�sI	[hǼD�[�w�n�)F�x"�.2Q����޽�***�VUM`���<�/�(( rY>=q�����{�]�?��i�W�f>�Q9�0v�h����f�ۡZ��Bj�8y�}�K��H
�����1c4f�`v�G��?i)�\.{��7���v���1P�Nু�
PB��,��Y�7�0E�%8���(�>"$d�2��G(i�cSD8}���|`Fzp�'��05Ŕcl�1=p��47��h�uC] 2�%�>�v��T����,kij��������c�� 3o��fv>M���̱o�15������Pa�c�!��1Pz�5c�*�#b���|��5��8"w�������r������	"�*&���(��Y�Ϛ�:4EL�����L ǁ|ǡN��HЁ.){�c�:fnؔ=��+�1����o�\����\���u�����a� xf����I�+V�n��V۳�ʦe6������߂�D@��>P(��$ �bqA�q���'Y$�*��Wxn(L�ï��Դ���O[��K6���B&*�5�1���ܴ=�BI�i�R�l/�����G�%Lc���n���m�u&�] Ml�V�L,��u����Gl��).N��X�c�e 
j�D��djC��ig&��oQ�i�î{�y���\�ϐ"[B��x���'�b��.����Sg�#x�م"�N�3��b�)��X6�'_6��2�66sc����R&g>���6s*�I��.�$Ñi��G�4BY0���k��kט��Wl,�� 3	>�`���9f��'��g2�׍�L� ���)�!�f��
*�Ҁ�V�Vu9����PO�&T�:�9�;Ϝa� �8r
�غ͹�J`��I�%K��n��v{�A�#~�1����A� �p _�g3t���c]-~�`S)��.(�3|O��]�3��B�I%I �y�
���7��q	�I���"��LR|��#���T�V?H�Q�	��c� L�֦&�?�K���i��&�ut��T���wٴ�Y�X� fOBR�s����hE>�-�%X� ��7�U�|����c����Fǆ�`A0%6`��Ȳ�0)ar9"�Q6 �����gp���3����e��H�z���g��P��`RJ�{�9b}h+k�3ά�a��1�XR��۠r�����ىk�CI�	�	A�����Dce��#���>�H��:b�]����h���������f���k�lr�=�a���gQ�0E�I���n��vHo����p��.�T�H0�(�z����!��x6?��#�&�tL��� P>"JF�&"�в�7N�5L&8��	����P�~��T�`���i�=�A}���v�2�E�#�"|=�����aZ�¤�z�!>v->A�c!0�
�`O�;�GZ�K�f�m�{aߋ����<�"�?.N�� *ݳguye���G���'U�~Z��̙5����*�Rfs�~�|�N�<R�"Z���Je�~Zt|E輔�&�5p^cV* ���(��%"9|2dNA ����X@���e(�25B��>��~0���"�1�8f��W�X��TW\���lf*
���Np=L��w�8��2cX�|>�LR̦�6�̑���=/��%�3Gnm�B �	3�C�}Q*\Rl��G!�m{;SD�L3j��&\��>�>�(�ܷP��f�"�i��n�p��� � �P��b���ُ���&�k��4@�x8�	D���n��3���"30��Y�l���@�c����==�W�BZ�r�g P������җ�z>Z����9r��))�P@�� Ǽd��
²ZZ��m��C���q�d���	�)� �E�,9ބ�����cg����F��y7|�pDc��@�g��K�<����C��f<f�Φ��QD�a��G���ȱi��%����8|9,8��p�kh�o~����L����&� ��f����2 B�"�0#��Ek��B�5�@��q��������iy�K&3; �%x((�	� 8�4����N0����5��������P6%�g�G.g�H��o��)��"~%ʂ�cɤ�}C�����6����)e�\G:�r!D�G�D|�	�gD��"���Q!U��|� �^� 9f�}0��2Bo]Jr��ƾ�����>�X��zvQ%:�9�����P�0�EY(% 
�a�R2�ڀ ���D���ehǂ[Z�EKN(C$�C��X���
�/8�q�,ǑMe��k�k�Q���s?Eat�/������xf�`C�&[�cO��� .8�'Ň���h����;���g͢�H\��D%%%cv�\]QU��o�#�.�A�<�71��oP|�̈́�Z9|�\ ���8"$�p$�"�6%��=���B��Ǧ�vv�;��еP>��2� �d�0��1�.)"?�#��k�B#%A��8 �(��H�����	>�W|�u�2ٳ҆�\�OR[Tx6  �>̙כ"�iU����v#��)+�I�M�{���v=W�����X�&����(HK$G��	D��嬦l�(jHtl�D g<���8�10rK4p_���B)C��pL�>(�m��g��{��!ӏ7���!���@#"\��f��� נ%�2�l�j�)D�9�'\a�r> �G��YBĞ�Q�|�P]��4��6�4��Ddud:u�<ߟ����� ڽcǪ@Κ	"ʊ�c� �~D4�p���H� B��N�ߩ��ϱ�F;�vP����e8�v�A�@���Vșb��e� �Dit/�����俢���7�h@�j�t,=�U)-�!������r΁�����hI�@���@G�B��{�L�Y����C�9	^,�:����$e�@����^�"~Q'� ��Q�-��
Rx"����Q^�I���Z�a4f�=�)%2��7��t��,!���GxS�~����f~��>�� �5@�iȭksWD2�p,�f��z��);�t"�g$�O�Oע{e��9�8f2��M]jk��	�Qn�(��Kb�ț>�V	^bB��\կS�Dy�wo���V�]ܯ�B�#
�"�s�%G+/�ɯ�M'�麼IC&~R^i̞� ���s���Fe1ecߣ���ъt�$�w��:;)(Ǣc������j�~䤶x?��:"�8Z�O��3�� ���t/�|d�� �� ��&�&�|DBuǫ!! ��L3��i�}���țf���5c��x���̚p�5S}Y����G�y��}5B�];w���{���"�C��H�~̀`F��(��A�oFR�'sùH�����O�q���x�B�!G7uv�l�k�>(i��=�C��@��l<���D�MТsh н���+?XɄ��3�������`N�y�LX�|/�Q A$|�^\ݵ�u�C1B�D�@q�h����F��ߘ.�ٱZZxZ!������r��4P1{�T ��B����Wg�����A/TW��	��;΅���������w(":�/K�HqKl���Hȃ�LE$-��A ѱ��ܻ6l�P� ڽcǊ�ʪM�RDb �ߢ�e����DB$֨���}ܽ��A����JS�eC����M*�Q9o�	���Չ�����Ìw��*������K3r�ˢ2	N��C.k����R�)(��j�F��2!�]݇�4;V���G��rm�	�"
4�\)���ߎdnP�!���J��|���4��2���s��kA��{s�3�D�P���?WוjZ�'4�<Տ�{�Ã��<�\�%��q�O�ă%�wG�@��g#���ڃ����#������	v�?�;"5�&�^�=�B�V�+�[�aÆ���>߇D���+***�"V�P!	%��Y�@T�7e��(TBb�H�����9y ��7��	 ��rw]��8B��� b�b���LRa$�.� v������T�l�����`��G֕x��@|r��ٳ����@�H(ՙ��E��Ö�o����L�ex"1 9��.fA�y���W�y?w�$��de'�!"'��%7B�D�x}�""U$���Ď�
"�#z�)"�(��`�#Q��naG�AD⏡�=!��vp)�ėc�=)"O 3-·�y�r^��a�	J�zd�
_2b�,f�H���&������$�\�=�Zk&�4,��N ��M2Ͳժ�����6m�̗���9^*"_���0͖U�W>VYU9���������8��I��������Po�ǽx͎��+H�<��Tn�����]���3DR���3�)�_���#������ ؄`G�$UI��>�`�������%����D�{�,���z<� �7��:�����7�O+�l�;���$��<D��@|���X`�������]�=]��[B�O���sL:ǆ����/�P��|O<�����)�j��7��#�'�wTHA���uiey�"FT%#aG�I&6P=����.�������i�{���Ϛ��Ηڽ�)aR�7�*�GL�(� b�f9꺂Y�+�?�~��6��� ��ʊ��TVVN
�i�wB~������\�̈)"��o�k9w��H�>"o;��k{����pw�+S��'w��KQ�b �ay������p�s�ٹ�E��{7�p֌|DPDDum^A!Ѿ@��XY!���.�ꪞ�j��h��^���B�7��!DU���@�@W�3�su�]�G�+ �;r,�t���L�$�aw�B��0_��z�CRa�jn��;�$t��u����l�ֹ�Qf�� W������UHѸ�V��\O8�R�>B6f,v�g��ܚ̎�1��([��-�/X�~����h���h���#�ݲP��zR*��9�W*$+�B���Y�� (�F��+XK}n�輙3�����!:��O{E�����#�Q>�\�@d�V�2Ǟj.r��{"�J�2�}D� Q~a��7ES�D�����V��V���T�־�sVK{�x�����vuzKS����uqq����p����:��O�m}aGf�oV]�|L�KE��Q����'�A;��GD��q-#╾�>�M=8�_ "Ad�yE�4r��&�0o�"2��:I�    IDAT�uaTcbo"O��Ӏ���t,��)�G���A���7�U��}���f��D����HiJ�y!�#��l��|�B���yE�{Y���
���ߴ�4�������5�o�<�Ӳ�;�U�'�z�d4("2C\:sELO�}ޛ� O'��� ���H]�D�������y|G�'����/'��PB_���_�VB��)���p������6��@@*X R�U����oZ(���!ё�;�:���z�$������T����R<))_���<>'�A�wZ:�
>N6�����<J�0WL��0�p&(	!����oRP�0-�;�x��s��D�@��Q��mܸѾ�v�?!��͛GV
@EDWo%O�ơ'��P�)�2[:�*���P
�"�d�I�� wSߋ�4}/E�;�ҩ���i֓�����Q�h�;Peؽ�V߻���Y3��X�W�t����}�}�g�D%%%�ۋ�t���"�o�oO3�ӿ�ao����iq�+ "K�=��'��|��y���{��C�x�S�b/BW�*tЪu�{���b�r��/�u�"�ʐ_��t�ƍ_���B�۶-���OD�ȿ9��"�1(QF ���^��0w�ܠ���
G0�%TE�<c�����C�,O�)��\���'H��2G$�y�W$���"�kď�g��6��-ݕ�{&���5Sr��lڴ�������Y�ѣPD���=�H��_�f$?���r�N� b��s�����C�9���L�	��S"�E�.���Ba��r�_��^�q��G�����,��ܼ/��
"_�%��N�L3���"��\����|,��k��DA��FT��[G��Mũ��]�����Ďw������D�-�:��F�_X�$"A�΢��zݓ�q2ۻ����M�e?�j�p �dm��M�#-59}XE̺�2��i�i���"1�L�wr=�q��2C���yF��\� *޶�#��" �?l� }�2��G�m�a�?��{�݌�g
����*��� re���3���?�	|�b�;���J��v�ŵh��
{���E�i��������)"���j r�1�<3=T�;yz�(��- ��]�B���N��?W��>_�q3����|�usVG4���m��A����X=�m��s�i&�v��H&���	�yxV�QUD�!�=�������"ڔ0�!�1��.�D��>����:{zј��і-[F�ݳg�1
"g�����9���Aj���X'rX�b�}GD���M?G8��~�ma�j��]��ܽ�<�x�E���յ��yj��H�1���/���{�����?��OA��~c��D�P�6��7�����R���� ��؀�z�P<sX^��*�!�X�@�Tk��
1}y� Ѿݻo7�O�ƩQ��Q����
gJ���(�^cȏ���Ub *��[�K<�h�Π{:
"�}G*$�1Ʉ/o��MP�58�'��D��kqDCyѫoqƛ7o^~��|���LD��'��y*3t�Ƿ+��������Qm�]E^�@G��y��JA�ꇮ��\�K}No_'T���ȷ�L0H���Ԁ���nܸ�`(�"����#�-��<7�� Ə�WW��{�>5 E���.��`�ƍk#/guD�;�TyR~b����?��>�_���1�[;��?�/�������Yg��i���5s�
a].e�;������0��8QC~a�����K<����� Q4���`t�N���!�2���R�=fh׀+�T�c�yH��;wR�c���рF�M�j�^���� ������#�D@�e^A��6|�{9���f���9'A��Y��>�= ]:zok@D_��ܰi�No�����vC�<����ﱋGt���M'D�hjaI���UD�t��9C�D@�uA^��u�����9�ʏ]��#: 
��	L�I���EA䩆�ߋ�(� wՆM�CQC!��<�о��CDn]��DW�h\�y��QE���q���yy��=�n{(�|P@���~g4��	�i�πDy���*b�34��и�@�Y$������Vox��m�xސ�����w`;�(���,���E��^#|j��
���\�غ�P<M�Ath߁�:��@W���ׁP:�~�hygk`(�@ޛ[ETPp׆MoE�)����F�-�uG$���F���ך����֬{lݧ���;�A(�î�٪�D�߇�|K�C�~QF �%�ˈ�h���C�S����azQ���p�M���7lZ�%-r�l�g�-���OD����F���ך����Hyz�8M3��Ic�q�`,�d#�S�"O�ğJ���u��H�i�+,X2Ed���ryh�DA��}-�O��+�8d@̇�Q�A�k4A(�A�_+R���'�`Q��9�W�>"6}5�D�~�^�0	%e	��f����Y�VYl�0���� ���k(|DCX\�>�T���@4����@����n7����Κ���Ox�@�$P���Dyyиs6X�N�>,z��ض���*�h�0x�(�\4sV����A�} ��1��o�6� 
bkD�v�@Dn@�7�6���qD�n58�)4O�׊n3�^gm/�a������UD���h9�j�g�:�1���l�g��f�a;��2ͼ��D�+�n�!s�� Ri��

��쿡x���~�v|v������`����'���e15Ry�RG����/k���Q��{�yyK9\J{xs!>�����>},�����]Y�3z���ᬿ�T������l����3W�D%�K��<�}�0��@�R}1��9�6:�f0��� ��)u�H�t�O�z�kH���txŸ�f�3��İ�t(�Q�T��/���M��k�{s^�A��mK����R("$�w"_;�7���ul0�9oD;�"��`ݏ�����TN����8�:�v��F!�T*����{�=�n����󠐂h˖-��l�J�Q���`�����;��I_O{��ݛ���陽���3���J��M����`ׯ'��rE�n/(ȿ�#k�	Ţ���h����>;�s�A��h4�D��=���x��/f~0���v�AUnn�@�����y�T��zp7���ܷ/�9�J4�h��#�((��YZv�,��RޜR�|���ť�~l4��1�@�
$�:������=���Vv�ʑz=:�S}y2a�X��襂��t��^�������~��i-�ҕ�>�G������ŕ����y����o�:�x3��>��p须�z@t1@d��UDR@lG��@��K�4�T灺7O r��\��C��3� ���d�X<��o_V�11�M�l�7��?��}gӦM�=��R���AM̚}��&�N���`����7�}?pv�ޣi&�#���A޼ �w��2�F�{Bc�$�˭0��gڗ�s�v�:����������=+?y��q��og�A������*�uD����yw�A>ZXߞf���]�����ǲ�z^�� ��}D֘��n�Ri�/(��ڍk��{�b��IC
"����s��J����6���Ll�l�\f�������ـm ��z��f������[F�d��bbb&�l��Æc�Ç��������
�� Be{2M2h@�4t.SlV++��j���6|��������3�yLLL�\&��`d�rY��&���l16�����v������h���g�@ZM�������c9?�@�M��&��cP}2ۀMfg�5k�YmV�Un뷎��.���I7n�H����7�KA��b���)��z�zE[����1�]�����u���c��>�c퍍����Z�1#�������d���n�;�0�1�bd2<�����3���
5D-b�d?�����cb�z���`��V�����U.�ad�Ym�11�����޾�qÆM���:lذx��7�U����7�kR�qqq�m2����#��m=�F���;̬n��`c�kE��e�1q�2��;>~dkfFڧJ��dӦM&�]3 �D���xab]kݥ6�m$QdE�<F6\&����cX���˭Vk,�VLg�i�ә����v�9�700;梱�c4(ހ�>:���r�������]r�.�dۥ�'�������c��;������a����o���š��d���rY�Lfu���0�j���X��ܶOl�3�Hl�����X�5�j�ϸ�~[���x�,�����g��������=q⛹Mǿ�7&&F�g�
�x9�+�p"�Н9s�墱c�uјq[.;�\d��d#�e1V�U;�g=/_
�CǇ�7W��W��翭g�@Qqqv�Z����X+:�<66Vn��Zc��X�<v V>k?.�c��d�X�����i�a���6�@wOψ�������ל<yj���@
�)��$j�e/޸XV�����;>v̘m�.����L�P�=z�hkggg���7&v�([ww��و���>#@����zqll�l�XӦM����v���_y%�ر��o������Q�F�Ύ�	ހ���@B���3gX�w��i�O�Y����P���ԓ7�N��*1wv.���6f��E]�d��dX"=	��������NY[��ZE���i	��[r�m��5Ծ�����?���g��^����7n�l�ȑ�O�N������P��*0�ͬ�ѣ��<e�����r�-����D�y��k����z��dyy�4�رcϙ���'�x�@��I&���0�P�ɓ'Y��8qb���W�{�FO���E������?�f2���舻�K����Y<�u��c�^&�Iv�ԩ��Դ{�TY%,�ۂ�y�嗳+*�ovZ:sǏ/�yE�	�}J���[�njg
��/�u���w�}e�P�a���ҋt��?��ҭ��ԩQ��Naoo2%����������	����w�ԩ�ɉ	���Y��ƕz�[��:����Θ����.�&M��N����va`w8M�}N�>-kmmm�Rf?xշ���y��uK��p:�o/�mNE��׺��2�_:^6f��WiD��d�+���K����[��n��	�H�>��Uw�Q0:����/�5������'FL���s@�k��z���;��ӛ4�`�X�"�`���I��.Y��`<�`����(a��Cm7�_��|��K�'g��A�|Y`��:uJ���r*K��h�̙�����m�l޼9�������纻�&L���4�;`�ڧ^�� ddtuu17�|	��)˗-[vď�Cvj�)�����U55��t�5'O�dfL3Ǵ:�E�L.w�i87$����}ʔ)�)��W.]�r_�Z(�UT������&��j��01hP��;����%��$'8�����-w��__3s�+9�_���u��555#�ݻ��_����{��ɓ1��T뤼��wz������𷉓'R�'�X�d�!�չa����/����֠7,9u�T�ް��X	oAD�:�x�@��[f����I�ɫ/_�+TD�9��+�).N߻������V� x�w���b�鳧y��/�� (��f�J��ݕ߾��+���#�O6�%>|xT�Ѹb����vuuM����/>���(==�ga������W����SI�)+,X��J������iZc�﫪�O�:%�S���(�)6kF�ϔ��!�;�"hk�O�L�0����ikV�Y�ӗ{���..�>p��&S{:2楗^�nW�3��_���S��9�O�1Q�R�z�ʫ�>7o޼�ī��JJJ�4�5�9z�l]ww�x�U�f�;����E��w��2����Ί�4i�195e�ҥK?���8?Q������i��EPD� %a4���aw�%^~��?��$��k���*}�d2���4�1��GtF�R���ܫ�����n��S����*Ï�=�`WWץ� �A��|)�� ���&O2�NW,[�*
")���1G���P�{�J�]z�ԩ�@�������A4q��֬Z��3�o|��k�.���o�Lm3���M&��̩@c��&�?@�Y�����F�缂���p���p�tk ��R�Ѳ#����f B���)����PD������)���ӧ/[�jUTI�Ho�a ��=^U�]q���X4�?����B��C�$\v�]+|�no�{(����V�"��1}ߩVk^�sE�o���o�r�ro QU��G	�4c+K B�4iRu��ԥ�"
�k �Vh�ku+�,��������x"�ŉ��*"NYfir��E��CD~���Ç�U����ѣ����$ �|D�p���S�K�>"��߷"a��0�oo�]��&N��6-ᮕw���Q�@����5C��9ߚ��y�N��#��YDe?9r����`�f"���A���X�d���{?��o+��� ���=n��B��k�� .�(`��ĉ�	��w-_�<����6����>`g5]��fOeC��WD����9*�kW\����>�g�����[Vv�������v�Ý"JJI^�|�����^3,A����Z_U�"��\MߓpҤI��� r���L31�---=3Ԛ׮̿�H�ѣeL�4*���&U�&�JWDޒ#�Ǉ����]^U��MUeŊ'N��� <�ii2�Qt��:���c��qDp���i�j)�w/Y�$���wnݩ<����9}O�I�Hy�""i4���ʛ���ot���r�iؑ��������@D��|_��p�I�_�!2���/�NNN[�|���"
D�` ������jى'ؚ(�Wp"�+�*D�,�@T��H�{����X��8����2��fy;}��U{{Q�Z�׹W���>��{��5��)//�b�0gu�A�o�?�&9Y�,
�`PH&��QՓU�ڥ� �<|��7,Q´iuɊ��X��8H�7(�"��5���^qUd:� �Qyy��P�h	5))I˗.]Z:(��ˋ��iVY[�;m�n	�s�iFKhe3�,\)"w�{����H%&$D$�vmߞu��ȔbE�:{n�cCr�^�`7�ģ��������4_�P��X�x�I�1���A0ܡ� ��J�^.�h��BBo@D�>����:Ezꏖ.]�c��-������7=�5op1g�Ӭ;G�y�p���Y����>����b��ba��0�hm%^��#�"JNN]�t��("�A���l(_Ng ��z����ӌ@D+�ݕ�/|��!^���ui)��/_샏���򥾤�SRT�y�Ё�<�H�4� ��ξ��gu�F�����_E$^' ������lc�@>�^:�:--e��EQg��1��1,��J�۪���B 3tA�����;�آ���f]9j�˅W�&RAt���eee�X,��>؊�@4a�D�B��l�ѵf�ID��'���V�G�Y3�$����@ěe|�ܫ+E�Y3��a����:EZƚ%K�����*�"B���Ȣ�伜W0�7������-_UQQ��b�L-�&��K�,Y�D��4+--����>����L�H�E+�]�!��3"(Q�G���i��Y����Eښe�E�������8t��&��0� �t���m�����reyy٣��#B��O�4I����tٲ��T��PD�vJ�0V�A��� �""pD�	5��Ի�,YQk͊��ӿ8���m&ӜA �K������|yYY�c�eb0�D�'O�&$$/Y�lay0�a��KETQ^��N�e ��="���8��<9�%*��ŝ�W,���� z��d�"� 2k4�g����o���h QYYŲ��r�hR0A����'O�LIIZ�p�ª��[R�~ *)�Vn�|V����@ӌQ�AdHW�ݹh٢�R+8�۵m[ځ�_�f2��1�:�j͋3s�~*RAt�h�Ҋ���C"8�)g��ɓ�S/]�@}0�@����+�*����wx�5����!�T��_�G�OMKa=y�    IDATY.ѪR;�D�.��J���Y�z:RAT^^���� �lE$ �II����n����Q���Nw�^L�2%t�Yb�V���zI�l�"�c�l-Q�~^��v��[��Z�y�ʫ�>����>����^�0�xM�2�49y���VK��y\X���R��N�]M�:���TMPM�Ą����Ջ�/:<���ݵ=O�D?/���d�vD�ծ��D�SW-Yr{M��(x%�%�*˫���tl��@�*�ܽ�-p7}�X��H[.S�R��ჯ����D��c�������3���+��♨"��Z��F�IMM^�`��Z�J�Ya	��򪧴:�"RDBg5m�(�#:������dr�ܹc�KQbByzrڪE+m3�j;��H���C��L��D�t+B�r"DG��/����}ה���;w%�>����fl_��6և/��]���w.\���@\#�eDA��Y$m�>�L���jɒ%e�n�P��@t��WLmm�j)5�篼z�����B"��l��LOWܵ`���P�%_��W J8��H�iAbR;�C�l2��͞[�̵�^k�~"�>���G��
 k� �@*"�:�"���i�
E�E�5�C�FA�%��R+�X\�+����S�z���~mDRk��q���_,��uM����K�]���	�o
�M�v�6�"�GQyn'��`qDgu@}D6[��~�Y⑴��U	����d2]j�r���)|6R@TYY�xgg�Ty5.(8~��D		ӊ��24��c^8H��"L��%�\�ti� �WP.���(���_����~}D��b��}ѯ�"�@�vx9��������-X����=Q�J
;a�}���Y=�(RATz�ȟ�L&�H>v�X٥�^�z�0B�+z��Ud�3pVG��Ⱦ֬raee�o,�5����p���O��SQ��9� JL�"U��*�Qɧ%I?/����tC(A���ҡ�Q?_8���H4� ����;��+���@^���*�(��� {��%���X���"r7#!ek!w���P��F�v|�c��#�����
DR��R��l����F��+���H��/**}��/UUj�tY�@eb�WW�j0g��|��ܾe�f4k6mڴ�i�mezs<@D���@D���4]����t�9�xLO�HE}�š�L�����Q�9[�~ifn��n���6o�A8��t:�2�V�HwW�$!� OQ��������wGM3O5����vJ0�˟A) �/#L�B砿�'�U�fh�v895c�����Ejo߾=�p���M��B��l������'"1C������Vׯ�tk{�{&�G�+�@����9Et���p�&��吖A�� �4 �X%��+"��z��\�f�g���Z�y��i���b��h��YD��QRRr�AW}�ޠ{����̛AE�4bL`���iӶ��+�D�7��ű �Q_��V����GD�Fh7Z�D�������:�@���(���#0�n�"r��W̜���[���š �^[��`�=���{)�ȑ#�
<\��s������B���;�xD���[���\_��V�c�R�b�+�o>|^D�Řt�Bӌ|DH����x��/^�ƳV������.�Z�׹��>� ڳg�%��ڻ�z� �;@����6Qqz��Ψ"�] ��˟��t�K��7$��\9�i���>���ăɊ�;#D�y��d�%�����f��|��o<�.3h����Kt_��1���� ���w�4�#���hGVVƝ��� 5��}��WU���t��d¾f��+g5��ݾft�Di)i��<�6[`|sPD��n�F�ڬ���"D[�n�����^��������� ���!$�i�vfgg���HR-zо��k�����[��!L��.���ȴN���W$TA��uRG��4SDӧHMK�s�z��|�Q��d��å/�ڙ"�	td5�D0�P���<y�w+U���̟�H������}��5��X,��#�"��Uh�?=������ӧ���Jw	"��P�ܘ�s���Xn�+))I�6�<o4�AD��B�sL��*ru��,��& PrR��dE�]",�r���(U���f�m����OH�4Cq$�������5ƺ�kkk~z%�L�J[�$��Ur���@Quu���Vu"r�3����=pc L@�(izҾ�Դ�n���V,)��v�-�UD=�j�����
DRl������[WW�3��rQhQRIrj��E�~�G�~�k׮d���BMu��PD��B�����+E	�@D�l�%$N��7-=Y��x��*��苃4�ھb��	�뮻�d�b�BU�%%%�z�Okjj�7
"��v�ٞ={R�U�?V����-�DR�y�S��@����;-Cq����Rܠ�����Z�z�켍��� "����ښ��X,���"��n;�۱/UW�{�X]}�
|���4K��+5�)���aȃ���^8�#D���XU��y]]���|�s�K�C帒���c�K55��	9��G(� �i���T�����a�3��64Et�HW��EM]�}�e̅�����s�;�ڵ+ͨ��SMm�5BEă�O��?���μi�2zzz�����i�k�ϟ_�[uͳ��L�[C�#:ћ�V��_��!M����Iu�����'� ��395�Ψ�:HcnO�tm������y vy7n�����X'��H�%�EEh�&%�$�P���� ��:�S���9��������(ߘ=g��k���UJ���1��œk�5��������5z�x{d53EN�y(ˑ0���S�;ҧ�����Y ���2JJJ2���jk�5 JN�\�`���b�(�-�0͞7�ڠ�<��U�>��/[�|=RATRR2Š�~����n��2:X��K��nW��{4y�ԁ��q �Qo|����*��;���,��Jͷ,4��QRrrqJj��Q��b>�H�zc�������vo�=U[�{���vM��2*� Bd5��L�(�)�]<���7��ή�ֿR[[{%�@D����BB_��5͒���'��h���\�75'~�*�Ѷm�.���{����`��Z��"M�5)9�G|/�$0���R �j��/�s	D�iP�D���DI�)���S�#
�+�����L���i���9��E�"������ښ;-��`("��$ і�����Jj?���n�l�ΝJ�f��s��7@D�`�(99�SE��|Dq������Y}Ŭ+�ϻi^�`_��N��ر��}��5u��C�Դ��g)�ז�p�Dh�^Q�!e$L�&�v�("[rrҖ���{�%ٔ�g�QDR+��q´, Q��fmmm�P��f��ԏ�3�ȏuw*@d�_ihh�����)"W ٲ��]�QJr�ӓ�������q���H�z�ܹ��U����Q�R�?�?��R��`���bg��$'5���X%�>hdڡ���AYܢׁ��䏒R��_�����h��6@t���?��n�~{{{���lFl#
�T��qׅ�P�x����+5�7g��]w���[�~����S�%%%Ӫ���u�ս��#)1�T�X>���lf�f�i���NN���(��iA7�
M3L�C�iG��(��Fq�FRS'�F����G��ߟ����E���ϟ����y;�����g D��z :s��0@��D)��pz� #e'
�K!�Z[[��3g�9w��TD�Wcc�Cz�~Uoo/�����t�U���HR���<��B�9#;��n�%<^�a��J�JT��+�5�l��]4�u��:����ƹPF�G���l��TE�;)�I�v�mғx�J��W�e˴C_�?}���6!����o��R��'ŉ:���ٯΎ�8����������F�ʾ�>"�w��
H�j��Ϝ9#;q�,..N����fRJ�C�����K3���q����B�JMm��� �ި|Z�A����<U+�!�;��`B�q1hd2YO�"�LU��HKk�i�#?u�t���ۙ"�3P�II�"�k�!����f �jF��g�)��% ��P�pMu����~6}/�r�W�S]�/
RDDiQ&+�_��/=� ~� ��i����-z�z�aÆ1���x��740��(,zu$F�ONN~/)e��,X�S�bu��G���Sm���ۇc��@�ޤ|GuI��a���Q$�h˖�i��ڇjjjW���1"!�}缉�8"��aÆ������HO}4\v�;a���J��,EV�"�*"�HihaR4�5����noo�5)9�CEZ��.X� ������M*-/����Sw������Q_���=����ѣG��Ń �l����W���� ї�5������GB�c�+�/��&P(=`&9>>~ ##�Ĥi�	�B��;�ܹ3�����z�~ �7uv0d��h�Ƥ�0ZkF�ı��53#㓌���.]S�R:0��":�{������'N�	����͛�]D¿S��P�Fmmi�-�;���W�Y{�M7E��D�4�1֮��t+:::�Q��Ƀ7�~w�ȧF�/�l���̵��Y�D���=��#�VVU^���"1b���܇o�
D�
IiHzk�4(�e�M3v�ؾ���Og��i������֩{�y�믿Z���4�on�K�B ��7#���wC�0�1Sͽ��μ����H�GmO4�����Xt��iV�T�baR_�q�I�]X	*��ߙ�a���DEEE�eG�^���^����� ��<|	ht���`{�������O�UY��"
��?���ޱ���֖'N���I3�B���[�w(0m酀������K±O{ߜ+�|����<x뭷F\>��mO<�/ߠ�j��L��x~RD^Mۻ��\&��d6V���PD0��*���t�Oo	��7�A�� �] U�U��7�F��GD���R�
�B������f�L&�fdd|�Td�d����V�V�2��ݻ'�+ٳ��ɓk���Q���,�a`�Y�+ a�?1s�G��(������7�����}���\�634D���z�~��l	�����R���q�F(u��:����T9�������?�+z��Owf��+_���f����i��&xD �sA�)>000����QJZ�����J���p�t�]mmm�G�zŇ]��<�!���4�J�"��w;y�uVn��s��� 2�˺����҄���w�6O����_rV�^q�쬬wU
��E}DRk��㊋��Z�˵uu��4 <D(�Z���LBU�[�m6���Y��{뭷6yy�C�p̚��|�#mm��&�)�j�@}ȇA�AX����hPϘ�z���#UU�h�W��{{{G��=?k�i���6�_�0�0	ՙ����J��e��Fzm�y��`�@��~�����0���i&v�%!��	�}��l:}�mU{{;���ج�X=�k�H��liiPj�o͙1��pys{ӿ?���u�u�z�Ҿ��xW�b��R���=�N���+3#�lu��� �ż8V"Z}/\�!�4^Z�3���V�զHM��"Cq$*����>r�����2Hy�r�t�&4R��l��۳�g=��f Qmu�z�Ѹ���7�h��]9�9�ڧ��*��+%F�����V)�.Y�Nm۶-�Z_�J]}�<8<�*">��ӛEl��y���100`KMQ�'=+2A��dj_������B�x�?��ci��n����l��Y��"r����P�^o40E�n���zꫮ�ϻ,�Ym���edf�����@�Y����P�DX�
D�̚����^m6E����H0�	Ѿ�{6�>ݶ�WD���}p�pp�ߤ�����߰4 �9���̀�.>�d��:�v�D#'N����>�*���?O���7qK< ���3FA�M�yq,@��������;"�M�o^��H1ͨ��k�-s����g��$\R+H�V��<�P���b�Z���v2͚��;���a3`��)���}U�n]mMͲ�����'O>'w��[��kб�oL�;֚ɲ�3�LKO{(
"_jS�90�z�����ADS�(B*�����C�jLߧC���d0}D�DN{�VL�ؽo����"Q�A���b�Ѩ�ɝ]6�S]��D�Z��555+B���7T
�CQ�7-�ű[��(��ʗ�s"�(�W8�p�Dd�Ǔ��0%j�Z��.-=���	"/�J� ��=�7����<s����Ls�LNY�9�g��z(��Xkf���f RE���w�B�6
"�����nݪ��/564\)
m'DSͼ�Hh~	��\�㤮(Z�k����i
���
���%ٔԚ-))�ppo�����5�0}��j���Uy~�f������G*��Z�C555+C�쬬�2��k���RG���1i�/544^��	��ۭ"�V��TL��J;��y�i����OOK�W�*��6h ��ݥ�;�g�YM ��<1r�(��#:D��~���z�=�`�(++�oYʌ��/.��"�V�RcC#SD�*����f�K��Ԑ+��� 6J���܌���L�P�"�hr ����c4�H�iPy9Ї��nA�`�y�p��BgufV�_���a��wX�H[�{��Ѯ�܁���(4,?���i�4�J555D}����T���2At`ׁu�Ύ5f�y4�*A� D�G�W��p���x?�#�2<X][�*Ԧ@����.\�΄��lْ��2���XõBю�i&�8B8�`��q����wթ��%��AS\\<���C�;-f�fL��
i"x�l˖-�j�5EA�'�%��:��΂���!g�7 �Q��4�����T)�F"�J��_��i�QWW�h�����Ό .4|6�N#knn�"z7/B� �:c�յ5�Q�h��\��H�,+;�/��룊�3}:�qD�N�,t J;+;�H��c�֭��8��ZKg��@$4ciF��Y��F�n���^w�u�� �Á�����Q"~	?�TE�p�a����[�Rn��ScC��d��D=��oe��ֆK�J%=@�����;;-����<k%r��f99���)| � 
�@Tm�}���vuOO�(�3���Uр�(+��Դ����*�@TTT������������(#���̴���r�)��<�c����,�N�h�+ӌeat1��'�l���sg>�?a�#�7���G%��Ԯ��kX���3 �M3�nD��� �@T�Cd�wC
������7�3�#D{������[	�ݩx�SD�O��d��F�Xcc�}}}#D��2WRDٙY����l�v���O?M�k/644�9���F��]8����3^OQ$���۾d�� Ѯ�K���+������{��f�*�|�Tc�y��ر�`�Q�[�A�LU��w˼�P�a"�x1�/644�������f֬+##������ :���_�� ѯ����"� �H�n3�PDYY�/�R�7DA�w��� �j}���5��32�����1A������;�;O9v����D*��ssg�2���?������j@��ռ�:� ��efg[VV�+Q	B(�m�R]����������c������eP&V�c�G___WFf�k�)ɏD"�v�����y���<�"���YP�X$W��ZZZlJM�?��͍H}���DC����Ǐ߁���z	g�X��?�͖x D�X��(��� V4��U��~ DB�x�xw!���������>�i����<&T�H�Qn�-���7�Q�x����?�I�6�>v��W{{������B� �@������B���c��K��Q��� g���yogg�Z����?�ϜI�7�N[�+5����F$����i�5��}}��E	� �����:�"��	�e]4ι6�;����t��"�G���N6}o�(ٸq��yr��iFp���M3�湳���n�����C���7|����h���{{{G�Ze)3��>,fx�D��r����c��?��h�1�    IDAT�&蛏�;E����wv��X��"B�JQDb�#��@����<gFd���?�̠���t�8������!A������g �Dd`6B,y�?�Yzz��G�������,�1X��4 ނ����7Qgu���]����y�#z�������m<�uvzUD�$
;m�p�e�5�gya�`S9Db[������7#1�z�֭��{`m���G"("|<�H���..}D9��wEn����*��6o�dʱ:݆�������Jefe�����5͂d�s ��l6�Rb4�#ru~��;3=�ʹ��u��� B�X�ż��'�H���G�;�U9�������_�U��̠� Ѻ����
1���2_N�H�p�7��
���a��*���;v����N'�x�(�y���D��)�C��.H�����E�� �s`��l^c�XF�vB�r�������xE���0k����w^a��"D����6�mj:� B@��8���6p��Z�T�|Lf������ã ��>�u�֩U�?D|�қ��� JKO3+;#�24�-ٳ�l6�j�g�>(�3�g�^{�>u�!|҇~8Y�5���D��K1�O�9�ς(�崌Ԩ"
V��iF��b��b�|D�l��򽸺'4"o��[[��Goo/"����ʌ���D;�>b��X-Q��Q�YE���9�� 2�k�o�"C�H�N�UC(�Oũ(;;�ϊt�ƨi�,(�)��g�}����%.X B������%+;�le�#�ҸR����6�� Q�s�W1���r���@��Q}xE^�O�禛��R�P>�)"�������/����F�1���UD��炨+��h�j�F��&����ȡJ+�	DV�լR)_R稟�7o�)���K>.�����M��3�B"��������~�1����D���_7����7�fؼ�W�A���R3Rׅ�K3�� QEy�3_��;;;�h֌7�(��� B����l�Ł��3��ٜ�9�^y��������44Q�g���+C"�F�%�0��D�H�gByv��lĈx[�2��TE��(��I�g� �M�@��� ���9avg``�='G�L�̜�>���|�"z��yf@4j�h�%_|��ͻ�?Z�4�(?-�3��믿���k��yӌWD����b�i����Ç۲�������-��K<�W��#9�G4�|D�����;Y���3r"D��l��s��͝�-�H~�^z˸?�B9�"O�j_�ZD����W� �F%���'�Lіk�9���l-�A"�7$��%�k���ah֌n>��'O®g�Yrj�n�q����mٲe������0/���r	"M	�X��77L^e��������6ofqD뛚������ɝ~M�;�Mf����G��"D6�M.�ˡ������N���x���	�nA���� Q�J�|65-��HQQQѤ�%{��i^����JEA��0�Z�ZC����M����F����e:������g*�����&�"c��M���yAI�-�Dϥ��?� �]G�yaD����� �}ͣǛ�����DN�0�J�H����LU��y��󥴕��8��?>�j�5�|� �b�����Y�R?���x��k�m��Ƈ�	��œ���}G������CYU��y��/k��?��Դ���d0|D�u��� R*����Q��]�A��f���j����OE(����4/���J�fh�Ι5��kn��>X}f��ݼy��uƺ'�Z��<?+��b0��J�z5#+}]T	kڻ��v�A�8"�'��FRD4;#��8k�1׵�:BED� r8��Q�)}ҫ2K>)���ޝ�t�ͷGA�Uչ=���ߟfl�~����~��P(@�R���(M)&�>��75���΅��2�<�f�"V9@��y~WWװP*"u��hv��{#Q���H��m�}sK�m�}��"ad��"�G� R�T��g���V��v��B�����Cl�����G���	D��#�J��x�l�m0@4+�}7�xc��A&n޼9��X�Lss����,��gIxfDj��崬�ނH�e�rH�h��Z�皚�o���c�:����g!� �������|D6��C�V=�����{��WWP���B$z`׾�:���D��m�y��D������him��j���|���?�@�O����(��+,��'�%�r���`>}p���������	�ym�I`�X@�:G�}V��{"D���?��k�s�(6
"��v�ȱ3��MǏ�ј1c��Y���"�J�Ez�3��#
���۵�N���>�H݁(�0��n��VB1au�D�/��6�h�Z� r�za	"���BsSk\�f� �Z�����(��÷�onN�i��cKk�w�VkL(�R���Y���\jX�Ƞ��csSӭ��2�lg�*ͳ�i���l0A���)�/Ȼ'�;？�XW�bKk�V�UQ��fz��Ŗ���Aa�(">1L���f2��Z�L�"�P�f��'���'v�{ｗZ[S��֖�k� r_ǡQD��R���|��J�ǖ��[���b� �Zs����pb>�HVD��ڬ�m��ssK�5XJE�5��)�9 �i�/675�E��ja��`)"�J�tjZ�󑦈��w�͈#�~�LB�F��Zڛ��w��v����斖�DJ���陊��8"	�ӗCD-�-0�b`��is���{��J�~J��{!A4���#u����K�����������/zu�+˗�����)U�/�g�o����Z9 �W�_jna �D6�\��h��?}���v�Z���ܙ/D\��OJ��ڻ��3�N�5��Hh���挚ƚW[ZZ�1�l�l�)�9�^sMa4Ul0Xā�Y���֮R�?+o�#D,Ȏ]�֢�ܼY�Gb@�ﾛ�P��ז��+Bl�(U�/�5���Ν�r:X ��(䦙�֮Vi�����R$�h��Ϟ2�;��(�$@����˪5ֽ�z�u6@�R�	�i֟��|N��z⪫�j�����̚��Gd��4��3f��S��ȑ*����~nrVR8;�'�����oo�n���{��,�Ƭ�D�j˷�������O��%�.\rg�%�0}��҂�� ��ξ����L*��	�Z��y��}�*C�,$�/ݳ��fs'rV�4y�jF�Gy��~�������ʺc���8q" �"BWw�!��!�z�J��sf���=;<6zK9L3��Dmj��	�F�r����}v`����]]���b��r�f����r���7N�h�1��T*哚�� ��n�ά�$EԦRi~���~%�@T\\<~ώ];���]]]c�^}/��EL3�*G��3y����RB1auQcݛ'N����?E�ޤ��E����R�6+ᧈ6|��F�R뉖[���c0h0�O1D�� �Ֆ�b�漢�~�24�V�T�V��i *))���m;�0�������D�(>����G.���cd��Ƈb����X��'N(5����z��o�����_�]���lii�g5��!W�%�m����УP?��0���{�K�ƖӨב#G��Jկ3��^
��v B���?���[�f3[�4 <�(�1P b��lߨԚG�3S_����;�h����~������LG�/̝��"d��z>�8���pǀiii雑�����܇���&�3υ"j���'O�Ob9ҰaÜ��n]�H%���&�>�#;[�XFvڐr#�Kgv �d�'S�uڧ�[Ztww�Y-��z{{Y�����*�r}^A��s������{*))�ߵ}���3��,�T�':>_�&uJ������ Q�:G�V�����_�	_���-�pw�����ꏽ~����� W�<�)#1H�*�L���6Y�ȑ��lգI)	���K3�@���O������r������ )"���m�X1�vB6��Z�z`����k�eop:����7Ն�7\�i6���ݭ �>��к?��������b�R��r�f�o��횰� ��>�z�-E}]��N��� 2@��{�W��Bӗ�����s��}�|r'@����m*�rSRJ�ߢ �ż8��>�������Ǜ~a�X.�/���|}a������f�L.�Wkf��S?�*�$������ׯ��0w���l�b�ȑ,w����GJ4?�F���Qs�7�3^�B=�y?�g
TE��es'����c_�x��������W���C���T>�H"�E+<��TD��'��Ug�弙��g	�����SD�_�<��G��L��d2Y�2�*�w�y��UL����*���Pe*�{g�Ա=��wB$	�պ���Zk��W��A����ڧպS@E��ZE�즥�CQ�ō��OY]����	Z�-������%�$q�O>P�w��33�9�̙3�}�,�k��gJ��Z����fn�޽"g��ZZ-�"0w)guYyш_��������������مw�m|��R�b��B�H&��Y,��G�#�i��411� ��W���I���	�F03�u��׍3��ĉ�թsO]kp A���ʗ?�� �L���+RY�Ո�A� ml<6|����qQO5VW?7|C�K������3`� &�r:s�B}������ g��'OdO�T]�xa٪U�e2��;���E������>�n�
(..Y�`2lll�ㄐ�I_���N��� 1"T
�~
p/..��X��Q#F~�r���uӫj�������߹S����Ѳ�}�:YZZ2QC���=:[�(@Oq���'UUM�zE�w�{޼y:3!�n=�k�.�k��}bfb:����
d����g���L���+�H�Hꏎ��x�:~�)n�޽����WU=���b������.���'B��Ȭ� }�n+������c=7.\8�Lo�$����m�f{��ͅ}{���21q ' 4 4����А�A��3�u`���Pu%I��UUg���\�cǎlCiXM�9K<�%�^��8����dB��� y>�9 ��|n���������4�S��>K,w�z��ߗ.]����b���������@�ȇzB��G�B�HӇ�����������{��c��a۷o�� D�RE�ACՉ���cW�����Gs���9�_�@�T��9�U`��1��!������p����N̞=ۨ⇔u�����R�th����-s��X�����r�������G�.�>"lċ#NM�2� ���z���V%w��1���x}�D򎕕U?l��������ӗ�Q(��cfn
`gTUU�|����݈#��b�A�4��Zn�t+�V����5ò����hWfw+҄�@��+����}�Z|��W?���錪ܫ/� �����-������D_��g�ep- }��=����￿�<y�w3gάPE.�r͚�k^���A�-���`F_�W������ߑ���H[�3e���8�����:r	{'O�ܚ�C_:���f��ڲe��G取>����߿?��`��Z�ŕ � D��P]])�I�b3dyhh�Ec���'�?�1�a��������������eŲ�`�4�dO���0p��?�_��h���x�޽�EE�o�VW��X�P\h8�����#��C=Y�U}MM���W���j��u��� ������^����j����j`��������\�$�[|{�p.��D�*�%iii}
�^�}��g�ff#�{�j	ģ��t�+hS`6<}�����ʣ/����%Kݩ��6~T��9���?�pРA6���A4A� �_��\C^R�r�w�ޛ�\n����Z}��h@BݰaË�����2��Y/����A����r �?@!g62�@{�U������},�_r{ic@p�s7s����d�y!kyCC��T:�� ZQCZ$ݔ@d�l�J{�2˪���43hf���K�>���g?Vp��3Sӷ͛>T�"ԑ֣�_a!�(�2V�?4hз#G��T��]�<3*A#�ܶ��K�/�g�A/@ ��J4*rd���B>"X%�������dٰm֙���
U+�� �\�q��w߹?(�^^V�2��d����E�����J}V��7�<�1b�F+k��b�� r(�%$5/޿��ӧO_-/��Y��ߣ�#W��Ǌ����%��
��ׯ_��f5��r������q�	�x\��%���  Qs,5�Ì&Yyy9��no��C�CZ�x��m���������Ƶ�~7o�}*�Jy w ��u"��z�$c�kΙ3�r���~>��c�W.e�.))^hccc0�#-�-�O�P���d�nll�n��d�H$�[�hQ�~��j�2:EF~k�����kg�O[6ۄa��FQ42Z�?���������ƿV�֏�Y�պE۫��~u�x�>O[[[�W��R&k��S��lKKK���OS�N���X,6��g���IOO79�v<���[�\�͐!Cڤ]�/��>����ܾ}��Q/�=v��B�Ai,��~;;���l�	="je��v���Fލ�GB���_n(I�5���MIL�-��߲���10H�D� d�!��r-))��K$Iӽ�.���Q��P�2Ftmh��I�����\�=���e"�%Ґ��r.--eܹs�x��1k�]�6��P��W_}549!u���:��a)6.�i �~+eyy7˜�D;fD[�!m�ojL*;&��v�T:��Ʀ�"�D��/�� ��d����{ӦM���[��dgr߸q�k���s8��t�倬��a�,,,�������͛�i[}���@�g�7i)q_s8��8�@��!�4J�����}:�ż���,�U��9�M����a�$�|�`2����Q B�D�uh��`A "%�$����L�b�{�4��M�^��������	iD��z�چ+**bz���nxx�qM��o�'�R���q^�r�m�� |�h`��ՠ�:9�8y���N�8�)�2�0 =o�����9�mgg�j:��F�� *--����%�N�]<E�AD�N�&dg^��Ύ��yѤ��)V1n��ݻ����;�n�?�NC5:�۷O����5�˝��r	����W�h�&�,�xĈᛧN��5Qk�N�N�N<��!����r{�>���iȔ Y����d���IS�OY,��FD���͟M������m=���'�[Ј���绸�,���H� �C	 �����4���F���a�A�8T!@V"n��E�-�����ћ��G��}M0�o�x<Sؚ z�E4h�N�Q�RI=�<�g�b1ֈڌ�����g5��>��rh!�~���Ν;��]��߼y�=�jW�(5�f�����H�E���gL�f��2GGѶ�K�utt��-M#�!66�{$�[&�x���QA� p���;��$Z1������Ɔ�Ɣ@ߙ�4S�����ʼ�����^dkkK9��29�C�3�8�	\RR¸[Xx{��{�ƍ!g����v��-LIJ��Ϸ�`ooO���F�n���i^-*p���/ރW�Z�w|t<?&���9c"��fhW=}S&��! Qyy�T�(K��3�f
�	{;#3s�@ �@����F7����)����`�'��@��=����ޞ��2!M	5p��
�/g~i(Iǻ�bbb��c0r�2�c��iF���D���1���g����������B������R p"�B�E���4�z��5`ӬuC��iD{��%�'}���_VDw*�]���� jb ��؄��+��H����A�^#��������A�f��hD��tD��n���V�����?��)��<�Kt���P45r�"Q4�fDJ���G��;wPSɤ�To?���F�V�a!a�2��v	��iD�;A���1?dc�im�2}��(A��О��GG B�?�`�ycF�    IDAT� T��eМY;�F��ED�1q?0���5҈ei� ���O��ܦTQ6��B¼2���� "�We2��4��H_0���F���o�@�ipT�D�D�5�� �ɤ�cӼ�-^�iD>�YY;���VN�N�;��]D�����QR|ߞ�	���7��1c�}�|UJ[I��ӽ�-� j"�̬�<�#B�����SO����tJJH�����C��) Z5SE#� j߰4�f�.�˥��>~>}||��i��j��������\ p�Dݙ���|D ��Ј��|~���~ %�����gii#?�,���Q�q	 :w��d��f��@�^3�;Z �Y���G ����3f�-���*�����p!@�Q2��~L������A�բ@���#��wSD����������B�4����&fX��=�`2_QD��6�$y���k�X,.зw������ddfn�D��ڭ�u��C��F��#�D(�;rVw����{��H�27��:���)+�"	�����|�;��]X���33�2 Dv�����c���t�5
htwuo�.�oW�2�E#h�����]A#� Ҿ� 1��=�f�Q�t��!t4SI������򵯍�6+#3s[G RLYC7͚"�=燆�7���ֶTD����;"���%��9��G��n*�5iD�p���svuŪ���\��)�;�d2!����5�/E)!�z�y�ņ��+���@�L#B��o��{,� ꊖ�A���'����]}DD�qDM�j
DeB�`���_v�t�z=RD\.����@��a �)��W�;����V����>4tCx`fV�gH#���P�;��n�{�-	�����yw��5,-��O<.���i����� �)�M{�ځH٪��F��8�o����M��4=T������[����~7�j$M JMN�L#	�/g�Ļ�i@�(&�{�1AU�`�/I	�A��C�n���ya�@ {^�6�v��8"���ݻy��և�?��Xѧ���G�"h8�t�+4J���}�Ӏ��D�� ��A�5=UD�4k�G�A���		������"�|Dt ���g�S<

��<�懄���O@Ѵ.�������i����#:T�k��Y����. �;��`N�ry&�Ȕ��HchH��cQ�p��|DD*K�/l҈R��흑��g��hG����	�]�fcћ,::�����Ʉ�h���%��jl�u��C7����̌PG#������p��7���C��ٍë�e�Q+�@rt��#�4�/f��Ʃb[��(.6�;AP ���:�ĥ��C`�Q "%�����Y�vk	��n���bܑF��ߊ ��fw��:88|!�9�ی Q|l·A@��6 ��>*�5��<�+�	���ځ� S�x��٤��25�6z�9�P@���i�irF'�6��_:t�`� ?|�4����;�p�[�`�M�t�2�}Dͦ�Y�>�1�ڎl�efdD��{e����j:�
�A���D��K����3�[Ad�01a����ѝR��a�4�i�'N�W���}%�Ę��&'�!����JKK�$I�i��z۸%��۩
"T*:��Gt���c~H���=U?�6z��=��4"�GQAaA��A��4�)�0�Z;,��P�����X�H#�D��bH����8�����ꬾ{���}�~���4"�߲j�G7��<�AC?�����8`�+�X4L?��MG���� �7�\�rVC9*�f��<�;�wAw�7��|a!as�_8![v���#9��
�^q�p�,C�����V#�Dp�4�j�f���h�j ��&�}� D�1�_1	⟚���4������ ���w]��� #��)!k2����W�уHq�@iD���@��w��-ޝ��ȑ#��k�~Rtt4'>6�+�	D��Ԉ�$�����.N�ֶ�)���Y l���Y>"����f]v�p��~��,��=��� ѳL3���޽� "`V�7...������@t4q�b��	��34�)�E�FU���f��y�qBD ���Faa�%7OЈ����0�t�cQ�����|D�/Ӭ���@�)`V�wD��;��8����X 2WW#j�Y��n�E)nz�_���Ft��݋�.n�ׅ��� �C	(���U4�������������'O�~�ĉ�z�z=R% ѡ��{	��� j���I� �{���G�K���2�2"(��A��A���{�RH��������jE	���I�'� j��?I�Xok"�$O�/��z���٪�iB��4�{�nn��:W�uꩲz�4��k�"�����A����b�X���f�111�#1��,����$���}��f�u%@b���LH±��Q�u"w��u��.f�j[k�Qd�SB\�/C�u�p8ԆWd��y��|�\�h�ѣG��'
�nڲ�&�)������uDGcb�M �P�G�H�t�# D�99[�|>��ں%?2������.~� ���#xu��K��Uϔft ڷk߰����5�P X�y��_D��g���$��g���}Q7Z���+����윜�|>߮#!�2�z��[�n�e-��7�5��\n��ժhD������� j������j�ՓW�6�m������ωSу��<\��D]�H`� �M���A����DB��1ͺi$i	"X5�f�����c�5��9��D����+ӈ�ę�d{���[����Л[�D]IQeRܵk߰�ĸ_�k"�@�v����#��M+�pE�����-++� R�~r����qvvv���L3��� %ſ������=��^�A���C�����3<!.�gM@T\Rr_(�����3Q�|�������Ad�fڂH$�ۼu�ODF"=u���?�����YU����F��:P�J��b���4Ո�WufB�4�w4�#�>��G-g�_������Ϸ�U�4C1o�����$���u.6��J���'������$A���v���`~ee%���쾣H�~̸1?�F����=�(���y��7v"xʩ�b��_TQQ�())�quw� �Q{輘�ۿu�x��|�X"݈kD��#����t�3�g����k����g7Ϲ�W/ǫf�o�K�D�!��Q�0�(jD�"6��}DX#Ҿ7v\���������:*m�E���H�U�._����TV�έ;_L;�eo?�҈�x�A��F�q�i6��q]��p쬦	kD���YYY�I�I�9��a|>�F���n�!��jT_-)��t�kD�o]��	�@#��fM>"���"���A���X,��EC �ĸ���sB;]#��D�%�nn�W�\y��a�ѱ���Ǩ��t� �����B�#�Bώ�����M�$Bcg5Q[��
"�VԈJ��r���1{�ʏ0����۷o}���( ��k���������`�=zT�(/�A��Q)��C�X�5]�� j+�k׮�����9����ш�2�h��3���r=]܃��^~Mǡ�u2:�HDh����AԤ9�Dk�7��-���D<��e˖U�8�F�$Ӽ}��ǦY�PD�~�Y�{1'D#Ӭ�,�kD����G ���c�����@_�F58�����cF�#�Zi���}l�$m5"��2��Y����5==}�+�L������\7Ol�������۷�}�Xj�� ::�޴)��M�͂� �}o��ܝݰi����M�t��|*�iDp���4�"G�hu����;1����fg�n� �<�G�`2!�ͦW�)׈�M3�4����n��A˗c�nȡ�Rvm�5:���(�;@D?`4"� N`������#�
������0����� "��3O�>�H��m���|D����3pŊ��h7:g5��؉cQ�r!�-�*�H$~�9������D�A����)�`2feee���G�R@ԓ}GU��h�޹s���ND�x���|�L3pJ�5"�R��4�� "$@ChDU[��0�4�\���"���+��ʊ
H��
�t_{ݗh ��@t2�d�ǥ�x@�|"�j�R*@���ay�=�H�"|s�!݋�pK�DI��,���i��4Z5�@TY������K�i��#k��=/�HK��*���FH#����@����q���z�r=T)-A�@J$iDmO{=�uuw��lٲ�=�-t��nՈ���ѩ3�G�X[S�� d�)�҈�<y¨�xxW���ѧ���ө��0-��1���Az����~7''{=��2d�ja���nC�L�&R�$0i>}�4g��1�Dz:��m�6����~�eێF���U> ����BG��u��K��3� G�`����,b)�LYYY����^�����[����1cGcu�@U�9[���������v R<��F3�H(\�v��du�k�׫���"9C&�S>9���p�Yj�f�VN:���K���>��ʕ���������X�A_}Z��H�m���@#:���A}����ӧ��ʊB��9�
��D�H��Q�HP� �v� ]�zm��[<�vz_�D.�˖-�>"M���ٱuǘ��N�`cc۲���ظ@�1LFuu�"�֭[��43��d��FԪ]*��$���K|||�F��H`��M|����`�Q�&�i�pʻQuuu���D]��-��m_�M?{� 8���h�8�Z����MQ�]�@���k���1ݯ����]w���?-��[|������V��q�c�򽞎4J#�����P �p통�^��z*S-AD�$��5��� JM>�ޕ+� D��ZQ#� ���J��m�b�f�EV+jDPҊ���*�9
EKW�_���i��2��$%�?��i�*T QJұE׮]^��_5C���R��f5�5�cǹ.]��k�
���4;��vvv��lvKFFz/E�����񤪪h�СK�nX�������D�~�K�b�}~��Z��t��d��]h��D���=`�u�%Э���Ъ�����i��<-8`)��� ��d����D��MOO�<u������JX5�L�A�u#XG �:R����"U�F����"�@�5"�k	"	I��޾^b�
�ܹs}S�R>�q#�c�7@���ªYhD�Fկ��T`W_�	� HMM|�DB�Gk֯9���4��tVc)i�����K�K�w^��e "++�vѳ@�<f|��?����q0=Dhe9�A#�/�f55�E�"��UkWaQ{g���	IH�$) 0��iӦ�c��:�F�����7�Q�x@5"��h9��*����!�DB��������q��5+�FD�7��z$&6�E���*V��A�?����P�˚@tli^ލ\.��L����ks@c��+[�+˦5�* �;��a!�)�����H� ���>|t/�b����*��d��Y�K�F��Y��ƍ��0x��NM��D*�\�/�D�f}�>�e4=p6l�U+���{vg��5��X�/"�HV�NO�0/��'�Ҁ����F��h);��w������8"�GDh�����4gu]]]����ҕ�Wѷ��=)Ը_��%�Aoq�\35Ӏ`�HI�5/߃i����P�GD��i#,d5`PfL��Wk�jsǿ8;�{r`t��-[>w>�繃����������i?A$rrZ�jՊ��\�V)GGGs���L�?�\��� ����=@�~2��W<Dha�3D�������Ñ� �nr��A�-�[\��q� ��igg�NR�j���uuu%"'��+1�̦�i�à@�A��� D��#��\5�x|��:-��Gyy�D�;ӈATWWǐH�,�1�f/\����1J�����l;�DPOe40}լ���T$}����'6e��FLL�HL�,�x��嚨���פ�Y�`gukgjѲ���s8�~��i�`�5�d�8�q�.� ��!�٦���������(���l"�^3���2'GǕ�����\\\��{�R����'�|G�k\.��A�}#@@crb��7�/�p8};��gAs�/����1k̸�A�-��}mz����޲e��?3 g���M�t�� Z��?_����s�%�|�"������͜�kD�2�$�||���e��� �` ��Xl��<C�� 4"0�� �,1Rw��ƺ��a���'O���ȑ#I}}��Wtt4?>6� A�r�\BM���'���m[MU����N���644d�s�M���>/"<��BV�A���p�i�Q:����:9:��������Q��3��:"ݷp�i��ƍ�Yvd�A*c�Nj�Q�F�l�1γ�����t�<ڗ�u!����M��" �HUؿC[5{��(Z����A�*5 QBl�A&AL�H#"�o_�����V�?~���3�����7�Ͷ4hPK�FЀ��Ň�C�S�(�qv�A�=5����6}�q!3〪 g5��&%��G��^^S� j"�L3�v=��el6�D�dh���~:�d2Y�x�qD]����3;��kk�a�4�L#j��)544�;�D+��כ�a��@���f�/��j�Qg j3&���J�R"���
A ����f�r�����F ͨ�QZ��(���7_�� RQ����U3u�Ս�L�9��=�� ���+o��\f�f�8p`���ʆZ1�>+��rǹ�bQ�D�b�n���̌�6��N�@�b� B(���(�J�D����:ֈh�@[��8"�ADJ$���4����k�=[n�L[��h�ܹ81�n�D�� ��3s�4�@�x����4��Z*�V���V����_�F��.Z�H
�xh
"���)-==}��N��y�&�f�҈��0q���.n�A�gϾ�?o�yM�.�Q]�� $9C^!rt\���oag��F�Ed��5���Z�ݪ�q�F ���?�T�l6�\������n
fD rsv�8/����_��>uS?��������C;ӈ�4C>"j9T*�Y��Q$Z���w~rpp�ןf�ٚh��C&!�T_�w�Q��@�O?{�����O��˻��2!M�~:1���"�%gW��s�̼���Dy��nz; QvN��!�֎����A���z@C#5��=��VO�6�G�������4�y�M_�A�*S ѩ�������������FDҌ �v @�e�K�_7'h~ХnZ]��Ѷm/gedomm-� D�N��kߙ�N�R��{u��2�$����]�Ozm�izz���~�p���l6�@������7�f0]��X"���d���L]dE�|��dde~�
���J��@m��tr����oc�n�L����0�Z�z��	����[n�ɟ�f�	��i?���D #�����	
���X�˂�m�6!+#�[U@�E	��99��4�f�6�����76�;VSu5"9)i8�?K�`���E�lkC.�X�1��N�*�s�o�\3E������pq��sfb�~v��[�������"�P��N|��f��Æa)4mӦW��$yr���D��MHH��=s.2�v�t�À�^;�cw)��I�\Ǝ���oP>��,��m߲������� _X�`2�Ç[�5��$�������=��W)i8��7=X,�����k����=�~f�۷�r��6QG�A��5��`�͚5�b��^�O4F�����kk!�Y�L#�Y��<��i���u"�<�7�7����a�����K?�y;?*hD�4�V��Ȏ��q�&M�'�uչI#�1L	���сh�������܋@�� �ln�yF��x8|���o��6�Dk���+ D�N����ϟ�4"j�L1z��*��5�� D��0��P�"�M����c5d� ��W	��  �IDATBh��$S(���Ąj���jJ#2a�ʇ�ɛo���>��|�Q���M ��^ΐO������}!
�e�F���`�TVV�����^^�z�ez�JIII�gO���u��d�GiDD�$~h�>�1B��T�%�5Ww�y����=�:~�QiDr�����ϧd���b5�mۺ���� A���ۦ��jk!08ˆ99������������ѱ��g0����S����������͕���I�᤿�x!Q�P���Μ>�UaAZ�DH+���)ȕ�A\sus��b�3*%''���s�7�R��!VV\��t0��������Pkd��T���oOO�#8y~����_y	q�߲X��9�O�>- ��~�7�%����d��ԥ�X4u�T�nkґ$����������@s�8"��"��|P�	Ȝe����e��Y�fe�X9��
Diii}r2s�.]�beeŶ���@_40 B����ߠ�����2���0����,Jd2���G��k,�XJ�~&A�ammm
�C3v�&��-PB�/������Չb�%S�Ly�#�\z�H���P\\<��Z��F�:��wІ`�0���^u���M3�k���������ܜ���<x0H���)��¢e�A�4���i���/��ᇋO�"�[��a�bbb�G������X��@�03���yY� ߿������1^����ǧD�*�m������Q���ib��Eࡃ�Ji@,f b�X�>}�d�w�����*����4*��?y�dPfv���}������� &I�,�DB������4 fffd�~�.�=rɇ~h+�������PHU�_����}`�4˚��T*����ߧ���3&��<k�c]����9p����Y��߾u������L�1	�Twd��jjj���[9pРnc\B���c負�kcx	�;DFFz^�xe��Eo�EoҔł�"�44�7�,S���	!�6Z�d�d�y��QާO����	�Ż�����[��y����ƆF7�`0111ihhh�?L�((#�� 8��Q*�J�RY�	�86x��C�|�I���5m��~1�⌢{Es��z61a�0	��"X�� ��B�2��A*ml411������%d�`����ρwI,�5�C.cm�H�{�DiQi}�ܻbe������Bbj*�Àill4�J�f�9Sn*'�R�L.��kh 1�R���}�{�����_
�J;��ݰP]]mSYV)�����f�&��!�ɩ>$')�I�&L�D�`J��Z����ή��ۻ��D{�袅����KJ*��X�@�ϙ0&L�ɤ�[�I4J��F)S�hnn.%kHyccc�צ�����&M2����D�vy��Ȟ��rvv�b �&����&G�����O�}k��_�V:��Rx����x>%�=���o�%�%�+	`�J��,,�%�A�����XX�� ��$�����XD�߈%�%�+	`�J��\�����u3��jܪXX�'�^�uy����"�P� Qw	������0����K`	�0���p�H ����-0���p���E��V� �&����LD�`	`	����3�[FM    IEND�B`�PK
     C"BYW�����  ��  /   images/a3b4885c-2487-4906-a080-ee9b44acb175.png�PNG

   IHDR  "  H   �9�   	pHYs  �  ��+  �sIDATx��y�,�Y'xr���/������Ւ,��6���܌����G������@�GÄ�艠���L�0x��� ��`dO#ch��� /¶֧�iyz�z�]�֒�s~'������Zneeee��T���2�9y��|���-
(P`�(������/O�
"*0a	�6(
"*0��<ϐ�I
M��[�`$T 	D4q(�\�� �
�(P`�(��@�#GAD���=�(���X� �|� �
�(P`�(��@(,8CAD@>Hh�����
P���"��QY�9�38�@�IB�٦ODgϞ�=w���g�n������5͍���׮�������/��.¨�|�r]��ѐ�ˢi�M�i7]|g���8�iY��w|��x��թ����c��T��k
�i�OCû�,��a���(���=�u�Ɏ����ڪ\+,�-��͓m�m{~�1�m��^p~��C��rvi��t�^�Gu��Յ��vl=�����zDէS�z�;ť��9����^�X�W���>ZrK�k��]u6~�fC������}�U������ˮ�{�q�qՔ�����(�*I�����o<���_��g��lD�����p��lǋvɾ$�o�V���,�5dK+I�)_�!��+��0 Ieyj)�ε���ܶ�!�?�|g�!�һ���4�\zF�u�AW�`�ǿ�ɧ�ʡ�'��Q�Ne�j�^��q���~v/����Y��9����V����<'7|y}�E�C��<���uC�Q�B@�B/��ο^�7����;r�I.�=�3K��lK8���ɓ��T���4)05"��ٹ����akc��/^w��I133S������g��h6n����^^�"�����0�wC{�}ʠ~�F*F�j4�ǅ�j��������S/۶ݍ���F�yfs}��w��W���w��a@�]jD455���/��{��ջ7��������RI��u!EB���hJ %��Bؚ}���R �$� �Xӻi0QC3�٩Mmom7��.��Z�����!"��f��s<�U))n�3 dD/��gP(���㛂�va��^ ��1ޤ$���������\�TK���ZH��*Fe�6�s��ԕJ�"��2$�6"j�>�����@��"���"Q��D���q�q�1)�ϛ�I����;��R+��QyTC=#��FI�0H�"b#d�B��1	� ��h��1HG�Ӕ5�N��Ѷ��fZfE���e�<�#��V�����T8�p��ɨ�
�'0 a:��O���0� U"��[�y䑚�:UT:�����b�I��i�~W��d�0v��ȱ��;ٱ%��Ʃ;N��TD��""�@qЉ*�~�/0�(H�w���Ɲ/���D���OH��s�D���b�Hi/R�n/P`R�5%m��y#���YV�"����3���&��i������b�DF��qK��ܩ�J�:Y���,���m'�(��d�E���4�D��x(H(Mtyx�⩈q`D,*F���)[�A%Q`$H��U�%	i�2���2V��Sx��l�}(	ϖ~����q_#-�4R�8���aXX�%"�N��P���9�2E������.V='�me�zS�=Z�G�yG��f������:W?�����c[��gCF�4CA/uս���4!�1"��(�s~/���Gg�f��}�AO/ݮk+m��)�5~^�D�فp��� �l�W���^l|�BB� uE#�iF5�o��\�@u_}V��X�&�.�{�\[��h���KB�ϻH11������hy]�ҥ���~�I�#�i�]"���t�V�Ƒ����=��d55���t\?�H�H�K5��F�����\��^R���g^����]�#�zy��!���.t�'�c��;�t�N�t�
IhggG���7M���[H�I��t�7�I��4v�\6gffԚB"Z�5�D|\*�R��8�IL#0�ē�����u��FG�Dd:f��n��C�'��h���ٸ�B�#a��{k�ʕU���;רն׭Y�Y������B4�/�2|ջ$/[.���r��_���}��l��KE\]�pdjD�(5��[j���ԉ�_W�ZtL�a:}��t@<���V���F��]��Vg��w�w|ef���|i~UL�)�4��)�x�|u��V��.o��is��cL5��-ól�nK�jj{m{i���έ��Omnlܶ���Oާ"��iJʅt0$19�;��?��P{E&�!��!��W"
vM0[�w�
	%=,Ba�C���޾���y|mm�%��=������/?y��^�Ї>�1`̿��_����W����~gug�G�M�Z�d��:�MRJZ���U5�թnY�+9 ! ���\/�ǖ/�l Q��({�n���̓g����Qu�γf�v�f<���o�[�C���\��lmmm���]����������cR:Y��_��ͤ<��4j��Gy�����W�k���������|����K��f)%-�AF�� ���G�~�g��lj�l"*fK�4zmX��:��JD0l~�k_�D��jYw����5l�	��ă��2eD�������!�A��0Ѓ�+WVW_Y�r�%�4�fi�U_�������b�_��_����ދ���̃���J嵿;���_^_[��r�r�����(s �<�'�{B�M%�up�}��z0jp}ts��}��_�<lU&Z1
z'=���	�}.�"���:� �	��s޶�o���;>3;;����7�&F��|�g����C?y��._\��,�'_��ˠ��Q�Q��8��&Qh^C=�=�~̮�y��_����ӧOC޷�:Ahu��ܞ|��s�=�s���,�����5$x�vd�_����g���w����PvDp�}�]�d�&�z���?R��>(���5E�L��얄�>c��Uv>Q�1l��{�~�HQ�&�>���S%���S4�=K<p.Z�M�����O�Sw�X��-�iԈ�$y=��L�u�4�Y\���k�\�׿��q�w~Gd
�� �������K�.=����q���K�	d���H�L(�Rv�K�$�Nqs���g�],)����1�Ża�*�J>������,�C�Tq��T�6�����GFF�gV"!��N� �M���R���p������5�a|�#����?z�c�_[�__���>۶V���^T?r:��ҳ�f���KA�d�#ӓ "�
蚆ٔ*q>%"?�����r�AXI0~�d3�5Ge_��Ȩ-�N���X���ժ0L�Bɲ�v����9r�ȓRꨊ1�?��m��=])W�������Ӳ�W�ϐ�<��n��2��%�L ĩgz�yR6U��1	�u=��f#���*�j5WVFQ,P�°��ywS���02(Q�( "�`�������]���[n��9�=!Ih$�B��֋���g?��˯5d�N���}�l�xF�>�()��M�+��������2�s�J���:�ao�-�.R%�n��q�ܹuW8g6�7�1m�D���g�b������=��6n�^��MH�$LG�NX\�%8���MD�E�3d�^�LU�a~z�?��ȓ��GǊ�A,�K_�O_�Ա�/ϭ����T���/;w��:L�Y/;7;pW<����/�@M*��l8�]�7`�H�T> m����t]g�V��KFS��T�F�Gy�l쇤�P�p���3ۑ�T��K]�J`�G�tۖݩ��<��;�׮��w�m6���|���V���_�C���������y����%�Lg���(�G��D�c�A%�]�(�J�pp�ʿ���[���?�	�� ���k_;u���]�xq�f���C�d����'�aN$��NR5��x�\�"$��ͭ���z��i�R�l˺�!aX�z�Tw��i�J7�4m�J���[DI��	ƛ�3�(46��l4�3\㑻�{��v0��_S�����{/~�s���;��{�����Ҝ��6�S˵=����5,�ёM��m��\lG$�l�T<���˦�065%Ӏ=\�l��f�}�
6,�r�N�1}��\�p�%!�-g�
7|r.�.!R�ЉI�k�k���g�f����[�w߇��9 !e�yA>�O�^�� '���F����	_{%�a���Ɵ'�!	U��K���f��5S��>7;װ�*X \i�jKM����a�؁y �۔s���m�-t)[��SC��A��0帑�H]Ķ1��<��Yw�U�q�M׿��^��H $��pV��}衇��n�I���������~I�19۷� )�z��Loccû�{�^�����?���w�Po6~X�""��Q���ձ%?C�'�P��+�����{�����ӌ6.��f�o��o��o}��O�>�"���4���נG��s�%%*O��Ls�s�\s���x����� �AI�>�lIJLJ��ғ+ǅ�������;~�xs0V�0��[@�$�����c��cL=zԁ]N� #!"BP�T�曯�����T�J��Lv2
F�F�&�8+�m�Kv��A��kWV����o|�c��U�C��}�[��g?��W�<,�d�x+�
��pz��^��`��w���k��k����]9�H�hԐ3��Ey��t;Q�mE��D}��Dc���+K���7�t^�����~�?:}���.^�����KJ����^�A:�G8���:r�$��)`�4��YyL0�D$EZ)����Ab<ͪz�X(v���|�@Ґĥr���쾗�������\����lm�z�$�#�A2�m��ЋnD�ɛ��~���=��
�L3Y}�0�D4��X�F����9���m	IE{�`<J�KE�J0��/�۷ߟ�ˍb�I��ԧ��z=��(��"���t��MB����%���%�Z�&��+���`�8�>mD�O��5�����_�ʍW����o�U�!¾}��///S��[�\�rB0�^D�3Z���vz�E��ǻ�`�}��ۮx�LÐ�5S�9#K�X"���*���^-��;�#�����nll?|���I�$&��G�|���+��l����e[d���:A���t��v��>��u���[q�{3�� 3MD�jpp��|�:�{|fj&�^�n���O���K��>�����������z:���u0l'�ݱ��&���c��s;3Vo�[�������+=�����>����i�&���A�$�E׻/*���{�g��i$�<��X"��"�eZ"2�����^�j��l����>z���D��8sٴ�3�}����n��8�����A�����a�n��3��%"9�3M@�#� ��LQ���ǖ��J��Y@ڳz�\�V�S�%Y�H�h5yP������y�Ƣke
KD�7��=@�р��W�*����\s S�Pڪ�������³R��nnn�#�/"m�L��O&���I灖���˜5Ox�OOO���5���g�}v{i߾omm���V�!Q&G�EH*���)r�LA���Ѵ�'<1_U� ��T7�}�{���S#�'>�	���OU����|���h;"}��pT�e��Ɩ���eZ��[J��DNs�\.�DBy��W/o\�0��z���Z���������%�I��t"b�{��tjr��e�Ť����937�㺗]�[ًaZa�>+�Xk�R|���ܥRx��J���q�)_���>�ϬJb�dY&2r{"��)C-�v"J)>�n�y���$šH���fgg�*�ҦeY�.��v��Eu¸�\M��ThlU�A�Vܑ=�AnL��)�O�d7�.@P�T*�aZ5�'w�p���Ҿ�\��勵�ѓ�l�9��DK��aLD���R]m���T)��/~�c"�%��%"$�7���Lwڸś�ɡlۍR�p��#ۇ��Mr�!��,�\YY)��@���(�.iW�ŉ?�Li��m�Pj��l�����Q�J	�G]�QX�&���e �k�����>n�n��;e�M��ڦe"�ohk�Br��``-/6�<߉%"��+��-��	�Ѱ�������y)&b�/�'���=Ca�����s!�XL�јX"r�ie}G|*Sa��W)���>C�w�����ӜÚ:=+@$�oF���Ǯ9@u��Dwb_��6:�薔�f��S�m��6�����r�9EE��r���p���Ʉgda"숸��rY�i-��6?��g�uZx����R��dۋ�7����.�1i��`��h�W���pK�����N��ѣG�w�yg���hh\<��\���Ω�%ڭ/�X�K���y��fF
�>&������{�|a�����S}�/��myx�v���M���'����7bw�K7�{@�30�U�Ռt8�X"b���x�li�J��r�-���w�={�"���	H���/|a���'�i��}�zd$�e����gbJO=�\���sꄉ%"�������`֟��2��{����w=���g���#��"��6Vo_^Z��T*md=�m(���L�occ#��+
9!���-HDj���m�(fy����������˗.�o�ʾoȯ&2IZ�ј�nW�Y�_�"#5���hy���uýp�B�V"B�STN���'�83��5�qHZY���>w���7^�p��xJL $A�X�}H�PI7�{ޘ<^%��/��/��"��	���~
,��#n��<=���zfZ�uM�Y������o�)��P0�Y�k_����~���J��j��dG�d�*ǁ���B�DR�X"R�j�_��Ӏ��1??�_*$w��������(�A���<}dk��ϧ��P�jZ슶���p*�{H��&���ͦ��� *���a�-,,�����^z�7~���=���7D΁�?�����'~FJB����(����10W2Q��hґQJ�Z�ʏ�`I`ss�ȩS'~qښ~^t��ɝ���z�����9 ���ICA��1���Ҁ��&���;�9�qL���|�F�5H�ͺ����=�����ω�Vv*6 ��G���̷�4$�T	dڵ�4�������f?�	k�fD4I��AC���6/�BF�:7ʇ�=HEr��f�Hu��Ӈ:*�>�;f$Nn���Qw~R��AZ[F�Ժ�@;Dy�F��������hqDHD��Ğ`^(i9��8B�3B5������{��跿��/��>��m�����W�����S��yaaAIC #��E���\y�H��O��n��{�JҘX"���r+�Jc}cS�NF�T+�ڻ��I�"����ŋo��c���kW�6y�o`�/�#<���}��w�;w�g%]�������t		Ȋ��[���M׬��M��ݝ��c2�ȊJ�ԑAT�����A������mlm~���^:!OyQ��X�^<���뛿^*��,�j��,*	���,�I��H��.���ً�db�ȸb�LӰ��^}N^Sf�؏=B/�N���P�V�R���Ç�ɿ��'�Y�w�׿��o��ocIB��'��q�����T.�KJBS8��x	%*ulړN��h���DM�Em)�7���Ȉ�+_�JE��eD��uK��|7�a��x�����ޥx~���̌'�;��x�ӓ�����~�{���/�?[�i�ac�Œ	����׋D�q`F����>xX��/��n?������G>�c{��-gΟ���͍{���E�z�]:��t���(I��^!�&���/����������'�eu��b�D�ݲմ�&�ݮ#�x�s����� q̓�w�Y�����>��TcGBD<����W�A9��H"��������~�د��B\N�S�1ixt�cj��C�bUk��y��i�Nm��S�T̵���O�=����3s�:QJ�T���P�"��	�� O����C����/=����O�?~��E�!�����c/�/�1�'KH{!	��Π?;NRIbo�m<U-^�{;;;w�x�䯿��kg��9;;�����n��^�g��%U��A�M#�LQ٦vlw��5p
�R�G��Wd�9��������_)!u"��7���������c���}���$0#����T,�0��C#r ޣ���=�!£E��Im�vwjUHL���y�N�|���4��� q+���P ĴS�^��v�_nV7�����RB<c�5 !�$��^9����Z��� ��� #DSG�����Z���UC�$)������; ��`�z�2]��O��4ղ�H���&~Lf��e[ج{�҅����#kG��p�wn��:I�w=���A����r[p�Ϫ���T�_�/��A+ˢ��$M�])#��^�s��"YY�#���?����5W_��`�%�l����>�$����z�öe�#g��x>�4hqk0��fa̒d�u��^�
$�(��0�H*%�dXqTX�sk�Z�.;D�� y�)Ӵ�Wx6��Qɿ�[�w�@O����x�4�s��I�q���} W6:�|?�]��Ĺ��������w�����d��?��?<��˯�ԙs�~Y��7�\Y�$�y��8�qaDDxǤ�;M��7���'��؈`�Mq���n�� ��v�T��EOR
A��tC7�ND�����r	:���Ώ�dQ�?�kaaAE_ˎvP���g�?:��+Ǿ��/|�~���3W��������3o���_���O>t�F9HKxN$�!u��eE*�+��t����O���$�`<��zs$�RW�`�7T�#�(D�H����*:F�G�L��C��&��w�ҥ���>2]���O����u+םx�O��2�u���җ�t�����776~ڲ�7�����,xQ_A?��g��I"��E��rl���~�u��܅�m��֜�:9Uǔb��$���I၅�$ jv��%����]+k��\ʣ���ϰ��۷oJ�k��={��������أ����o���7=�K��K�i�Y�������g/����������;5=u�$R�lyT/�i�"�lX�J����MÐ�H��ky�7o����ԉ�a4�q��@u1[(�:W��?|��E3+���j��.�ZY��C17T���S�N����/�j�[�yOe��g_�������Ͻ�=��:5�����/��w�w�+�����"�t����9@D R�GP@�T�$�q�nv�mnmwv���c���p�DdaR�=��;X/�d�+ys���Kq(A���G��Q�3���FyM!
�m��#HWmmm-��jG��?!�������)��N�-ϭ.//oJi�~�j��������P/I���;���?��;\��.9�ݶ�k80�=bT^�e�5QpiPo��?COg�6h�Q�W���ʦ�,��0�پ@�K& ��ѡ�v�HD�+umNP��NH{���y!pه����Tax,a���eIמ8q�$��\�]�m�:�0w����c����;���65?uɶ�w��JCv�ڑ#��j��(v��Kkkkp��������ʋ/�|�����p�ܑ�����Zu��h.,.,,�<X�^=�q��#z���Ϗ�UbM�T��[I;F�Յ�\o/�Ƭ%��5KAtV��T�!g"����$�n��:�!���+r����RLϙS�~�̩�krY�D�f�EaP���ݔ�y�q�E�uz��/)c���yIPKN�Y��UYX4�EcQݏHP��eA�}	�Þ�"��p���RF�Q�5�i�'��G-�$�����Q�znw��r�2�����W�\Y��յ$����|!(��!r���ǂ��؈��@���ЄA��nu�L$0��z��5�H��%�����^~�w��J�HY��I�f�Ψd�(
2!���7�����6�`GZu=�>��d��[`P$��0N=����~>�0�h��:f����Q�Y���E�J�f��Hd���F��1��LD0<���E�'B�e�se��qr4d*�O>�T2u"��ν+�2�r�ɀn��=�p��x#����d�=��l(;$�>�͢��� Jק�Qp"݋��]?($���t�)�_>������z�����y,}ǽmD�j�qJ<܁{%�G�s��
���R�x#�8"Ǌ�(z��G���)��G����8x��T�̉���] u-j�L�T�h@��I��Ӹg�D�zjw�V�!��A���嬣� �|���m<&�{�8x����{r��$�WD���f��D�����H%�A�Dd�*Zt����vۻ���D���0C�����S�ȵ�=1�r���Mtn�,R��N8cйec��䓈J~��Z��Z�S�T�E��L��P�y���E�T5�ݞH(�t
�H�T����C�J�Z���㈺HDq������|Ϭ��|<O�3S��;Q��E�> d�^���q�;��^0��A����'c�g�U@cd��P�x6��,����`<:��(ǪY�S6���<�(J:J"Τ@vQ<׌�ȹD�P9c���� 9���϶ʚ_`���l� �O�P����}�G�+^1��Aцy�k4�Զ&O��ʮ�ވ�p1�
���̘_"r��

���ծc:�U�2�1��(P ] �i����2���
����jZ���/=��uT���!}�S�0���̺9RȨ4�BS�&2�\R�Gem�\�)�e|��x��[ƛeb1�ϥ�lڹW�&[O��}�<���Ȥs��m��P��3��Ar��f�QIcF�0j�U͚ͦ+����@��c,gϛr�����ƚ`"ʀ�@z[��0�����FGdx51�(Hh�0�$��q��JD'.��ϟ��p��E���.Ν;n�����r����?i�%`+��v��<���<���ea�ުڹw{{[,--8~�����t�H��.]�T�p����ӧՆ}��Z/��@&0�;�8�OL��ñ/����Ry߁�����<�F9%"Y	��:'=�u�f��0�5�-��&���3|7�%&��m�c�#�=��"�H�A0���7�V9%�n$�nh��e���鴟:@ic��^��n�~��툓[�xL1��[�;�cԢ�RW��ul�湼�ݒ��ڳ����Jğ�~W���G\��I�����ܲi�U�ԉ;G���>��x�|]5�g(����.�+CDd�8�#��_�>4	��]�p�F"0F-/�DTwݦ�ِ}�K)�x�M22��Q��凌o�H&0j!�W2��=��XV��1GBA��'���1�8"�.�Ү���{���>��u��{�{�+ :>�63��:Fh�|�e%ռ��e�/�x�ԉAR�[w`�v]��#���V�"��h�*�����`a[�ηg�� �Ⱦ$�w�x�_�|�� x�?�-��i�������ݴ��m��N���%���v�(���x��$ŗq-�� �ݶ�eY��ʑ�DT����vB�b�3�����F�?�O���'%��>�P_؋$5�����ӺM�'�Ã��h�,F"E$�)�����Uy'!B�V��N����Z��DLRX���~���g38�r�Q�u��+F{Ǽ�ƓkM���QkL�#h���������͐mh�P_��8:�(4�]��k߃=(��P{����@�"I���Y����M-y�]y�O�D=����ހ��v�6�(e2J��������(±�h�u
)�נq�*�}m���笤9�D�����$��P�^c�b��;��o�0�FWɈ0�Q��X!�_e�`=P��n:�CD�m��rR�bJ�K�笶�$�
�/UQp$���A��e�ѼZ��ȍ�RWɨ@��G6N���?��YHD
dQA�ʋ��m~4,�J�����t4\���PҚ����%#w�8��S$��G`t�����А�-{pܤ��̶mF�B_�_ޖu�K�F���\���]���2&�4�|�/0�H��ND�F#��aF��7�!FH�G�]�8��GXK�X�xF��DdI2<GEQ#A�'Mm���M��(2�+@��f�w���f#[�x�P����z�z�;z�jv/���R�{�!���t�:o2C!vL*���c��7�¾`��{@G"Z5�7.*X��̳)H(���m7�l�0�hӶ[�	H<U�#�ߎ�
�o"؈V#D4��+�d)+j	ey���i�Ш�-	�?���^`;v~%�\cԣx��/�7���;$�P�j��o"*�
d��L�i嗈v�?�s�0%�g���=J[�v�����E���Og�Ì�Ѿa��M" C�?�(���ژR�/�h:#��tC���hD�� ��7p������mՉ��?'�^��n��6<òF*y]>xC�&
�3��JR8�
�M�^2=ۤ�e���
�Զꮿ��IZ KT�V
�mE��$��Z��ڲ��ך�e=��.�xF��*0��Q��ED:��)Q��ͦ���$&���Nk���pq8m��{��2��΁`'˝_��8�Q*(H�@�p����w���z]}!�3H	�("JDB�rYLMM���ާ5.�9b�l�P.�`�=�� �ulv�(P�A�T!�ύ����Y�X�"��`�Ri�^e=�^3n��g8RB�9���N�s�&ף��E)4���R-��b�i�K)����m)�8.#:F(����|��5����2��Y���ܓ�s\���@�aA�!���"���?k��%��#���c7 �҉�*�K<,)�aI����ÞJ-��m{iъ� �𜨫��2�%�1%����}��S#�>�R"ک�US����	�G����u"�^V{�p�p>�^h>~��{�;�l�n��s���w�5\ñ�)�>��C�j���H*�88�Z�q�� ���MjI*Bt�;�!�KP!�D���Fӱ��c旈d�"]����H���]����n�ˮ��ɨ��������B�D�8���lQ�B���;G��%��%��I�#=l�V�rSc�ԉ�4�F���@�1��o]���hܡD2�r8���+�$#����ID� �b�\�C�z�D�k(�y��&�~㏒���N��e���3h׋і�lP�hw�Ĺo�؁t�<4z��� ��@��_��fD��I����T��i�R�"W�<�]i��L�Z�piEDPH>fS�c�mT��h�\��ZO���Z3QHDr�a���r<��5stQԒj�8�2�{^N��6z	8N���
S�0�P������5�N�}���[5~[d�#����e�H����t��fYᶢ��1sl�6M3�i�M��d5�KfX���x�N��9�kt
��'_4IHY[a��(M%�Q�W
Qz�k�	��Åg�)4("J�_�^G�g���EO�_l[����_��%	��F&L����V�Wj�qx��{�H:{���D�*�h�}�50 ��M��D��g���<�p[t:;}�vT��"C`۞Y��j�+ݟ�wO�W�V9��(r6��ܝ�%n�&-��$�Q{w�@�t�i�<ј���L�t��R�c��L�#��;��S[��(A=��;Ma~�|�#~֑ee�k�(+���j�_�}}��昈��d�8�ȥ!�:uZ$QLm���i�A@I�m��UJ�p���Z_D��H�R��꘺��:��{Sy�{z��DF�^��d����8m`;g��-F�2ȿ-W�-PՈ������ߕJE�[�Ch��QD;y�!�X5CB�ۈ�@��I��$���A�|�ӬN�����ߡ��2�%��k���ELD"tE,�2�#
4��ۛꁿK�z����R�FwwI�$�ׁKs�-�zϘݣ�t aQ�X�:d��%�$4���%a#�*�BD{\��2@�3c�R1<�@�v�^ �����4�H�R3:#�X�{"�Q*C�.n�ߎ㪁K�D��Z2��V��$@W�\hj_��m���%%m��;tGH?t���n�m�鎙���-IJ�hٚ{97�;�JD�a������%q�6��D���q�6z���C��� �*HFW}���Ɉ�E��.t:W�7�O�
I�^FR'8�&E��K�a}�	r5U��2��D'T��V���,MK^�m���|�.�~B�v�*��t���D��p�*7����.����m6�M���4�h�pc-:�>�u�$�k6n3h@���,O3=6�4A��&}Dj���\H&�Y�Nz9�p�����EYq�����tt)��K�]��}�Z���&����wQ
='z��>^D|��.QZ�璤�G��t�����N�4\�!���\����X ���177�|�N��{��������/_�%�ѹ��+��ҒX\\T�/'�bkkK��Ύ�x�o�
�{���������}ggg���������"�݃6+D9����1�"��s�XYY	���AN�^�$�Cٝ5/�kssS�	��v��!I���X1$��F4��T��w|��t�t��Ȏ���M7�7����n��t���@<v�x��'�/��fߠs����UW]%n��6q�׊���Z�A!P@ kkk�̙3��^Ǐ�.]R���k�w@Y�� �k��F����P���N�\�Re�����buuU���+�.�Ν��,�'cP[8���C��؏��"��@7�>ǂ��m�P'#�I�����}�1.,,��}���զ�XU,Qq������KD<Z3IU�F�L��7,�i赑�������������=�y����;;ڗ�o@F��A������c�=�/7N������[no�������Dv��,��� M�F"�]�rE�������o�ȂT>H$���5??�^o|�����o�QݟT2��%�Ar�J�;}��z�lt=��	��c�j���׏������>J��Z���Ӎ ��| 1��o|���k���`.r	��Yu=�L�=v{���4�V���@Q��M����l��,�9�]�/�\��
�����9��0h!��Ƽ|F�7��"��܀�w��۷o�"����m�@@TD��{�) 9Э�@�"��� �r��D*��kC���!E>�T@�?^D$� L�-�{��C�������n��V%�}�k_�?�|+��#����=����w�lW�Lbn�a���P��$�]�_�����E�?K}�{�L����N�X�ki�OD%R�x$D�"!�6S"�;]R��Dĥ.!���;?'4E(T���sXv�2�Y�k^$�3}&b ���-oQ���_����4C�2bӴa[rЛb��~��r@\���WR��
2�B��k�@~�}�{�=Q;(�XeH)�� �	߾�x���bV�YID+�,oz���#׊�gψ�.
������f'5v/�p��d�OP�;$]a�r(�, ~H`d�'�.yG�'.e7ph3���aKzڵ�XH�]�\*�S����T_z������U��"(q�����e7�A��s8I͠0p��	��$؄��ZZG�?�oll��_]�b I`PC��db��Y
�� 4H<�AM#	uF���:)u]��$آpn焘*�	U:HU��<��II0~;�~y=ص��.��'�xB<��ӡj�<� .y��xW�mD�Œ?�]T��3@��w�0q��,����u�A�Y 
���{E������[ۈr��Q���n[Ѱ���t|�[
B%Q�N�`�/n
��RZ0�"��54I�@�i�>A�h��<  �qo�D��~�/	IbRe�l9ȶ�ju��)���/+�e��r�w��C53b�C�����(��)�|�ΡC�C�~��5�u����3g�)ma���5O��}P�����<�&iB���$A�&I�XR��x6$V-�\�x���~���7��j���ia�-a���9��qk��0L���D�"d'2\/Y�}���Gi؉t�l�?�9�P`�� ��	�Ս�	t��A32l%WIiFAu��T�����g�_|�EE���A[��r�+���mB�=�����GEF'N�P�!@Z�dt��%i�U ���2BC4�AYQOj��C������r��;Ҹ/ID����w��zd���l[(�YTS"$�5PG|&O\иbM��x�X�ԬF@�\C{�!4�G{��r��k��n�W�#�H6vb�H$�p���������ns�i�������ة��q�\��c����^ �������7�����D�����஼�3�<#��/�R�Y0<��/B�� ≀��yEVd���P�h�:7Ρ�p�ɓ'ţ�>�$0�������?��a���%����q+�A*(�Jv)ܓ��΁��v��?��8{��z��?#���J~�ύ��a!�hRyb}==��0�h���%�����@� $cj�w-	��#��gL
�À�`����=�fd�f@� y��ێx�0��`�?���.0��;�>���C�tb����2BH(���x�7l��rq]܈��	�`jVH�A��DP֋/��)�!�>����p=��$�R�'U9�1Q��w������$
�} "jk""2~S�;��xqy�^���_x�{�j��gJɷD�pV�������XK�f�!��^.:B����HM�JH}���Ő{�.��vΖa�6��A�A�����:�s�K
*euv
z5H��	;�<�������
b��'���@����H�W��$�s0�`k�aS�z.�j��j�ᙕ�@"c��K%35=+IFn�9�l�������ܙ�b��e_⓪於�����q��c�Vp")˩�g��){J���EUo?�׷�]U�~��K/���7nx���Kմ��VmMhR
�@N�ѳ�G�rﻎ�u��Tؿc��.��;q*��?����!��񹹎Ѡ
�䵡MW���;ID����FҎ�Z��N���P7�|����ep�T4C�4`ky��g�;�*���$@N�OAm���{��p �����Ž�ޫ�\���;���V$)��u$i���k\/�ڝ�5e�B��K �����(+ �%�s ��Zv������FDҘ�u�aU�oK�[}�٪n�	uB�;�����>�mv>"�����g�zYu����| ��i;ۨ�2����r�3u���mJ'�8��UG*gTnnk 	�Vo��P9���,G�"x��9zT�Y@"�jH
�4����W_U�$�c��� 
Nʧ�~:�s���/G^6ٸ�.	��~�4�N*H��|�9��߃� Ł� 2(�I$�6.Aə��Գ�ŅP�$Ւ"�#�vC�\	r��kյ����:����):�L|^���%>����d�i��U���2b����_"�?at�"����đ��<Σ�����%���6�S����Ȉ�,�$�`��5����H"!I�V���6$^ZA����O���)��Jj��ӕ)E��.
ւ����P#��@�h��A��7�	d0�ŰdӢ�%a~���Lτ&~C��s #z��r��R�"""�����UDJ���Uu�W� }	V�'L� #/���<��Ͳ���i��A'#" �~Dy��~؝T3��Ħwru�G�E+��s�=����x!Hp��.�AB�0*I�?�@2"���|�[��������f�N�R�
��ɜ<_���Az w9�Q}T�-+�=��������7�ئ����8فx�������L�y��":�ybƘK������ �"���TE�������i�[[$�'���{19�cC��~l�VF��ʐ[�Lv���ɬ_r�'�����Üi�!M�ݣN�SN�������y9����593ӂP��8M�:�&�M�DR��","z�#O����\ၴ�kA�"����(�GPi��� �긻�x����
j(h�r'���Ҍ("���������IKo@*t-%V�ᄁg�k!��"�ٮ�$H�}��ԙEE3��6=_���I��C��ўʴ-��Ͷ\*��%�� ��=V$�2RFWfK�ߤ��泵�����A�<S�R r���J
F$(*�� -*C=�K.pM�;���b�PbҚ��Q��HUM&��*w�>I\J�5}��$!E� � ���	���eU�W��"�)��Px�t�Rq�� ���T[��~�F��Ob��,�9e��� ¨���ĉ�Qe�Z�Y�D$#Z̾��O�ѣGū�^���'�'C5%4R�!,ˀځc^��R�u߻[y�`/��
$(\e��d�g1�EӺ-��&�\ɣйt�	�b��g�$�Բ�!`�Mp>ȗ�u�/��2�D��@`h�[�x���젮*d@��*�t�P���\�ɟ{'g�0��>���M^�*�c�MϢN�:�uېސQz0��X��A��0g�na\m(^�0���c�ó��TK7�q@C��W^S*E��M��$	�nw��;Ԁ�`S����i�OA>��@Y�qa���'�U+�4~����w�S���A��&L�����D�_�J[�p�������a&{���3F�څ���0��d�F�$��AB�	����&�%y)��r�k�;"n����Z�+\��$�9�W�i��Q/��'P�$Y���I$�F�}�H�fkH  �ŬTԬ���1x@�F&�6O&���1 �
u�7*����8����~��/֛!��G9�@6���|�H�sj ��	�e�1]I���PO�l��<��`M�=a��Gy���;n�'�T���BZ���CQ6'�{"���W_��e͑�M�����;q��V�kh3�!R-�#�NH�gӉ�A�I��2Zg\��r�A]�ԭ�++"�x$��1�c0��A���Cyq��&�j9��\� S뾂[eb�o�C�Ad܇<Q*�ځ�JX�y�f?ϑ�~I�V(�A�l.��`�Q��lA�0Z~����\�&�:�(h��lj rF�"��쑔*�b�(&��a�:y�8q�a�{���=�r#	�a;���� ��0
��ѥ�Kᾼ\���I��lA����gU����y�����7#B*yw�۞���P��5O�� �8`�B"�e��<�0���GL��<A����42�#b�{Z+����� I6 y�Tt��2��y��C܋��៤%���{Q�#��#�#��Q�~��O!�.D���޻b�
&�	��^��	>����	l�AQ� :�'�B�`<H�
�Pw""�F�Bc���T���l�ʝN��15�,�����QH5ۤr��c�
HH�t�@�"�8^��w�`G�S�b�{r�q�]�$D�&�2,��uC<�!5PW�B{��+�C�hw@m�Ԑe���N@`���'���6�v���=�NRz�hvzՌˀn��fP��q�=YTӢ�E��ADʣ�TR_0cC-�$�g^�HC5H��yds�e�&�	ĐD��J)<I�<8���|ΰ���HuRe���T� �� :�
�E���� ��! ��o�|�)B*'��㹫�jHi�$�J�����äl�}O4 mD[*��Y�c����J�US%"����H=1N4I<�8�@d���Q�ٓH�T3O	K��@D����C��K>��[<��D0`)���P y^ɴ��nJnF�6��o�#-��C�	�w��x(�I@�CYq�)����5a�[�^�&8i(LQKKK�Q�6Z�B��q}��@=�2��#[V�p�#��b�*���"�@�U!l��'�A��I�K2J#P������羧w̂�Ss�-�%��`�a `�ap+׳���FD�";
�A�$�jE�B�sefZTf}�TC�:(�N)���T6�
s]�=�ނ2�4q�HFr�h��`�H9� ��k� -��j���� ��Fs��}��~Y~�ͭMq����SU!
��[�x�莺�=q��!��=A��K�u�i���h���k*�4�)q�=�AF�M��C�*�KI{0^�]����D��H�؈�ma��KBQ��vU\������w*��!���������T�����)�J!��ڝo~��i9Hq.�2�b�bl@���*��d��Z�N�|��i��O��//��c�?A�%�)������xí��k�� '��q�>?�G��V6�j����UB�Z]�ť��"\�(�����0x��	î%7��������cW)�內R�+C�"���l�N���P��$h�8 ������I�����<�DF��b���!��k1I��v���=�GFD�N�<x/�ql�q�İo�6�Ȟ�:��#��JPܐ�h
I��`j��ݒ�hMT
$�4�����A�6�(KANhx��oP�b�@>��킁2�@t K��ǑV�ȥ�=`��z)�< ���������O�|���2�K�C#�"Z�J���6WVо0@�syM��qP���I��y��8Ժ9��%�\����A����@���#
���%ʁ?D��G\
$Odv������N�;��(X���I�@E�B�	�0K�*qX`W�-�i�����G��K �a�cwW�Heܐ�@��Pq@{I-�\�@����0 �@���ArPY(RD�?+$�mTʍ`Y� V��i��dt(Ġ�]ci��`	�"D}?��SJ��hf��6 �� �n�Q� ��uѡ�x�M7���ZF9�":<ؒ	R�w���N^7J���$�.�(!����t���f�?�K��pwHKAl�|J�J����C��;���s�ҐL`�1��ː�Z�nP��Ԭaك�?���b���!��E�M��&%+O�?�=,нA^�>���7���Ɇ�=�� 9�b�@DP�@Z���ܮ�(�d�z]}�5-	30x#Z�F��!'X6c�i@��6��M���o}Kݟ�%�Z>u.�N*�x\=%���l����eU8���d�U�7T�T�hu\���H��Ä�T��[ξn{�7�x�-C?�4�~�)%=�Z�(VGE�r����T#T�j
Է�}N|ʇ���qSy�L!a���nyɿa@��/	��*�K�B����G !�8-�N H.��r@J�5�i�4 ���:�"O�E���u�J�ĵ{�1%ݡ�  ��/o?�$xR�5bPd�t$�Q�fxѐ%��i�3~���� �1m?�-$R�0  ِ{]�z6�1��h��.�Ka�1��� ;q�Z���w�;\�� R?*,�>���c�����IP��! Ik  ؉ ����ϸ�J%[�:/_��h[_C҂D�-�pHv�Rʲ��J~262c�W���=�6�u@�J���a�ލ �%�x�'$=,yѢ��I��J���s��0��G-�:�^�Qѐ�- ��a���qeǡ��u*���
�P���]�m[� %!����]-�<�{Y٠�x���S�iZc���^��M����� ��zZ�O�yԅ�@�x�M����(p���> ��}@����~ w4�P���VYO��ǩ=��ӊ̰�ȧ�@L8��"q>�ܓ��Ƌ��RVG� ��}�-<.��
#T�H�!�nM�,�����<�/�!���ևݞ�ЌI��^�: R_h�TR�"��>�����M�m���U"24�r"%���1d�Ȋ��H��Y�z�Ql%{#��A��o�l�	ISP!�0Q�"ΧEQ�싁�����'�F��#r�k�X[�9���A���ݑzd��TR�  �:�8��.t(7l�2��{�(�<�ȋ�Ô�[�k�d�4����h�*�`�D�K��R�VW���r��DC[� �������h�S��|�y"W���7J��c���w��Ì��`���?鷊�3<����F(�P� ���NC�˶ݶ��Hh�i�'I�<��;��	���=�$�*%ث�xL��]�HM�_��K����4 �c� '�JُTv"�;U�#�iݖ�M��V����8�.�����I�����=���e#�*�׾+*I=�ۦ���"T���lz@h�m�Т�-�c�xݨ��D��Dk/3���}3�by^��-���k���\���������A�gr��Z݊�8���,0���x��*uE���#�n�p�$�~���ep�ؚ�x��Jצ���|��$���.����/n�_��D�$���+5�2w�m��cQ�v���KK�F��#����VOK�홌��X�٘ȑ��g"��v�VG~�#�Nt�h�]q9���M��v�ɈO�JeUj�h'C=�8ՙ����v�5H�4�s�sU<J򙪔۲<�IWI�é�"#w֚4��5mO��iڢo��� 4�p�Yx��[y�W-�Pq5*��\j�}�V��$�pYaMk�ԅ���1���:�g>h��K�Q��K;��)�t)��ǥC]j�DH/�Ֆ�C[�AN2�����㆒(�Ѳ'EIDTn�=@�f�j�N��+y�!%��Ӏ�oG��~(,��$	Z	D��C_�#�庽Cu|��D�7�]F��w�v��q���d��cMM�2��v�H�5�E�� �Fq�.#�)���d%�Qui�`6"���M?����qRGZ��(Ծ��P?�^���KD��N�<.|�p����iF�&�.k�@�����I��s�������^eo��� ���`����KK���"^N�G�p ��g��d�f32v�'�.�3����N��%�=��~$��fN�FJ-���=���n���q�~�1�1��DYC�H�K`\J�8$>��N�q�:�ģ�y>�V�T$�Ƨ�k�H����Z���̈��0@+��T��1Įl����g��4��Θ��`~�VL��9�6�5Z�!8��A�����Lx�_���Kq�:G�ޢlK\�ӓ����"�г��䫮��Ӱ<�m���JCa��JA�k�3W��:�P/d�#N�Z�|ۅ�lb�3��ɭDT�׽aو }v�g�^D�4�ʖ`�!����M���k���s�};�&��v���~�Ѝ��l��(GP�?���r��X"JZ5�d l-�EF��=����o�v�a�k�����qd�IU��x�s����î�)��ثf���$�$���ףs������~��z��t���k��ōj�^�5j	�WD�dW�e5�̪f�;���	f�ҍ��Bu2#���W2�zN�ב����1�~�n�~��K���K���"�4l�QIՆ�hM�ʴ�JD��k^�H1;�s��;j�6��=���^��l�h�~=@}�;�`�!�6�u9��1bl_q��1�U�Z���#�+rc����t���8��C?��g;��pW�V����:��Q�c�uCķC��N�Y
1<�ɬj��>�$���sQ���a�W�}�(�QG׮>��c�ݯ�ۦ�Wt{Ɲ�b�_b��q�N'��0)��D��Q�f��k�6�V�C��ߝ\�Q&�x�x،����ۼWt�9�Dv.DS��:���P`��u����.DЯ�:m�Mܹ�;��@TQ�ӿ�O<J�$<�p�'�=J���;�Z�&H��n_�&*>�������Q����AT��A�a�L�Dg��j�ѹAx�.�� �S�{��z��-��t0D��D/�P�	�$ٖ�v��L]&�����y��g�~d��A��:y<�0N6 �g��*%�`<R��'F����̨1�V�)�v��^������#B����2��jܬ� !�:�FG%�G-���δYU���	�.�-G�mg嶍[r]�~��Q?���D&K�3&٤J��ax�rY}R��'~�2
F�����6�eS#��%�GU7���;>#�25�a�%A��Nm���w"���uP&IL �|D�Ǖ)�|`Eͧ�^�R.�ޢh���vu,�M(�`�gLIG��R�F}z~��=x��.�5�R)l5 o�(x����}�E�a�D�ft�:��q���:u�>Գ����$<3��AG�M�ID=w~#���ۊ��b��w�¦�G}VO|�߳�{��l��3�W�V5[YY��J%�q����AWI{	4�&*�;Nf� {/�n��P"
$0Rj�M��wb4�Pg>���c�A���Lz�ðޮ�����q��C[�E}�z�\_'[͑2zKý��9� a�G����&����[�k�Q������;^�З�pt��G舕O"�p�o��d�%�ٰ��Q��W�;��0/Ң艉f�����
H�Д�Fdm�+>+ހ�tup��.�6�QbX��4[�����Ԃ|����!�\"�S��o<��j>)���`d�n���mD*	�y�@��L{��h��=%��&�Ҟ���+��-w���.&���ύ
ZM��t]�2���\֐�Z�.;�N���8l�L�����h;i~\�^'�-����wj�n�@�pԧ�w�ʯ%�ؚw���s���Ku(�o�v;�|�3�wI�Q�#�HOs�A��[j��u�͌��s?�$"��ȝ1�֭���">a��N��ٚ3zq����X������,SXt,�}�m_nx�mW���E��o��a{�}�)�4�<`�7�=�����?��T��Z�z���wC��{��E]�w����7�Q|��#cDϨS�UD�!�W�������[j3���T3�T!
Q��IEQ3*�1QШ�Dw��1�D�Mz�1��^��&N�N�/G�k��;��f~��5��1�ޟ ��I�j�^��� �Mh�N~���̂�D�{�8k� ���v�R@r<�
��\��:�-�xss��%�i@_	�D�����^�a��D��kQEV�|};��U�:�c��?M�y�����Q�I"!`�����7XNZ��H���6dv�Y���镀&�m0��l��׭��8�E���D��B@:z�eT`�Яp�_"���6\ARn1zD7ɦ[Φn�Sx���__%5��F_"*�+��^Z�!�1l^��Bj�^>%"�5�\�۬��� ݰ#�s�0'�U͐��t��v�S�MB㴰��XA�U3��Yv%���2�� �Âk��Fc�䡌Q�=^$U�S��a�["��z7�Ƚ���h4�8��"�IA'��5rLDHZ-
m+�E��R���旈��fI���}=lI�ZY���*[nך���܍��U��BVIH�l�h,0(��ì��I�'ku*0<D4v��8::$Q��ԩ`���F~%��X]`�(H(�H��z�l�N�^aZ�X�x�Ky�EO�P"��Q��]�w')�k`'EB2�.��^��5v�yR��X�/䌄����A��E����-FAD�H9�
d#�^��`�l��6�J�$T`�����t�[=�~�Fwݳ`�Y°���I(m��j�Y]+�+P`0c��?�/HhB��)�P>�B�(�}L	y���%�b�rE�a�8y���W���tʻ��ԉ��5��.���7���cYO�����<7�k��Y��>|{�$��e��ZxQ����ʆi�Pm�WX߳]G�>���uO�s�ݫ��:�ߍ�A�	���fQeu�ξ���瞯�	4��daz��O"dEKRD�zޛ}*�-v�ض9�`�@����p��A�@픲U�Qi��ѝ�LK2Qj��*U窦l��`�h zuC?3k7��Wt}�Jxi�f��~��~1R54���ۗk&�%0FQNrQ|'�JD�͒��DY@�lU��*��n�T9`�jG?��Ȩ�5c���{�Gܵ{�P�����w�0�p�L��!*����/��CF�Dd�6��=���H�~+�2Qw������+�5u72Hj�哈�\;I��l,�FҤ�/�j=�	`���C�[+++��C'"��_�ߚ��x�N���!�=Rɵ�>��B���={�&����IS��н�7�;[�#C[��M��|�wA?�U3��.՗�o|���C'"�,K����6O��s�q��*K%MZUy���T����eYm���$f(NDx�<�ݡ���2D�D�W���Q͜]��5U�(U9��{�n��DD�~�S*��8A�ϰ%�n}	����7J�o��,���1-qܴ�k���>1�
p�S��ٽ�ݻ�����������Fӛ��T�e1�	;���l �/�����s+��I��{A6Ԋ<6�N���r�,j��h6���$ѩ��b$.LU��[�-��d��ߔ���X�u\��u���,��PL[�����"�gȧ��s6<�s@\^�98�{)Y�s�Q=/ Dz�h=$�u�D�ɶ��n�$���x���ayVEN���j7,..N����z�6�`iҧ�ڏӶD�RQ����lX�}R��e���]vkNݒ����3+劰�s�5xj[<jC3F&L����g`P*b��
�ml���?W��o��u��ɅC^�Ãp�u��t��lֺiZu��YoL���j��a�W�B)D���A'%[v=��a���e��l���*��Z�sk33�bscS��k�+j�8��tY[�.�1�v*SS�����n�i1Dp#x���O�����>��/�+���\FCv0��`#O%D����е̭�+��W�dmc�6���;�0�:6�
�I������u�����SSSg��<����}W]unF���lZ�Ri�M�f�p�q�7۰mG�Ӵ�U�u>��;ήk8�ݱ�V�>Hy]�u����=��V�k6m��)�]���n�n��v�ٜ?�һO�:�1�foB]eg�A�H�R�0�>�n}}�����_-�-~ey~����¶lQ��,�aY3�l�]#U�a �nQ�e�;�o�ώ�����,���o�dKs�1˵��ϓrr������^�k�����^��t����O\�p��mp�)ڕ��0(��xf x�)M �ڧ���*��_.8���3;;�lmmY��̌���#g���0��@���Βe5����O|�M�F���7��o^�o���?��gO?~�S�O�e{{��w`����ds"�臈t��J���������k�9�՚�>.R���}@���O<���[[�U����ܜXXX�I-3��ۊ�M=�{9 �����7������������}lU����~���zn����`g�v��8���t8�A��7(_ZWZ��榺���ܱ���?��w|�����8�.U��^Z�غx��yO�z�8�D ��t����3T?\�jii�^<p`�c�XnH8������b
:��9ž}����8t#"����ٲO��)�2K~�(8�%���k@ �����ӳP�U���$jCB?E��v�1���Ғ8p�U�Ɓ���#��Çݹ��r��qC5㈌z�j�5����;
>�lz�TJm!`Z�˰�%Y_�ڀT�n36I:�����v���2+R�Y��]�<QZ�-0x�T�mɌ@��Å"�O�t}��573F���#"��].ϕ�A��6�F�wq�ׇJFD%�S�S������R./I�5�.@���[խ�y��g��e���kI��$��z����:,��,�b�x��ҳ�:��i����4K�){zzl�u�h�4K���S�2=զ>�ԋ��u2R�hИj-`�)g�ZSxR���iz��N����U��$7��z��{p�?"#�<nMK�N��!������~���:��>�$���k�虑F@�����i�����)�֞��m�ǭ����#�jFĥf���MRW��$>���C�	�D�@��cO� (�gi�-o�Ύ������,�� \>)r���{~]��UN�B5s��a7�!_B��x��t(6"�/ň��k�)� ����w���Nmg$[@3R^[2�eb�?�w�z�yxW0d�n[��{)Q�ffQ��� �p��F�1�m�����s�Z��� �YWQ>����l�U ��
3Q�~?���F�^�Nz�y���H.�Y�rn�PFWy�Jq����8r��A���Mh�e�R5�V6b�1�:�N@�/IE|�q1xd@j;"r�\��Z%N��W!��5������l�m�d��RKŝ: ̐̕�?��nm�[�$"@���X�$��Ё����#*��m|�h�H���$��"�Xۺ(x�'W1D�cpk5%Y�m痈��n���L���좆2:L��h�+�/��Q��'/�S�CJK�a�Y�|� X)��C#Z�)�Fn��C���3
���t	�CFtp/�Ƨ�#�Z�aI��M�(���,ґd���f�#�W�x���l���$�q���v�#��� ���F�!�B�bC�ÞiU�ܵ)�_�֪^b$�G�u���f#�<ǒ�|�79"�5Nk��0f�IEЖ�9#ǀ���X� :E��>˳�F6;"2wL$1]�30۪Ŗ��ȗeZ����s������>�qZ�w\��jes�U�b���hs�$�6Z��ݯ#��i��&zv�C|��^j�/\��������>�b��f��C"�}�H�CcˎZ2^5�2�w��jf�d�C7����z�q#!��狂�7�����}y�$�YgDdf�;�u�tO��1F6���?ؕgAX؃V�4�;f=ZK�Y+aa��`K��-��5��첒A� -B���\�c�a�\}���]U�_dF���̬��<*��Ϯ��eu�����	�.��N"¼�A��!IF���=AV�Dn��p�,+�z��M��Kצ6\ȵ>��� �xk��`�R��\iL�L՝�R�mr��FD=*�E1|�о�2(ʄXW���j~±�_��?w��gjy��el Y�GWY ���Ո��%����E
��1Bf�kaF�8`�ғ���V���U����j&3<:��zF��Cs���N5�\3T ��������	�����:/�d���jY/jᲰ��$�ū�_�O羦0����ѦT�!H�(պ����,���ǡ��'���1���P�0��0�0��EeQ��utum��+�Vi��M��W��^/D�!r�W���9.����y�.눈��a��Pg�=t�#�mA=���rn<u��(W	)��2y��E�t��ȍ��M�����%���5'���|R���1��(�D���3=�C0L�#��e��z�jι�^������ཌྷ�5�DT��D�+_ƿ/���b�%����^3Y���O	�D�.��e(����6z�M.Ѻ`,�K"�l���:MFm�,nN���Z�V�$"��-�L�0b�K4C=�?Fȓ�[����̩�D�U���Z!&qz��ID5ǡ��
]�c�U���Ȼ�[�:�Mc�Y�W�X�{����<t����7iI�TQ4R.˭%D��*{�eEE�X�6�?�N�L"�f��$�VPǄ-$"27�OO9_�{ͺ������7JHb���h!p�nn�s�\M�h�hk�԰ʢ4 xhSyOD"`�ID| ���d�7�(ûPx�Y���\aW��D�Q_�V#zR�N���Գ��vQ��,k��J"�,pO"�@��^"jY���^��s���Y���$"w��s�:[���R�ڶ��.��:"��J�x�9Q
YK.�B�]3=�\6���h��E�A�d�����eN�#���������#d�=⑃�ݍ�G ��[	�"�O<k�\n��5z���"x���Ō�?�7K�rj�(�8�_$�$��~5�������Ɂ���#�7b��jc�5=V��uD4^�E
.81�c���zY2-�[��/4o�V�[�9tU":::"4�C�4ZV��j�e�Q�{��]4L�����ZY9YP%ȣ)d6"�JD��*��7EE,:q�Ά��d����A*�L�һ	v3;j 6"�[�=	��6�"ˎ��%f�в��p{��U9�E�N5�D�Vf&��&-��������f=�g�Vm�E %"§H���h�5���W��hd�y��1I���q�`O6" 9
���4�q� �h��{�Z�����I�:"J�DV���u���Ee�S�p���P��M�Ed�fY�h����l��`i#�`���+�w@����5��"Q���HE��-��0k��5EB������j5℆�9Ojn0w�� pV(�D_OjV�2>�C�#yBg�JA�!���ϭ#���S�`����WQ�c��^pM�x��]�y��YX�XǝT�y^�v���u:�H�J-���*�?��M�����qD
Z1��s�̢�������D�ZGD$��2�U��ԑ��`~N~��?ݭ���u��5���b�<��J""͸D�P'ͣn���RfS���GvT�c5Bn������l��A��׬	�x0gU�΁�ޠ���$T�Q,-Ɯ�*S�tTCT����;�,���?HfF8!d��ְ��I�X3W"��^��ٿ\�D�K�$G.��@��lDve��GD	���@�����M��*�h������%0AVM�������c�hS�"��u�5k��J~���YA�d�#�4H'��}���Y�Y�6���ad�N�����H�� g������U�9�����p��`DT���4��;�����:τ�V�	�Xɣ:#X(� Fd��(�ZX[+@�&��:"0��<o�ib�7oC�]���W�?�zGYR���X�8�^5k��j1�)�W���mt�p�\�����*ilD��[b^5�Eyb-.lU?q���/��4���&2�-�[�2�S˚�XSl@����C���JS!�wzm8?e�x!���E��5�{1a�u+3�!+��A`�IS8�6���i���AeI��u3֪�Yu-��k�ߩk�������uH��y�A ��g�^�3v�PTs+�)�j�ZID:�Ж�誄�2�ũT`����W`�C��޾1شpS�0�6�xW�S�ꁧ�9��o���-:rx�h��Nn�ㅊ�D��� '`,^"j8���I�SH�o�b�|LY����q��@p�=T�:��Ms �_�`��k�*�1E�H�n�2L�Rɥ"c����Cꤺ1��a����\iB*�1!<��8�F*���x�9KW$!�B����Չ;o�u	 �)R�O-�LK666��4IE�8ե��i(�g��)0?����q��O�Q �)&�WGk��F���҇f����R��:��x2)�&�6TL������EQ�&H�����c��EQp$ƌø)�L'h@U#�{B=���Z��u)(p"β*���q��eb�`��D�#��Sd	�#"1�0��nH6Op�T2��ɮ�յ���)�`�p���@��K��O�g�!�I�އ��������D���H�qOن�$"e��D46FB]��#"�1H��ã�#$�9���q�p=����k~��Ծ~���ܝw�����Qb2>�b<9�V�����N��Y��wj�ܸq����Q4��S@�8M��>X�@���X��t��y�=2�Ά�0j�wta����)9:8�����͛7�RR�3u�([Q��lʕ�������a�|ūкc��k|m�C���])EnllL�`z$�
���&����lFؘ�o\G�Ѩ�Ͳ��	><�k�_�vm"��k�	�H�3�څۍ���^���5�ۚ�&�$ӻ���8��6�^��.�N) ���ؘx�ѧ;�����+<21�1�O�:%�t{{{���%�")	
u �y��q����$��/'�3h�yA�v�_ID��4CY�]��1�u�_�|3�X���h�a���ٳgl�k�Dպ%`�{�':��l��&��Qc�67����H~rlO�>�{�A!� w^�> �Oy5Ằ!��@͍� u���	�c`ziW��#��5\oEIt�a�}�+jFQ�a�a�SUޔ�LM�\3�Z����4b��@l":p3�%"���B�X�y�������6�RAR���1�e@�5�'X�}��$)����Cw��o�j&NQdI'�޸���6S��1Ll~]ק�;�#"�m�s�b5�*~H�#Zzp$ ����d�P��G䣤x�k��D���HH^c���5���$� �|�(qYլ�+4o��'�*0�.6�6��QM�Q�ά!.�ғ&�F��d��a(�*ף�u��l���6uO�U�`�E�$" 曑ի�����&��v��(�53CW�5S��93��]�q8vV*������V������SP�.�wlS�'�H68��'�y��i�N����oDWĜ̻���1y�c�$��q�7~��(�k������D��\����4�������kcODm��ʛL����<���D1mGr�D��f�O���q+;��^�H��mw���3؉��vBm�\ʜH�:���DE�#���T��>�Yې�PE�`]����Ԃ(:�xv�ۿiJ�����I�e�΄E���!Q�l!w7�c@�(,=nHO%*JX51o�M";�>�j\�#"y����|���W���f�JYA
5���#��������P���ˊ�Y"`��Q�9�Cj���B"�: �trMB�s��Hѯ�{{X_�JC["7ϯ��W�<��K�Ά
�vN���E����jV�P�M���H"R�oeP�?#�i:tn�H"�ɽ�f�<*�ñ��)'H�6������ųT�e�Q�8�\ua�ɍ4T$�5�7�u�rycu�P#\d�)��H��զj&^p6A3��o�c�n�����U/�=�p�,�Ъ?77W���x���]�w�)�,��]�=�mʋ�h���o'�����ݲ�&�c���ᦍ�Wo�@o�P; ��g]XGD 3O�LKX��ST-�L$�;-1�2='L(
�[	�ex�"X׀�b�kf��յU.G�8�˚�u�X���|�q�h��!j?
�ȉ �j�El�M�zլ=؀���@"�b3�a�lCx�=ID]9�h�z���:����
Q1�=���wy@c�������P<��ILӔ�w��Nm���H��W���I����5\��S�6�:�$�iB���)�f����y��M�^�B��♋;I�&�.��p�3ZLblְ�26k�nZ�V-%�7M}c��^3�ր͚Y
m���F�:pO*�mѪ��t���j�^jp�P����ę�����xf�#�@Z3s��C1��5��_w��d�X�'���,\e�.�IM�-*�e�;iv��h$˫�3�Rec���Z��QVZ���Y��x�D��Bh�ф#����)l�rGGX��d�1����K�\�#<��T5�¼�e��kY����d@!vX�o���#"�s�<8w��C�X�u1�V�_������*	.eF@=��ʛ�XHDC����M��G�BV4P�f���:T���
DҌ���F�a!t�ʥΘ()|����Tg�˻�����?�D7��A�*�Gz���uD4d�b�*�<�4�_;r�6I�nI�e�&e#�x��x�f�Q��1��&��m�&���n1@�\;Gl�%�阗�~Dp�6^�V�N��4��TM�J"�Z/'���)��sm�fR=��T�e���>�kw*9�	5W]O�}R7�lQL��V�D�|���&�j��i��5��:"����h��Z���j�a(����Pn��zD�a�70[k����0��v�uDD��-�M,z"�ٗ̓*����[(�[N{"�$���Z�^k`I������yIEn�EX6�� ~�ı�dT��e��T5��:"��Lﱕ����ٞX�B�v���� ����� &U��������t3+��Mj���ׯD$$�#!Q��X����r�6V��=�,�� YE�V�B��e�N�lDȚ(�%�X���5.p����H����i��n!�N+`35�_�JP�a;��r����������KτuShɤWʸ�s�X ���$x�f�p��3���& ?�ɭ[�u�<�X�*�J�)�*}��CS��r��b`��"�n/����ۆR"��9�_���(�*x�@Ó��&r�� ��sf�q���W�D3D���v$��s�ۂT��N�fw1���z�X�Ak��x4��Ao#j����W��}�e<#$��Y3�u�/X+$�u�ԋ�!H�3QQ��1��d���N"�S�9n}�z""0�@������A(o�8�λ5a�ţ�VX�X��G�k�4b�����q V7��5� ��̠�:V6���т;�Rodb�K���*��	i�G"�Ⱦ]Sq�$�}P���-x�-+�����jVw0�y1w7����j-Ɏ�"����	�]8P~�s�/�nm��[�*~H?a��*������e�Z���٧���1�+�cw%�l_B"Rk�d��2xլ��T]$��KDK�FK�l�U3�Iz�Ј�����p���fpQ�X �(Iv��?܁��W��V����k�y̅uDȽ���
�Ul�6W�G�<,�'�m*��D����~)���B��.ۈ,
�V���(+���˥b=G$Xh��f�6�n��AG�fO�L�p�G{O 	Q���ϲj>�!���$o�'�ڥ����A@�y�Sv�6L�z'k���A=�c���	t;�;��BM�k;��zCwPo�� �Q��$�YRM4��D�Ǟ4�25Jrr�C������Jz*�mcn��P�Ĳ�C"���)ݲf\�$���-E�˸���!�yۛ>~�U'�"H�D�������9�tk�Z�^�$"��Q!��w��'wo�Il`͆Y�X���k�!1�p*�*[+��'pLܴ���-���Oey�:9�izl��&!޶����F#kN+���&ղ��ʒ$qn� 	&"Zz�.;b�RgmDi:e#:v���S����tggǚq���p?Ѹ��2 �t��ԃ�H��D���TxAD<E�N"�)c,��A�M
2f��7C�|:�w���I@C5eO6"k��>":�~c�Q����x��"�eeg���1'��A�Z�U��Z7�zN�'ni`$�ڈ��u��ȓy�$L�W`v���%�vO��M�o��S���}�'@���ӝč���&3�uDĆ���PVa��ŭߚ��&�8H�8�fr�"�u��o�t_m�E��B�et����`Ql"JH��a�$�;hd$֏|���]y��i���\n8�W��Z��r6�Q8KSyz�I�j5AJ��H�0������6Mr��8:�U�y�^��1��h�k�5�J����&x*���О�z�䘏iǩ�j̛.픕�){]�w�']:��%�aB��U�l�#"��R��51������^V m���Op�D\����Ϭ�I�*���7���O��[����~[�ڠ6����-��k8���qP�z
i��>��E���f�6�fJ�+�J�K��k8�導����e1)p�n�b���\�E@�эG������^pR������0�4B�5b������h�z�c:��L?���q@�n��֥j���I��$�2*2�ߛ؇�Yy�*M�R�K��$��0>��:C-XGDɋI�+0���>�l�6�C��I��'�G��nFW=w���'���o��4I�J���h+I No�8ǒ9z��x+NP�X�ݷ�����_><<<�tG	x��Ç^P���tiRـ�o`�)m@}�L���xt����g�Z���.>~q�g��3_O������o��D"��9���Q<��/�����������ٍ��zno�*7���S[W[�����z,����0 _H������LX�j�$#���[\s<3����p�=��Y���|�ןy��߾�{�N1����Z覭hU��	������ߜ;wn9���O?��������Tt��W�"��Ԇ���8u�oϜ������~��>��O���[{�w����
��}8N��*�Lw���+����1HI�͉\;}z�o�^��d�$���ɟ����|�ww���(}������\N�8�'������fr��V6�-��ܺu�(�_��?��w��r�z׻.����~j��{�:u�� "�Ќ��X��τ�*U2
�dF�Q<FBU96��{_����o^B������-��m��GŘ�SkR����k��q��u�9���=|n�98��~ick�w~�'�vY�p]{����~��O|��~酗��������{���'q�w��Ő" �7�!q4��ׯ�>{�5���O���{��N ~�G��O=���^z�ҷ�q�w�q�|]' @]{�n� ��\�q��_��|���ί�؏��Uޝe����>�я~���^$�.]z���~T* !e�6=c�cK�;�V�HJE7oބ�}���}�'x��� �ZAB%l��w����~�r|y+���	)�S�мI5�S����� �����������x��j�p(�o$�������Ÿ�~��yy��cY7<B�l�8?��������� H�Iې�\������{~��՗��
m�b���jFH�Fkl�lw���X��š�|�/~����/G�I�լb ��[���ڕkhoo�ߋɹ{ggg�N�T��ô)�DU&8��W/�y�	ub�^��������"d�Wb��b�l(22ɧ���u�;�h�Y�������m���{����m/�A�_�������^~���:s���<�5�$K}͂4�q���C�	]���uYTs`��{��g?����K�/m�	��b����<z��W.P8a�!L�?��U������*�_S��7��מ}��_~��߼W���tU�H�(|6� ��7n\���~ÿ����Oϡ��|��'��/��w��W�\}� �;��&�+ ��D*�Z�Aa\s���{���.<�,�D�����o�������(^�v���p��e���a'9T*�J��8@D���7w�O}�Uw�����Go��7��M������/��P�cr������lJ��z�El z��ol���?�=��N0{�W>�������A��G���7@*o���)�"`����͛Wϝ;�����?���^�յ@=s�� �������|��_��W��s�KL���S&D���IH�l0��:{���<���^X��`����[��K����?��/}ߕ�W������i�JB駷��B�{�5����o���������F�m��;�>����\���k���z��ʉHيt�K�.'������Ÿ���/�:u�z��-X�N`����Www����| ��e3�Y��$+�=��{ϝ������{��S?�SG�Z0�������k{��$/�F��+��'8&��հi���_�����ŋ�!?I~�7��W.���B�|� �Mx]/���vN%�	��M��g�j�[B%{
Y�(I�rm�TLdh��i��1p>����n��K��/����� KQUnaQ���o��䓿��_�ꗟ��0��C��Y�w�mpb�y�Ļ�����Z��w������K��u���M�֫"$x]%���������~z�����Ͻ�{^���>��Md9�#"�F j�����tr'ڻy����?s�]�Y���t���vt#
×�L�J�̿GU뚁�L�0?��ÉW�t<��C�O�����2�Һ��U7up
�l���kb\�
\,�sDɄ\�i.�תj�(O�4�`�b����#�	��6�Ap��T��'U�(,��S��򾋢Iir�0����,�;����<�(�u��:��i(V=aj����.ѝS�4Μ9�|��"8��be��[U��N�r���� ]潉�JŸ0]�1M��^6z���$�΃sD$���'��Ȕ��#mGq,6M��\�bM��. ҌPˆ�P�?�З��) z����!!h��3�v��"˟1gL�(�	g�v�ɯJ�U�Ȉ���^�k2&�|,��������Fe���Iq�hbl&�����$m��!�D�8i�#"@�^�
�z�J<u#'�xbe�P#�B�XH=�Xn��L|��H*3�:I0��uyL�%q@S�MC�3� �kA �,/Y���ZW��d����(�J�	DgΜ�R�p �	`x�D�K��ɭ�"��z* E4L򲼀��5��|F�k��F��?�Ѻ��Q���&Q��*�Z�<z�W�Xx��UODHL��] �fUW���i8��W�
�Y�*��q���JQ2��W믲^p��2����"w3Q���`�U3I��lh�r�"vHU��1[R��h��
,`���qB�sD~~��2�Y��P��o����Γ�L�Wـq����(�(M��,��=�c� 왨D�C,)S3��)qf\�#" h]�����Ό�ؙ�mrL�S����$=O"r��t���a���[�+�8��$�B�eN��N�zu���
R��48����Z�v�2H"�%�G��42r����.(E���Cj���L��)�^5+�̬�tY��9" ��L�$M朹�������lΞ��`�5f2T�x"2��EZ�PTo�Kt��$��̪j�g_wYb� 9M�-����n�$���so�1!ek��Z�n�Qн����hN*	�C�ti��9�Fy��D��Ջ_Y��Dd�D�}�J+��Ψ2�NW��Y�1R����ƀX��6�BBh<�Դi�C���۬�e�S�����U�%PD���nI�n�fx��F$��E�a�i�.z�{�� f�lѡY�V	a'O"�)��*�����ZKWv岾�'"���{�I9q�� �x��k5t��4�H��Ó�|HM]�g�f9�puJ�Dd�
wEe7�I��r�eP�-�&�+�V�L�cuQ�isg�8�qf��'"@�]���vfr��Ji���6�ZX�	8F�X����F����ϊ�4I4*����W�S;� d��IHd0��Y����D�1��ؙ	n
`T�@;3�C�	a��� �ƴ�����E�No*02�&�)��ŠG�G�c�Z�􅩱����f��n��Z��E��r�N2t��C���9��q�Ǵ ,Z[jld��C��C?��v�Y���&c;�x<����5�ۂ���g^"Ze���ۈl�l���WMJ��q�Ip�G�,�ǈGQ�̦��S��,)r�K��R�eFW�D��ﾚ��m�B	�RT��mf���evf#�)�O�JΦ"�u/n�8ΧxX��`;�"���Ys�W0�
n�L��;;)�e,p�:ODf��^a"�����i�8"���Db���Y �LHD��M(#3�<�pvtt��7����,�Y]�<����C���ٱTĹ���z�X&��M�7V�!����T��I2V/�����c0o#j݌cY�KA40G����=g&�)��'+'����;��ˤ!�';���4�ѹ��M/c���>q0�'I�*��8%>��jT�)�N�^���7�t���B�'WR<�5%�j���gy�l�1̒ mG�o(��t"�B|���ρc0$�<�RQ�&�\�qf�/���Z�*�Ȍ#��'����8V��k��V��ۤ�[�/�g߯��
`�z�/����Q�$i���V��ڿ�:AC`ǨcR�@睇}�D��$p��V�Y�{ٱZ�ɫ_�鵰!��ϋ��[լM'A�DԵ�5����?Ϫ�yafy� �18���:��e�uW�L�	X ��ND]�Z��.OB���h5���XN�f� 3�7�KXcٖ/�ָ�A��Ѫ^����*�}c��{��r,���a�:���E�#�#z�I@�^�E�*|^��������S�\')Zy]`��6�z��=��i:y��[�f�#"�#�9:qD�a>����K��L�w�Z�U�����G�ҁG�'�u�Y7,�%w��J�0��yU����OB�cgg'���ɨȅ����<����-���o'�
|��Y,";��O�X{��(�$�C���I�?�:X��ze���Q-�q^i�i��V	�� 5����bc��^�^�Հz����?لߧ�K�س|!
U�Ɨ�3"��DT$Қ�>�X�U|��eN����H�noj�)�]_�*v �e}"��Q��_��I��A���U3KPY=GU�$��3���j�������+L�c�v��@���u"*2^�ꙗX�JlR�c:��6�Bg��9"T���:��u-��I�brh�E^W �a�AD�H��e��Qˌ�S���&��$�ÿ��?�k5��XIذv� "c�	*�ϩ��;��ÆI\{p���{њ#*%=鵬���5k~<[��{͖Cj���+r�:.�
 =� ��C1�{ar�	���+��֕-Bb<ݯ��"S����)����ǄS&g��(��O�X<D8E² GOFawg�pF��w����4�5(0/��"bRHN��&�z'�����@�j�g�ENi
"��*�u^��QPRA�|L���'�_��v� ״���^���c�v��X�I.Ք�P��(��ttR,�r�s�Z��6fV'���/O���jEZ�	�*�m���֩� �<��,�_ڬN/�X�{��c��8��1QU]T ���o��1�V�,y��:�{�&�@� ���9HDTS�J�Ji���R�q��*�h,����xy'����ۈ����_���c�ۈT��@���qw��f�8p�����Bu��K�?Fݢ=M�9"�]"���Vi���f���GR�"�:��7���6��8gȣqp����1���+�I�O�ٽΦZNc�U�"��F��t��i�Y��5�f=��F]m7���UZ�p8��!MS^2?,�I�8"RP�4L�r�A5� �f���*��@�������i"js��h5����\	��fK�Ѫ�jg"��D�&�9�k���\��3�WE�^ܣ,[���C�9ՌQ6�!2'L�bE����a�W6�0a���<I7U�H�UY����$��A̛|�1�sD#Nc�ӻ���~oB(�4�'��`���(�����B��.���xRȏ��;��V$�5ܯI��fJ+�dFVk���}֟�3���q��_��,�G�9Y���S@Bd���D�����'W���ժ�_��R���?��g��ly���Zc��T?4K5CN����|�2/Y�Q���ЍS� ���a@@#Es�T�k�7�կ^SI`q8GD�����K��;T�U∸'�BԵe����}d����ɩ"���&�mnn:3�M �U$"���x��t	I���^5[_PF�Y�0ΉJ4 ���W#���f��άS�~Q��L�i�l�z]�;�!>�U��Uԫk�.��ޞ\����kO���3m�<o��%�5F�;%�	���0��c<+���<f�U#��Xи栙�l!�(@�f�!A
�͑GS�s��BY#��#"�����N��+����h�X>��{͊�U{�n9]��F�f���ZYi������ۼ��Ā��b�x�R<�0vm@H��;GD ���4�S�U�=ǾQ�Xi<]%!h�3�.��H�`� ��+Х"� �'���Y�u���q"�G�l��0�Z�{�Ǌb�lEwD��:"&g��m�C�qD�z�͠��n���Y]�~A��c�%�%��:ʨ(�#���.���x�^$�q�I�a`?���$ D&GN�����x[��7�X	�-�-��!"+���`.S�e��P�Ώ��4MF�!�
�U65!I�1Gd�D��lMUE�T��_]P����'�6!�i��"
��^SR�;��5 �|�7U�����]u�,ī	$�{�� ;`A��)�&ZV-�LJ�b��/������aVf�]���G5FH�-�D^�40&�E��/�Q��:���tߗi>�Z@�2U3_0� �`�Ժ�xFǱu��M�����e���%������D����'����3P�QT=��k������I�9"�x���"�"I#퀑�G�PF���5�k�u�1ؖ<�+c��3z������r����V�%.��}�jc[������:�z��T
S�4�b\c�%"Ⱃ����y�f�S��̮�8����	�K��HZ�Ȭx�5�fv�50��#��e@�mY���#�R\�wOq]�F��4L�������Ҩ������SF�5j��������q����<�<M@R���d�)2:��8E<9::�G�=��0N0�0�j��s�P��Cޞ �4���Uti�A���r=�����D�=���G��ZHDMl��Hl�{؎�y��Q����)� 7)1q�F8=���~�La*$M�@mEDfYSx.�$̱��ګ�]b�8(V[��P�E��r�C��׬|�	J�3�SDt��	��dpxxHoݺŢ("j�f@��:l���͉Z���8f�@\���%i�$B_�~=��q2�]���J&nb����?�F�[DH���ޞ\�I�̨aJRR���<��ߗ������1rN���KŖ������-1aC�@0�� HjL��Qa%�A�M��q���O4qj��0x^��A,�b�Ȣ�0n
J�ԓ3�m,6����SOG��`<FqJ�M��Ęm�ahڄ�B���D$� ��������<�{�8ED=���'?��/���+������ͭ�8
�-t�$��6�f��0$����;I,^g)'���3��ѝw�����?|�C��o\�vs'M���~V��!R�	H��L�NņC\JS�^�������?���?|yLp����w�y��$�8��ч��q@!!p̓7k4k5�MGGG|4���~��/�;���n?��U��59ED�מ~�WG��b�sj���9�"�a��` N����<₈Ȁsv:I�s��	wN�\�:���#�<r	y��ox�7�Z��˻�����h�!�E�E��9���$1S�ǜ'������s��[�����+ڽqV���O>��p�o���vc�C�oJ�VHDBh�)�4��ؠ�A�Aͽ�;_>s���������K��M��	l<u?ϟ��1x��),�G}y�"_�߂�g>��3��Y}����{�+��
�h���*����$z���ŋ�̣Q4BD�w=<<V�s�����}�D����;<yxx�OD���I���� ��N<	y�9<y��P]�Q˰1�Ӫ���D�2����OD��������s�$��4+x"���(D�fOD�����t����5    IEND�B`�PK
     D"BYq���W W /   images/7c9bed20-c7d7-43dc-b689-820375f46db8.png�PNG

   IHDR  �  r   5)�   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{t��}������u�,K�,Y�K�6$�@�!�����4�%cH3�c�$�==s�G͜�4�9I�`;&�!mN��j�in��K�IHq�p3$˺��E�m����?d l,�'m�_k�%Y���1kyi���o�    �wy{�����B}.Kf��L���Um��To�jIU���^c��K3%%�L^#I.���0����r)/i���4��_�#2;t��O�u�h�ȥ���z0HC.�4���>�A��!�=��ߓl0;�9�,r��4�C2X[�����7��      ����+WU���+<_��bMII�BZ
fYM�P�e5&+X�5�� }���5~�ג̽���_��L��ߺ����rU���ܯ��
�^��_�:�[kX���ˍ>�Ҡ�!��d�2)5�I����on�|@���>I�if}I!�5����u,y�?X    ��b    e���\SSScP֤��(͒7e!4ɽ٤F���U/�,I��jcgOaC&fR�������i���������2;�I�-�,)�4wp$9�I������c��       �ޚ�V��$��4����nu.�s�!�2�u�LIu�>��je�)�L�kM�s�BG9��l@������}A��-y�{�ue=�vg
=-���(   [�  ���zݺƴ427UrJ4���� �u�)��Hj�݉�l��r����t��{�Bo��zf{<xo"ﵢw���ӱ�?v8      ��a^�����$�l��l�3�F3�-�F7�m�f�T+�L�f��I
��q�L�s�S��2uJ�ky�4�v��/Yf�z:n��c�   Sw   ��_S�/j~b�*��2͗Fo.�)NZ����}�>w�YP��vɽ�G���\}!�]�������Ñ�      �ym_�*f�s���T�z�T/��nj�L�f�����FN��4"�N�v��9���vȴC�vt�����۳ؑ   �d��   �N��k꫊vFf~�Kg���v�LgH����AIݒ:M�+��i��$Sg��d��ù���߸�@�P      �ܴ^���X��ZB��$���<�7K�d�l�ܚ}t�L�!�����&{:�=-Ϟ��t�7Wtǎ   &w   ���mkOJB�P���A�u�FOao���I;%�-�r�2e/ʭ+�l��v�;w}{�@�P       ��n��r�P�\�\�����[�B����u��I'I���
�}.=c�S�-X�M�=��q��y�8   `�1p  ��Ww������+���,;W��&-�dL3\zI�n�~-��z!1��S�U���Eݵ�;      x��6$IOk��TSx�����N�L'K:I�I�cg�ߥ'��qW�.��L���X�;v   p"�  `J��~M}����ȃ-�k��s�϶��2�OҎ#7��w�n���C�������     �i���5����[�|�曍���*�4I�q��Ϥ>���|�����oݽq�vN{  �T�   �V�u�GJ�E��"�](��}�X c/��)��_pٯ��7�*��М�ya[�ґȍ      ���6$��:�,���N5�i��ͤS]:U�<I�ȕ@Y:<zT����$���{:V��   8�   �.oϵ�n<�C�ăs2;0)uJ�&�w�iGRʶ�����~�^�     ���7��id�/��|�1_N`&�Nwm5�&ۜ&?������    �B   ��ᣫf&���`饞�e2] �2v���(�yw=mf�����?J�3���}Q��Y�@      ���ew�*M�H��p�3�~��ΐ��X/0U�$���2e�,}hw��=��   0�0p  ��hi[Ք)���/3�e��SR�����Y����s�BxƇ���+�c�     ���]���"�s<ՙ2;#Hg��t�ΐ4#v�q璞��!s{����{��;cG  ��1p  ��h��Wk�ʡ�%-q�ȴ@��	���H�M���-H�=���}�'�b�     L'uׯ�/}a�-��B�-��@Rk�6 ��i���ɥM�$ܿ�影�   P~  `l�mH��.3-1i���$bg���������k[�oWjۺ6�x^2�     0U���g��o��ۂ̵Ђ��6� �V�vH���&��������I   ����
  ���a��s�}ȥ��~� ��^���|��m�m�R��ӱrw�0     ��d^�W����������/�47v��6$�-�/����q�S��   051p  ��;|J{0��d���gJ ���ɷ�m[&�^SS��_�q(v     �xk\vGk��E.-r�E�Od�� $=/���;������o�  ���1   �P�GW�̗�t�Ur�+I�c7�1��]�c&L�+����;     �h��WkC��yJ�;�]��N�ΓT� �A��Mf��e��������A   ���  ොt������g�f�ߕT�	 �H��m&���[w�����۳�a      /=�=Y ��l�\�$�-)�n�1�I��K�V���x�3��   0�0p  �$�a�ꓓ,\-���t��$v L��r=������,�Gzf�'t��b�0     P�����'��J�p��_ �&�SRC�4 � n�[3���4�枍�;   �1p  �ƚ�V��Z7[&�"��! �lH��dz��	!<ҕ�~RK��a     `�rk�f��!I/ti��.t�I��� `�pm3�=r��]�\�   ���	  `����/�*T>왵���%�b7�1b��oq��P���}R��Y�0     0�4.��5��"���"3],�1v L!�]�[��{�߶+v   &w  �i��<4���p��_RE�& (\�j�G�푐�#]o�;
     L��mkOʅ���Å&]��cv ����#�}�S�b  `|1p  (c�׮���o��ZI�b� �4�W�Gd��+�I�Xz��o޺'v     ��jmR1�;R����Ã���� `���[��k���l�6  �w  �2Ӹ��$m.��2�#v @��i�f�oɤ�s���mKGbG    �7�|͚�����Z�E��-)� �]&�{y������  ����  �,l�P��h�n���$%��  o�d[M�c�~��?��X�;v     �]��k��.6��$�X�E��1`*�b�w�r`}����P�   ��   S�춵'�?��Ҥ�c�  NH����FOz���~䅯�8;
    ��ն!iɺ��r�H�K�Z,�lI!v �-; �z)�����b�   �a�  0մmH��烒-w�J�d ��a�&�G�m�����+�cG    0U5|t�̤��D��ʵ�LJ�� 0N\)غ�����o��  �c��  `�h�z���&�>)��= �(�2���l�+��{�O�    `�jX���|��>z:��2�+��W��-K�vu��|�   �9�   �\cۚ��[\�IIU�{  �J��~*�f�o��O����     �U�5k�{�ktоX҂�M �I%s����wm�eS�   �>�   �Q{{h�>������!�s ��HzԤ͒o�{Ŗ���;
    �1wӺ|c_��D�Xf���I��  S��Q��TUS��/|�ơ�9   x5�R   �HS��
v�I��uF� ���Jz���<<$���X�;v     �k�G�8��P��e�I~�d�$bw ��N��$I�]�,�  �Q�  &����sv1o�Iv��ٱ{  e̴C�˴YJ��q��     x���UMn�Œ]"i�K�K
��  ekX���e�gwu,�u�  �鎁;  @Ds��r�ґ��{Iu�{  �R�I���dY�e�ƕ�%��Q    �饩mu��]�Kv�K�� �(�������q���1   �   D�|͚�J�߹�&I��{  x��&=$�-�lsoǊ�1x    ���ew��'���D�Œ��_ &w�wC�g���'�c   �    �@�׮=W���5��t SC�\��f�@�9�W{{;
    0�4^{癉��\v�K�3���M  �M���=+7�  �.�  L��׮>'���\�KJb�  pJzإM��Ի��Q�    ��z�	�ҿ����M  ��-!���{���  (w�  �Q�5k�{N&��Ű P�z���L�ݵ��c��$��Q    ����A���$��	 �q�%s��ގ[�  P��  ���k�<3���d�İ 0�x����d��e��ގ[��]    {�V��s�_
���b� �fL�nB{�����  Pn�  �����5�i����)I��=  ��]&{P�[R�fNx   ����mu��]z���Œ�n `2p�w��O�l����-   傁;  �h�誙I1�'6:l��� ��e;%�ߥ�����]����E    ���Ҷ�)���u��+$��	 �I�(ٗ��>�}�'�b�   Lu�  N�M���}�n�ɚc�  0�vH�$��4���c�K��    `:j���k4\�IK$-q�|I!r  S�!�����u,�;  `�b�  �5��Y����\�c�  P&\���t��_̧����bG   @9�����bRxo��+l��%�bw P&�e���]=w���1   Sw  ��Դl��������-  ��Ԥ���އ*��?;
    ���I�z�e�%6zJ�bI���  (sO�§{6����!   S	w  �ct��w�.��/\�RR� �i�d�c�6I���n�X:;
    &��k��W�������f�n `�ڔ���y��'c�   L�  ��M���}�[��/%���  G��c�6�kS���G�ޞŎ   �X^3h����M  �����������Ď  ���  ���k�\i���tf�  ��H����OK���l\���A    0���>9��
3}@�+$��	  ��N�������u�<v  �d��  �(�h�ܐO?'��b�  ��ʻL��\���]�=�    NDK۪�4�.�%�ĥE��  �[�z(dي�o�;  `�a�  �J��yۜO���f��  cȴC�˴��������w�N   �7�����h��=��HZ����B�,  0v�&_���CO����1   �w  ��Z�־;�I��c�  �q璶��~��?<\|`߷>�/v   ����uեJ��Bz�g�~�I���  ��yW��g��ߋ  00p  �^}ۺ��e�Y���G  LW��?���٥V�qb   ��v���*�׆�Lv�ܮ��"I��]   ��YHo�]ۮ�!   11p  �Zӵk��k�I'�n  �Jj��%m��)�C[vv|z0v   �)�mCҨ�w�i�\��t�����  ����\�ձ�˒y�  �� �ii�G�8�PQ�9�n��  ���I�����`�g��p�(    �_�5k�+h�LK$-q�>v  �
�A���=+��]  0�� �i�y��\�V�I�[  ��5 �G.m������úky1v   ��^9hw�
I�c7 �)k����,����۳�1   ��;  �6��^;�����X�  Pv�%�ĥM��Ի��Q�p   ���ew��'����]W�tr�&  Pv�d���v��T�  ����  Ls��^-�$5�n  �B���i��6�v���d;
   ��kj[ݢ`���D�ߕ���M  `Z4�?��e�5 �r��  ����6T�7�n��  ���&=$�&)�AW�m��   plZ�V5�!wyp_,�%.] �g  ���W��7���mW�  ���/  �l5_��bw}]��[   ^�Ӥ�rm*&����W�;   �����3��Œ�HZ   LB�r���c�7c�   ��  ��u��}i�I&)��  �f\zҤL�`Z�����坱�   ��b^�W�a������z�L�bw  �����P�������  0�� ���x�g&�ΥE�[   N�Ӓ= �i���X�R�    �\�^���T�.5�.w��$�'�  `�2�0ˮ�Z�ñS   �
w  P6�,]{��_�4+v  ��4i�\���]�=;   �*Z�V5�%Kv��%.�/�  ���$�l���Ϩ�=�  p�� �)�����n��  0A��-˶��x��A   �d�|��9�g�b�~�x^  L�������Ov�  8<�  ���׮>'u� ���-   ј~%�.{�ݷ�v��T�$   `�4,[}r��e��R�]f�9��   ⱝ��u=+7�.  x�� �)kε�����H���  0�t��2m���9j�鶎�#��   ���|͚���Œ]"�bIb7  L2%�?۽��3jo�b�   /�  `�9톻+׸tc�  �)⠤��9S�`����ΎOƎ   ������E��K$�L�Hj��  0E�c���񉽱C   �w  0�4�Ѫy�\n��w�n  ��J&=&���lsa$���o޺'v   �zպ�be�����f�TR]�.  �)��Y�������!   Ǌ�;  �2���^���%5�n  (3�\O����m.����w���Q   (-m��\����er[,���   �̀�n�w�7b�   �  `Jhn[s���On  L�Nwm�i�ܷ��T?���n�  �)�mCҒu���l�4zB��s�s�   �tWw]r��Z^��  �Fx�  LjMm�g�W]�4v  �4W4��o��6[�?�}�'�bG  `�j��Wk�b蝲�1���+�!v  �4����z:V�  �z� �I��m�)%�ߖ��[   pT���ce�c�Qw���:����   ���k�:+���f�r�L�H
��   �j.�(��t��y�  ��a�  &��k�\��ߒ�9v   ��AIK�c7��H�����[�bG  `�5����$�BO�K2��fz��ٱ�   p�I����|+v  �k1p  �N�ҵKM�5IU�[   p�:ݵU��r�R��;;>=;
   ǡmCҒu���l���l��ߑT�� ��2����L!��f�p��LLvӚ4s��Us�2�X�����h_���{����!   ���  L"nMK���I�E��  P�J���i�e�5�m�]����۳�a   ո��$�\Z$�%��+�:v `zI�)I���`JB82NO��8=��瘤p��L��� ��Q{����e����fGF����R�*����Uʲ߼���,S���>0�\Z_S]u�_�q(v  ��p  L��pw����W$�h�   L�~I��|�����oݽ��m��   ����uu9�Γ�%r-6ӻ%͉� (fR.%IP.�W�����z���=��|��NTǨb)S1�T,�)��_�u���X�8-���#+��]�\�;  �{   ���UM��#�ݱ[   0i�ۿ��O%�txd��}��Ծ�Q   SY��>_�U�o�w��wL�H��bw ����M�$�'A��G�|?�>=��f)�I5\L5RL5t�-�w���<W�l����!  `zc�  �jn��mn�?J:3v   &�Nwm5�&m�\��ӱrw�(  �ɨᣫf&#�;��ȃ-�k���$%��  �K0S>��咠|��%ʽ�����z�d��0R�4\,ih$��HI�#%������U�ׯ�Q�  0}q�  DӸ�K�,��dͱ[   0euJ�f��n�J�u�ƕ�%�)Y  0m���g��s_3f?[���4̔��'����dt̞O�sA	�uHr������)ip����"���됙-�w�wb�  ��{)   ��ew~��p����[   Pv�Kz��[�����}R��Y�0  �ո��$�\Zd�.-�� v `�|��o��9q��J��[N[ǉ�2�P������h`�����t��le��+��  ��f  ���s��-��H��n  ��q@����gf��[x�nq��߿}8v  �Q]ޞkij9ӕ�'��]~�d�Kj�� ?fR>�9u��O��/<�t �,s��th�ݻ�    IDAT�������F8���d�W���)v  �^� �	5g��?����!   ����3A��\�P�'T
�wm\�d<=  &�춵'%�s��2;W�Εi��B�6 ��yy�^ȅߌ�_�>�=�0^�ԑf��������R^<��}�{A�J^!  L�e  `�4-]�g&�U�   �M4�i7mw׶ ��I���|�+v  ��?��ZU��/4��k����dͱ�  '�L�%��r��_�z��+w��PQ������{Y�{�g����c�  ����  L �9K���H���%   �[eR�K�M�Un�2���P�g���| v  �d.o�5Ϟs�_��"�-pi���%�n�)(	����_���Q;�Q���������e��w}����텯�8�  �7�  `|�mH���.����)   �8(�􌹞4�Sn�� =9�K�����Ď  �k^���UqV��r�9nv��Βt����} �c�S!��"�(��'A�|2:^��u�-K3׾C���?���R��	��U\���?9�  �/�  `�ܴ.߼����li�   `��|�L�ܵ#ȷ+�m]�u���v^� �)���5������m����Od?KR9 �&���8i�ho��0�ճP��N���i�W������!  �<q  ���n��rp`��]�P�   `��7�)7=e�oϤ����j���g�;�� ��������tN��� ���96��>v ����������|�p�:0�����?���!�Ǯ��ʆ�+TΔɶ&I����Y��	  ��  `̝v�ݕ���L��   �BRI/��K7=�rNY�\�l{Aw-/� `�kې�${Nv�oW��fo���n:Ǥ�%�c' ~[L�|��\�B>yՠ�"�(	L��h�����C�)ĳ��C��\�BU����\.� #w  0ָ�  ��¶�n�n4��n   ʉI}.m�i��vȴ�3�H�<�ױ|�>  &��m
�Y�<%�/�|��K�7�ΑT9 �
I0�s��i�Gy�O��ePֆFRu��ׁ���)x^T64�0#w  0��  ��v    ��$�8r;<�W�]�u����,r"  c���5����[���b��:MR�� �����$(�U�GOa/��s��`�����ۯ�b;�#�//��I���Y��\�,a�  �
w  0&N�rU����>�}0v   �W9$�s2�0��]��.�hn/fI�W�g���  0�4��nI�Nβ0ϔ���N1��=���f�n H�L�\���[N_p<ܥ�}�Գ@�k�j���G��<���T�Kf?��%/}��=q�  @9�$  8a�6z��C҇c�    8nEI�&풴C��L�K��i����w�����2 `L�v�ݕ�[�h������#'�K��N�4#r& @����_q�zE>Q����\��|;@�.���9�}�҈���G�MF�  `�1p  '�u��}�F����   `��K����^���,�Up������������"7 &��n��r�P��,I�Y�S]:�d���3;���\���	 �S!��"��p��z� �'�\/���ރC�S ): /���?GF��g##C���O훸:  Pn�7
  ޺��д}�7LZ;   @tC��Lڕ�:-h��;�՗ۥ�;Cf��f'/���ر ��3��UŬrn�U���[e6�M���>������-��' �4��|N�|�B.(����|d��`
�=0�]{�弶\Ti��or�~R��z����˗�t�쟘:  Pn��
  �"�9K׬�ly�    S�I}.u�� ^��L���;�m��Yg)�}��o플��`��v�ݕ�C�J���y���y�I����Ms�:YR>v/ ��^>����Se>9<fOT�O8�@��,ꅮ�J3&��Ӣ��=���GF��f�?���o�:  P��7  ޒ9K�~N�?��   ����k�I{M��f{\��2��=A�׃�����|޳[-{ձ�M���s��w�	����fg�}�)kp�l�$k��l3�vi��FI3bw �]0Se!���÷ÃvF� �������ܯb��N�v��C�������T���d���Z�  ǋ{�  �5/]�����    �:�IꕴW�=2�k�W���{C�=�|o�'-%�ܭߒ�A^6@l�W��Ns�����>ە5��l�7��`�l�7H6[R�F�<� e�c�ꊜ*�9��憋��۵���K�J��q}���}�L��kÊ��*}  �xp�  �9׮�En�cw    �8��'Ӡ|�}w�Ӡ��̽ϥ>s�I6����՗��\6�˲�R������mK��_ SҼ�/T�WV泴*W��4X}0�gf�&��L�n�7Y��UnV���ToR�KU��5:T���� ���OTS�WMe�1; ����T�u�S����I��%?�?o�U)T�����w�m�  �w� �1kn[s���.)�n   �)����2;$WѤ�L�L�/I&�IRf:`R*�C&q������((�^��,�3�\!;����>��l8ͧCŐ�6`�������3�(Kuׯ���
E��U��,�,�*	�d�,IrY��I3B���U�Y��*�T���j�f&�W�LA���.U�T)W����7  �[!����pd�^��; ��ᒞ۵O�s(���lt��Y�Z�r�L��]n��ǰ  �1�  ���,]��L���
�[     'lĤCG�����[�xwi`��P��U������f�Q��p�Rz�� `
	f��̫�����U��I 0������bg�=�J�������Z�B��tcφ[�f��  @c�  �T�5w.�$<�/�        �De!�����TU��xv ��K{�ջ��^�c�Ӣ��='�}Be�,_U���+��� �2�]h  �������ǒN��       �de&ͨ,pJ; L�,s=�R���i씲5VwI
U�d�ʃ�}=�W<:&�  �%�  �u5|t��\1���w�n       `�yy�^7�Bu��;	 ���ᢞݵO�Kʓg%e�z�軙BU�,W�LJ�{:��Wc� @�a�  ��u�9�Jߕ�wc�        0�̨�k֌JF� 0I���מ��3����%)(�4H!�d������1��  �LpO  ՜��W�       0�"����Fg�ܠ�ϝ�ٵ���`�h��V8�s<ؘ���)�yvN�F�[ض�0�   e ;   L>MK���\��       @LI0��V�~F��+�s  �#�5�U��o vJ��q��\�*�SR�𾞰g����"  `*Kb  �ɥi�>h�/�Wz       LSU9�4�蔦Z��T(��u ��*9�90$�Rn��#����z&OK
��w�X����}�'c  0U��<  ����/-�,�����[        �H�FOko��Tu/� Sѯ{���P쌲���H�����|�B�����������  �)��;  �$�^������5?v        %�j�Y��3���B��l`��g^�;�줇�HYqܾ��)+T4��vݻ�q�  �2B�   0	ܴ.����3n       LU9��T�sN��9���@���+�c5�l|�L����p���CK۪�q�  ���  h���.���       ��V[U�魳t�I�j����k��RWS;��XH����~yVz[j�{uy{n�/  &5�  LsMmko���;        O�U�q�,͟[���|� �8��*�N(?�|���L�@�̳�ϙ��_'��  `�^  &��k�\,��3       �L��T��晚3�Z��@�K��g�`��⩼4<��%�|�{j���Cۿ��	�(  ��x�5  ��9�}�Yi����n       `��V��P��
Nk���/��p1��Q6<-*�3a׳�������{W<1a  ��D�~  �l.o�YZ��q;       ��TW�����4n�v ���
��	e��ľ���ˋC5.���m]݄^  L
�4 �44gN�_����        ��B>QkC��j*b�  "��8�sLY�y6a�̆�+��|����#���]  D7���  D7g随H�ג,v        '*����F�4ժ��3�  �p)�����e�KÒ�|��|�Y�64����'��   *�m  L#M�|�K���jc�        p�f�Th��*pR/ ��֯���(+��yq`�/�T(��O3�z;ny`�  @�� `�8��U��z1n       Lq���No��S�g2n ��$p��X�$��鰲�CI0}���u�q"  �D�>  �����J~A�        ު`����yR�j*#�  �^0�c.��]���FN*�ҿ����  LI�   0���|���Zw�       SҌ����R���
�[ ��R�i����e�,�G$y��{:�P�:cƹ��?��{?�  &'� P��hռ`�1n       LA�L�j����T��7 ��K�8#첗��]�S�����5_���x!  `"0p ��]ޞ��r�H�; ����;��,����;�n��K/3==��R\d-�,QR$[�I۲�CJP,[�DQrl�p;�3�_�9�a�A����ț ��+��Erv���޵޺�9'/zHΐ�TwW���{�h�@�C9Uu�{   �v�tZ��=˱:?�:�1p?Y��6��G��mUU�O��YL 'w c뛛OFď��     �ۑe�Wf�3��p�܏G�{DT�ݨ���Y�[ ��c� cj�3O�����     p;ڭF<tf96�f"�R� PG��0u�X���	QlEV���x��_N� w C����g�����p�    ��X���#g�c��L�@��E��e��ܫ"ʃ툪z�̅gΥ� ���; ���?����Sw     �adYęչ8�����v �N��c�5;�""�D5�.��œO������ ��槟�dVů��     ��h5�x��r�/N�N`���ckT���NT��'7����S�  G�� �ș�>�VE��Sw     �a�N�⑳�1�i�N`L�t���Z�hEd�29+��nE����|���S�  GgT��  ���(���S�;     ��,�OŃ�����kk ���~/u����s�=�A���NUV��/|��: 8� ��X����BD���;     ���Z��s��e�K '�A��Aꌱ�5Gh�U7�r��+ٕ��� 8 �X��ԩ<˞�"�S�     ��ɳ,�m����h� ������3�_UF�{9u��e�ḫ˼������}� ��� c ��)�v     FY#��Ӌ�� ������A�ɐ��vꊷ��({;ͼ��i��3��9 ��1p��[��ӟ�,~!u     ��V#�N/�씽 �����eꌉ�5G�k�`?�����7ʿ�� �;Y�  �Ν�s_\���Dd��[     ���[�x��btZ��) �������z=ʪJ�29�"��+�+�Wֈ��Z/����x�sϥ� �� Pc�v���    U�V#:�d����������7"��߫*���vʬ�'�䓶q PS��@M�?񥟍*~%u     ��v��^�Vӯ�8>�vb{��:c"�ͩ�	���EU~d����L� ܙ,u  p��>�{��T�?FĹ�-     �ݾ5no�p���a<���(J�ۓ��(v�D���?kDcvm���_�7^I� �O ����ޓa�    �j5�x�Ԣq; �jX��ҥm����<��N]�Ϊ"����0+�a� ��y�  5���ӏG9u     |�f#�O/E��H��+�*^���A�:e�孩�	���GU��槟�d� ���@�TYT�#���     �*ϲ��Ԃq; Ǫ,�x��V�R�Y�Y�wQEy�Ud_����?�� 8<w ���O��_�"~<u     �U�Eܷ�3�Y 8>ߺܾ�5nY���}D����se�o�N oT?> |�{.���~��jD��n    ��:�6kө3 c�a/^ڊno�:��R{Qvo��xy4�V��<����[�� x.�@M�����     �����v ��~o_�q��ʚ����:�=�Q춋*�݈�AX ��Q�� x��_�������<�f�G#Ͼ�����Y    �6sӭ�w}!2O�8&W������(J�'iUQ�SW��rY�u���������?H� �7� `�=�d���ƿ��L�^�e1�n�T��V#��<��F��y�y���h7�h6�h�ydYD����������UTQEQT�����3��c0,�7(bX�'��   �I�j�����h6�8��7��ͫ;��?£i��,�ػ�����ḫ\��G�����v� ��5S  �m�+��Yd��0�ڭF�M�b�ӌ���?S�fLw��i�˒n��h��_bn���������� �{����c�7���A���   �ۗgY��\4n�X\�9����𩓼��D��%�F��n6���""�v� �ݹ� #l��SsY��QD�I����g1;Պ��v�O�cn����h5��˻��b�`7w{��ߋ�=�w    ��=��:?�:�1�����vc�`�:�;P���L��>�ḫ���co���|)u ��\p��g�ߪ���DeY��T+g;�<73혝z���u�ȳX�i��L;"�#�ֵ���^�����^/���QVU�P    F��lǸ�#��q��^\�9H��]Ț���Q�S�Ceow*��^D<�� xg.���ڼ���s�p�y�3�X����ܭQ�8\f?JeY�ͽ^\�����.�   L�V#�G�Y�f�34 �^Xƕ����}��Θ({�Q�wSg��|f5����+_���� �^� 0�6>����/��q4�i���L�/N��\'�̷ŷ��ƕ�ݸ��7w{8   L�N/��t;u 5w�/���~��=�f3U��y+3����� �|�L� ��% ���O?��DT�&|��#�l䱺0��ӱ�8�V#u��e\���_��   `̭-N��չ� ��N�W�����O��1*�7���x_��bDk�׮|�7�i� ��� `�T�槟�wU��S�@��[��\����X��J�3z�".^ߋ7���N׃i   �q�n5�ѳˑ�~����˸�s�w�?(R�p�������/ˣ1�~1������7�R�  ��L  ��槿��*2�v��fK3qjy6V��OZ�Ո�q~s!�q��^�vm��j   �1p�ڜq; �V�Ul�����A�v�s8aY���"��k_�Q�wO7��߉��6u ��@ �(��gZ7��"��)P��wF�F����tc?^��7�z�s    �K���os!u #nX���ߏ�^�t�QU��H�t�<�J�qY4fWw���Х���S�  ��� #d�F����a,̴㞵�8�2��FV�eqje6N����~?^��o\ߋ��T   ��,�ӫs�3 AU��c�ۏ�� v�����5�ۉ���)��7�M-�͈���5 �-�@ 0"�/<5�e��#�T�U�F�W�➵���j�����E�vu7^���A�:   ��pfu.��Sg 0"z�"v��ߏ�n�A�S�ۍ���:�P���~#ڏ]���!u ��; ��,��zDe��`i�������Ld��h�]�و�O-�}��՝x�Ҷ�;   �j���`�0����no��A����0�A1�׸%yk:��^D��!��^��i���R�  .��H8��gֆE�|D,�n�Q�ek�q���X����UU�_ۋ�/ތ��;   ��8���s��L������3f���q���b�ݭ������O���h}�ʳ����n�I�; ������̸"��gqje6��X�٩V�N@�eqvm.ά��   ���vӸ`UUDoP��`�~�a�E��E���_�<7�    IDAT٦~��lm�eo'oή���S� ��s� [��?:����#b*u��n5⾍��gm>��<u	�e/_ގ�؊��0    ��O-��L;u w`X���1������c0,S�1����E?uơ�SK�Ο���o���[ `��� ��U�o�q;������b�[��<��K"�<��O-ƙչx���x��n8   prf�Z�� #�,��U��m�6f�����۳Qv�1p/{;�hN������[ `�Y@B+�y��f�}="�畉�j�qn}!��\��a;�ag�_������K�   08���� ǡ,�(�*��֟���(�w��o�{�)uV�]�(�3%�Z��L�ؕ���� &�� �P���V�3aZ�<��\�s����L;��#���{��nDoP�N   [S�q;0V�5/�����[���u@^|���|�q�w�΋��*�����?��n��:��$��3Ql��8������߉��I� �ʢ 9s�sì�Z�3!y�6���B4y�j�(���k7�WvR�    ��{��ce~*u�����uɼ��E��ͫ�e��ۮ����[����ؽQ�㐑+� ��� ��0���̸����8�޻�m�~rwy�ݻ��g�W���A=^e	   P�F�s������9N��7�g�a�a���X�-��=U�G�n]q����ө[ `�� 	�y����=�����v<z�J,��,G�,�x���x��׺   ��+���4�:3U���������[#v�xaBT�+�Q�.9���ў��+_���� &�� ��0/�����_�f�Z�s�Scy���g����\|�嫱��O�   P[y��ʼ������h�[�ް������ ""�<��tT���%�R���њ���n�I�; ���O�md��z;c(�"�m,ă�����V��SUU|�������)    ��4ۉ�6Rg #lX���o���"E�C؁ë�(v�DD=�Ƒw"k�����~�ߦn�I�; ��FV�NDf��ؙ�n��[������eY��]��������FP�N   ��e�ہ�����������K���%v�dyd�����%�R���ў���[ `�8�	 'h񗾴���1���J�eq��Ÿ��Bd�o/I�?,�?�t-�m���(   @j�F��[��`rTխg��A�a������'�*�Q�]M�qh��b��;z�_��WR� ��p� NPg��vDe���X���έ��T+u
|[�و�=��\މ��v�/c    ���\Ǹ��;���8���dy3�щ(z�S���f���_����� &�� pB�|��t�RD��n���l�����gm.u
������/^�ޠH�   0��g9��n�A��2�Et��[\dFXU��ܿ�:���A�9������+�[ `xJ 'd0S�ZV�S���x��Z�t|+��[���}����^�[{��   p�ڭ�q;��`X~{ľ������C@�d�vD�Q�S�J��k[�5"�Z� �.��I�ē͍���G���)p��,⾍�x��r��mUU�s�\�ׯ�N   )k��qv՛aTUU��"{�7���0Jgف1P���L�qh���~kj����߸�� Ɲ���	����L�ScS�f|��Z,�uR��ɲ,>x�j�O��k�]�J^   �7-�x����"z�"�{��ڍفq�5�"�fD9L�r(�`ofؚ����oR� ��s� N�慧�]�e?������L|��j4y�8W���/^�aQ�N   H��g����"�[c8qUq0�5`�w��`ՠ��V�C˧W�v�o>�׺�[ `��� ���g��DYV���N#���V���l�8Rk�񃏞���rt{��   p����pB���W��{��;DQ�d����NDU��D�`m�X������- 0�����e�WR7��j7�#���L;u
�٩V�ࣧ���r�t��s    ����GUEt���;�Θ}0��p��e��f���9�jxU9�;�?��|R	 �����1:���ϗe���h�n��Z[���_�f#O��nX����_�����)    '���]�N��k�[�a{o������2y8���b�jD���@Yk&�ş���o��[ `\�� Ǩ(����S#�7��˩3��4y��Û�^��o��   81�Fn�w�7(b���A{o�a�$�z���ZSQ��jЍ�3�W#�� ��� pL�>�{��T�ՈXL�������Vc}i&u
$��+�⵫�x�%   ��Z����ͅ�0�*���y�}����0P+e��Ո��+0��|��Ǯ>��?J� ��w 8&��ޯU�q;�o�ӌ�>��S��)��έF���˗�S�    ;�᝕e��a��c�;�noeU��%@��ȚSQ��K���g����#⯤n�q�; �'��7���ZD<�:���l'>��z��^E���oƋol��    8V�]����;|�B�n�֠}�``��HU�ܿ�:�����as����_,�s� ���n�\�q;#mci&>t~-��g�:�a�   ��,��n�3��*b�wk�n�0Z�F+�ю(��S���ϵ�S��0u �w 8eY�Ff3�;���޳�:F�Cg����x��v�   �#�n6�3l&IoP��� v�����GQ����=e��(Q��ET_��|q�#� ���<uo��^��F��nY��=+q��|�����z=^���:   �H-�v���B�86â�݃A�9h��I ܆b�jD9L�q(Ys*bj�W������ Ɖ� p�e��a��ʳ,>|�Z�/ͤN����{W""��  ���iy��x�����A�toڻ�z�"xgyk&�^=޲[{�W��"�� ��� p�>�dscc��8�:ު�g���cma:u
��W^��_�M�   p$�]������pW�E���o_i/�*u G���ػQ����~3���ҿ��˩S `\�� Gh}}�φq;#��g�7��
���[�aQ����S    ��T�w��_��~/����w0H��qɲ�Z3Q�kr|��m�ss1"�^� y�  'Y�K� o�j���7���|��Z,�vRg    ܵN�4�,����ūWv⹗��}�z\��g�0��LDd�3�*"��'����#�* ��'�y0��'Sw���y|���X4ȅ#���6�٩V�   �;�gY4�ŘHEY�ͽ^�re'���x��v\�9�AQ�N�$eyd����7����� 0.|4 �JU|.j�r�]�Ոxx��X���Gڈ��ވ��H�   pۚM7�=â���~l��b�ۏ�J]�(��3Q��3�D���G���� Ɓ �O<����x5"N�N�V#��?��3��)0�v����R]�   jf�ӊ��.�΀˸�׋��^�R� 0���ke=�Nd�a֞��ʳ��F� �;��#����sa��h6���q;���v<~~-2   j��;	e�w��7��_��_�5n�=���	�V��,�_J� ��� 8U1u4�,>��z,�ÉX_��O�v   �K��WĜ�������+Wv⹗�ūWvb{�U���:�ZSYM���(��_K� ���A �Kg��W�����*&�<���\�����)0q��ū�ƍ��    �rjy66��s	������v7��zQ��� ܹ��U���ɚSSK?p����?�[ �Κ� ����W�2n'�,����k����[��� ����S    �W����񩪈��^\�>����e ��5EM�հ�j�"�� �BM�� ����WS70�>x�Zl,����y~`=ZM?^   �/�o��eW���\��/m�p��ƭ��PE9�}����B'u	 ԙ ܅�'�������L�O/����0�������1   0�2�/8BeY����^�ׯ�Ơ(S'0��V}�f]{�[�O�� �:3p��Ш�_M���:�:�^L��ii��YJ�   �|@��rs�_����x}/��� ��َ��3�D�)u ԙ�; ܩ_�UE|6u�ii�8��:�.�7b}�>D   ��c������k�݈�/m�`h��I��v����/<u*u ԕ�; ܡ���D�Z�&��T+>���W	È��}k�i��   0q\p�Ne�^ى�/ތno�:�	��j��mD��; �����Y�z;'����#nD���8U�f��54    �ƍ�^|���q}� u
 �,oD4ک+�*�v9u ԕe ܁��Ϧ"�O��`��Y}p#f:��)��X���N-��    �eU�N�F�E/]ڎW.oǰ(S� @���ǰ���/<�P� �#w �{������L�G�Y���N���8�+�S�3    ަ,�9��n?������K� ߖ��"�zLުa/�j��� p��� FL�B9QgV�������mz��Z�~�   F����x}/^��W�9Ydͺ��~9u ԑ� ܦ�_��BD���L���v<v�J��tZ�x�  ��;�?,��ߌ�7�S� ���Zө�����>�� ��� nSc��ň��G©�V#��p=�<K�ܡ�+���4�:    "\p���t��o^��� u
 ���ъț�3��E\q��e� �)�곩�Y���k1ݮ���]=vn%Z?~   �.���lu��7�����Ț��IW{�Q�h ��� né_X��O��`2�j1���z=�ݵ����{WRg    DP�N`�TU�k�v��k��? u���3p���{6�x��Rw @���m��柉�9v3�x��R���Z������   ����󦢬�K[qu��: n[�7#�V��)�Q>u ԉ�; ܆�
?tr�y�=up>pn5ZM?�   ��e�F@oP��_�����) pǲf'u¡�E�B� ��
 8���,F�O��`�}߽+1�� G�f��]N�   L�����'�~o�x��k� �^֚J�ph��ྍ'~��Sw @]��!����N��x�X��3�s�3�ctfu.�����   ?��a���⅋[1,|�����fD�J�q8� �����3 �.����|� �[�Ո�[M�����]�,K]   L���'��^/^x�fe�: �Lͮ�� �!��!���33�3�;o��_�Vӷg0	f�Zq��B�   `B�R'p�n������Qٶ0f�f��E���_z4u ԁ �`�����I���:�6+��y�ܽ��,E��H�   L ��ru���0��FD�L]q8E?�j�; ��; F��:���n5⑳˩3���3��   ���e�N�������� p��f'u¡UÞ�; ��; ��^�r;��������]�f÷e0�N��z{   ��+���ҍ�x��^� 8vY�>�(]��/ܓ: F�% ���������������X�I�$��=+�e�+   �Ic�>ޮlu���Y�u��U�^�l6�t� u��� 	�?�����l��ع��@bsӭ8�2�:   �0;]�que��_�M� '(���NqHU���O�� �Qg� �#��9�]�N��:�Y�F�;   pr��8��38b�� L���I�px��'�|�����`� �a��*N���Y���=k.6�tZ�8���:   �0[{��	!�v &Y֨���j؟�w?�� F��; ��<��t��ӣ���N F�����   �	�i�>6���xy#"o��8�2��}*u �2w xUT?����sfu.f�sA 8�<��7Sg    �?��~�:��t}��� ""k��w��p��U�� F��; ���_��B�;/�<���,�� FԽ�s1ө�u   `l��^k7v{�ͫ;�3 `$d��ܣ�����J� ��� �Ec��Saeȑ���btZ����ʲ,8�;   pr�mw��RWp'��z��m� �MY�F��/���I� ��� �E�ϥn`�L��q��B�`ĝ^�u�   81��������nw�\�1n����>�c)��ϧn �Qe� �*�����G�.G�g�3�����    '���~�n�~o/���u; |�z]q/?�|����w`� �`����I���X�����L��&ά��t��:   ���0��38���0^�h� �&k�S'Z5�7[1��� 0����T�O�N`�<xz)uP3�o:�   ��+[��	��n/��Ei� �Q�Be���Ϧ� �Qd� 2w���l'V�Rg 5sv�w   ��l��\qa�A/^܊aQ�N����͈�F��r�S� `��9 ��^�r;�������κ�ܙ�   '��k{�x�a�_��v 8�����Ъr���t� 5� �]�Ƶ���������X�s��3gWg��j��    &�~o7v{�3x�aQ�o�`h� ��5�3p�r�p�'Sg ��1p�?�:����i�ہ;�eYܻ>�:   � ��FYV�3�[���/nEoP�N�Z���	��,����w�2w����t,�uRg 5w��|4�,u   0!�2�luSgL�aQ�ol�A�: �'���=��'��� ��� �����j�����N-�N �@����չ�   ��ts/����e/��ݞ� p'���9T��S����� �Qb� o�of?�>rg;��G澍����   ����x��v�e�:e�e/\܊�� u
 �XV�+�UE��gRg �(1�������������12�i���t�   `��E\���:c��e/�a� G!���="�b��� 0J��-�*7p�Mw���4�:3�6|p   8YW�����ΘEY�ol�ށq; �F��Q?�x�f� p|��M�\�'+�SwP�֍P���2?����   ��y��N�eꌱV�U�pѸ �R�5R'ܖ�̞Z_�X� � �~���𵑻�j�qvm.u0���   8i���.ތ��R���aQ��o�~ϸ �T^��{DŠ�S�+ `T�����O�@��]��F��� �ԙU�   N^oP�K����q?R�a�_܊no�: �NV��{DY>�� F��; �)�ܹ;Yqnc!u0�y�˳�3   �	��īWwRg��ޠ�o\�}�v 8Yu��eU�#q���[��1��Wq 8&��Y�,>���z[[��N���x�]�K�    L�;�ƍ��������oFP�N��V�+�U1�_o\�[ �0p���h�埈�z�t��9�6�:� Ks���n��    &ԥ��ڵ����w0�.nŠ(S� ���j6p�(#���T�
 � UT?���zk���8�:�g\q   ��ՍW��DU�.��k;��ś14n����oW�?�� FA����q��M�@�ݳfl
��3+s�gY�   `���9��/o�BUE\�����  8Y5�W���#*�`���8 ��~���죩;��,sM8Y�fK3�3   �	��׋��r��=e/]ڊ�7�S� ���j8p�r����?~ u �Vï� p�v���������tL���3�	sj��   Ho�ۏ��v#�{��)#�7(��ߌ��~� �Ly�qUU���x5�* G�*㏧n��κ�$��8���   ���2���MW��bk��x�f�S `r��{DTÁ�; ��_��(eُ�N����<��Sg (˲X_r�   Uq��^�ti;��J��LUE�vm7^��âL� ����j�é  �z~���C����t�y�:�P�WfS'    ���^/����q}� uʉ������o�խn�  "��ܣ*[��׈0�j�U �ƙφ��}    IDAT����I�A}m��$�2?�V#u   ���2^��/���A�:��UUĥ����nD�7L� |[M���F��� ����hE$u��l䱶8�:�p�ˮ�   �i{��������(�*uα���k�݈7n�E5�������#������ �R3u  �T���d�8s���#��C`<�^��W.o��    xGUqe��wbmq:�g�����jX���qs��: xOyD��#n[�c} L4w &ZVV?\׷������(X�i�T�}��   FWQVq��~\�����T�-�D�Y���2.�܏k�]���,��_���R' @J�{b  G�ןiEߟ:�zj5�X[�J���(   PEYŕ�n|��k�ҥ�����b(��ڵ���W���-�v �����r�z�3O�O� �����Z�.�e����td����hX_��W���    8��������^/Z�<��:�8ۉ٩V괷������Al������SQt0"^J� )�0����g�ܩ�ג�ѱ2߉f#�aQ�N   �m���+[ݸ�ՍV#���v�ϴcn����_]��ck�7vb0�� H�*?_N� )�0��*>���zʲ�����ёeY�.Lť��S    �ʠ(���A\�9����v3f:͘�j�t�S�F��Ѿ]�7(b�7��n?v��1pD  �G���]6 L,w &V���(KB3�h7�3 �f}q��   ;�a���GD��yL���j��n6��̣�g�l��Y�o��,�*"�����"�����������^��n�x �H���G"�,"�rz &��; ��ןie7��Π���S' |����Ȳ��#N   `��e��� @-���]Y,m^���K�Ƌ�S ��  �����J�A=�.��0z��<g;�3      8U��J] )�0���x��e@
�0o�      ��,�����(�X� H����TUa��Y[4F�ʼ7L      |KUU��NU�6 0���TK@=-���kq����      �AUUN�  )X> 0y.|���Π���:� ޓ�O     ��r����M� '�����W�����O����T+u�{Z��N�      0"��w�*#�|4u �4w &N��WxqG\E�`ua*u      G�����8� L���>���z2p�`v��V#u      G �
 &��; ���]p�,����:�;     @TUꂻW���N ��f����]p��eY�⌁;PKs�      c0p�x衟��_V0Q��(k�����������L'�<K�p(K�8     0ܫack&>�: N��; %��+en��L;u���M�����     0��`�1��h� 8I L���p��i~����     &�8\p���[ &��; ���>�:�z��j�N �-K���	      ����=�����b��D���`��in����E�    �I6&��#"���R' �I2p`�dY|_��g�ӌf÷M@�,ι�     L���WUqj�S�7�� N�� c������8������r���v�ӝf�     �$���dI�����{j�@��,���n��
_Co}����+_����޵7��>��Z�@�#Hb P�5�|��>/(ɢMR@!3��/�'��!��"DdU�?ߓs*�0?�o�+� lw 6Ƶk�\o�J���W:�J^��     ��j�G��t��� �,� l����;Wr뺁(������/     `C�\�`���w���a����ڊ��n`=ݼ�S:�Jn]�-�      PFm�G� �� l����q%7܁5u��     �fʕ�sJ[� �������63W���;�~d�Ӎ��     �)��s�s�Q��/\g`#X: ��ۿ�����t��ƞ���v��n�     ���{i��^�{ `#��^9��D��O���v��gr��^�     ��l����?/�  �`��F��iV���t��E ��yw     `�
�]��c� Xw 6B��ߔn`=����[�}Q     �@�/]0wMJ?-�  �`���h~R���tso�t�3�q͟c     ����{���� �� l�l�Ε\3p�ܵ����jJg      ,ON�KW�]��K7 �2��ܹ��?.��w     `��
���ѷ����^� X4�- ���؉�+��z������n^�-�      �<�ҁ{�M���t ,�� �{����ADX��Ԛ&b����M�    �M������oJ7 ��Yl����.`=��l�N ��.�     $�z�� ������-w�doǏJ@\p     6J��s�Z� �j��5���+����P��     ��)�NX�&7?*�  �f��hܹ�����	 sq}ןg     ����{?,�  �f�@�r��t��w�M�Į?�     �M���G��N �E�p �~M��t�iJ �ϵ=W�    ��SD������o�ӿ�Z: ������_�����F��Ӗ�;P�k�;�      .�|�=""rL��?*] �d�@�vg���\�֖�;P�k�.�      u�n���P5w �����n`}�����     ��_p�H9��t ,��; Uk"}�t�����ގ�;     �6`�)�B P5w ��#\p�ʶ��T����;     P����	�4����mP�&·�y.������     �r��s��-�  �d� @�w�l�1p�k�     �.����]�)�  �d� @岁;W�#�N ��mw     �r9��=""r~������ �E�p �^���VD�Q:����ہ���     T/u��$mN?v��jY8 P�W��oF�o,se�����_�     ����G��~P� ���z���N`�ٷ���jJ'      ,L�7gྵ�|�t ,��; ��N��K7��rX�u���+      P����޿Q� ź�z����g���;P�]w     �V9G�t��䰉 �Z� T+G|�t�ͼ���VS:     `!�]o��h"�D P-w ����2��w�6[��;     P����� �2p�^�1p癤l�Tƾ     ���]p���� �(� ԫ��<��7p��;     P��o��=7��� �(� T+G��L�>�N ����     �UjK,U��7~�_���� �� T*7MxϦ7p*�e�     �(����,��� �E0p�Jo���x%"�Jw�޺�qo� �۲p     *���tByk��� �� T�O�[�X]�K' �U�     @}rjK'��$w �d�@�R�^:����.�ui��    �m��H���	 �� T)5�j��_�܁�d�      *���S��J7 �"�P��I�<��#�d
�#Y�     ��9"m��&�R: ���:�������}���1p     j����?�]p�J� T��-e�df�T$y*     P��o��=7� T���*��w�c�����T:     `���tA19��� �� �)��;s1u��Hk�     T&���	�dw �d�@�\pgN\pj�u�     @Er�ț��n��; U2p�NM~�tup��E�9�d�     �#�]�Ҟ��?���# `���Sܙ���;P�I�GΥ+      �'��tBq����� 0o� T��N~�tu�u�u��|a     �K�f���ى�J7 ���P�q�x�t��6��v@%��H     ���h������P��ԿX��z��>Rʥ3 ��x�^     �9u��s�m$ ���; �I��~yc�\qj0���     �H�ODDΎ Pw ����F��b��`4�&/     P���J'���F���P������\�����N�    �z����s�� 0o� T'�-��b�&.�kn2��R�     ���)"��+V��� `���N�p����k�b4-�      07�s��O�H6 T����lm���O܁�v>4p     �{�?I9�H Pw ��s�b��b�����7y    �z�-��J^(  �f�@��Nf��>Ŵ�Kg \��;     P��#����4.�P!w ꓳ���p�`='mt}*�     0��Qn��K7 ���P��㷘��؛$�z:NK'      �M�=�������; ���7�n85p���ț�     @=ܿ�i�f� �7w ���s���`�M`=�\�K'      �I����%���_�P/l �����N\p��p��x�M^     ���""��X5�kp����P#w��R̺�t�S9v�     �H�=y�����K7 �<�P#�Lf!cW܁�r|n�     �#w��	+��M�J7 �<�P�����ۥ;����5 `}���l�M^     �9G�}���.�Pw �2�u������X#'�H9��      ����"�g_�I[� T�������~ica�G.!���b\:     `nr��گ���	 0O� T�iw�Y�񴋮O�3 ��ѹ�;     P�ܷ�V�V�Pw ���7K7P���t�_ur1�Yۗ�      ���"���W�� �����4͖�,���c�շ:(�      07��9��I�7p�*� T�I��,���w`�����|\:     `nr�sگ��� ���; ��7JP��7N��vp6��O�3      �&�>��:M�� `���J�f�tu�̺���� _��ɠt     ����Ed��~��V���P�&ǵ���l0)� �m��     T$w��	+/7�����P�&�_�X��Co� �i�t9��      ����J'��&�� U1p�*9����¹���ώ/K'      �Q����+/���Pw ��le���p�qm�Jg |���(�Ӯt     ��䮍���5Mv����P���_�X
W܁Us���v     �.���NXM�N �y2p�*M4�,���t��'m<���     �.�����
O��*� T%��,�!)�J�\�N      ���G��t�zHa+@U����,��x]�Jg Dۥxt:,�     0W���'�� ���; UI�[,G�'�P����2RΥ3      �*w��	k��.�Pw ��;�t|1.� l��r�;�,�     0_9E�m銵��q���P�&�N`s��}v<�Yۗ�      ��ϯ�{���y�t ̓�; U��k�3k��] ��9ǝ���      s����'�4[M� �'#@ ���kK�;Pʽ�˘��     T'G�f�#֌� u��@Ur�嵍�2pJH)ǝ���      s��6"R�uc+@U��P��[�,��`}ʥ3�s��2f��     �ݤt���ۥ `�� ���6�*�W܁%J)��C��    �:�nZ:a�8@e��P��k�wx6*� l��    �Z徍�>yZM�4� `�� �J�^�X���q�Kg ��R�yt^:     `!\o�"[	 *���l��n�|]���rR:� ��Ϣ�S�     ��0p��&�J P/l T%ǖ�6�8x<*� Tn8i���e�     ���)"��+�T�]�  ����d�)����X�>{9��      X�۟A�4� `�� �K㵍2�.���tP���Q�\�Kg      ,Lj}�ze9�J P/l �%�V2�����_�9>|pV:     `qr��g�+�V�[v� T� ���p��2FӶt     ���n�t �"� �d��q|1.�Td������      �Z�� ���; ��K' y��it}*�     �89E��� �
1p ��óQ�ɣ�gwx6�óQ�     ����t �b� �(��]q�M�r���t     �¥�� �"w �9{xj�<�>;�iۗ�      X��"�Y�
 `�� ����I�g]�`M=L���t     �¥v\: XA�  p��w�饔�ݻ��3      �"w��	 �
2p X��\_�����M��      ����~V� XA�  0�vq|�qz��;L���E�     ��Hݤt ��� 䳣��	���S���GΥK      �#�� ��3p X��qLf}�`�w�$&��t     �r�>"��+ �e� � 9G<8q��z�N��:,�     �4�s� �j�  ���t�¦m��?-�     �T�5p ���; ���>�F�3�����h�T:     `ir�"R[: Xa�  v��t������K�I     ���z; ��� ,��`��i�`�<L��ó�      K��q� `�� ,�+���̺>~��q�\�     `�r7��}� `�� ,���(FӮt�~��Q�Zo�     ���v �I� ,A��\q�����q6���      X��#w>' �:w �%yx2��K�3�B���q��]     �͔�ID�� ��� ��O9�]�� 
M�x��q�     �bR;.�  �	w �%�wt)����)��?9��w�     �P���g�+ �5a� �Dm��+�Q޽{�co�     ���v �i� ,ٝ���]q��p��Y<z<,�     PT6p ���; ���]��G�3�;<ŧ��Kg      ��YD�Kg  k�� ��;��C�.G�x��q�     ��r;)�  �w ��.ŽCWܡFӶ��||�K,      �#w� ��1p (���Et}*��QJ9~��QL[��     ��4"�L x:�  ��}�{���3�9z��q���3      VBjǥ �5d� P��Ë�u.=C޿�g��      �!���a  ��� ��)n?<+�<�O�����'2      ���� �U� ��d�I[:��ǃ�x�U      �R�y�- p5�  ������������'�3      VJ��/� �)w �pz9����ur1��۟EΥK      VKn}�	 \��; �������	�N�x��A�ɺ     �r��MJW  k�� `E�m�?�,���Yo�>��K�S      VN��J'  k�� `�|��,f]_:�
Ӷ���QLf]�     ��#��� ��3p X!m��g�3�/1����G1��     |��M#��^ ��1p X1Oqz9)����K��b8iK�      ��4s� xv�  +�{��s.�DD�r�u� c�v     �����~Z� ���; �
M۸spQ:6^���b4+�     ��R�z; 0�  +���M�������׷�l��     ��ˑ�Q� ��  +*���;)��O9��ȸ     �I�v�S� ��  +��r�Jg�F����� Ά��      O"�� ̑�; �����M����>�[��ܸ     ����E��� @E� V\�r���q��ެ���?<0n     x
y�z; 0_�  k�l8�;�3�Z���_t�c�E      �XΑ�I�
 �2�  k��g1���3�:�Y��� c     <��M"r*� T�� `M����O�#�\:�1����hj�     ��lX: ���; �����ó�P���4~����̺�)      k'w���s `�� �̝��8:�΀�vz9��nF�{d&     �U�� ,��; ���ݓ�:W��to�>�θ     �Jr�"�i(oZ{    IDAT� �R�  k��S���q�K��Z�t��=�      \]�y�4 �8�  k�|8���΀�q��Y��Ը     �Y�����  *f� ���^����ur��Ν����y�     ����qD�� @�vJ  �l�p�$n�؋���h���K�ۏ�l8-�     P�y�  �X.� ����|����$�_M�x�G��      s��iD�Kg  �3p ��p���?=.�+��ro���i[:     �i6,�  l w �J�\������3���'�����h=�      `nr�F$ǅ ���)  ���?��[7�⻯�*�E|��q�9�(�     P��z; �$�  �y��Iܼ�/?�t
,M�r���Q��K�      �'���i�
 `Cl�  `�r���'G1�x< �a8i����     ,HjG�Kg  �� �Bm����d֗N��:�Ǜ<���:      "�ȭCC ��� Tj����b��S�;�ۏ��S�     �j�v�} ,��; @�F�6~s�0��q�ԣO9~��Q|��qd��     X�i6, lw ��]�f�#[S�ᤍ7?؏óQ�     ���v�=1 X.w ���r���t<���a����1��S      6B�9: ,��; ��8:�;w�Kg�SK)���;w��O�D      ���D$�� ���)  ���#���G��N�'2����O�\m     X�4�N  6��  ���(~��a��6����0����q;     ���n�z; P��; �::��>92rg%�)����w���S�     ���f��	 �3p �PG�����G���;��b4�_��O�i
     PB�ۈ~V: �`�  ��b���0z#wV�������c4��K     �R�lX: �p�  ��ro~��Y_:�5�����g�}�     �����ݤt ��� ����7?؏���l���l�|�a���S      6^��� �g� @DDL�>���Gqz�"��v)޹s���(�>��      ��� +�� �?k�o�>�ǃ�)T��b�����?u     `U��0"r� ��)  �j�9��{'1m���Q:���]�>;5l     X59Enǥ+  "�� �����Y\�����;��ó9�ǻw?��      ���v `�X* ����o�?��-�j���9���>4n     XE9E��� �w  ��h��/�ۏ�'��)����a��w���t
      _!�F�Jg  ��N�   V_�9�p�$Ά����MӔNb���]�w�$N/'�S      �:9E��JW  |��;  O��� ��6~��W�ƞ%���s|��">}t)��9      �i6���Uc� �S9N�_�}?}����ϗ�aE���N��)      <��"�ƥ+  �?�  <�>����8���������]:�B�m���ÓA�      ���� ��2p ��N.���>����[/?W:�%J)ǽ�����yt�7>     �JN�g��  _�� �g��)޾s����w_�ݝ��I,���Q|��qLf]�      � M�Kg  |)w  �b�t�����_���|�`0n��'q6��N     �R���  �J�  �Mۧ����?��}��x��^�$�`�����Y<<Dv�     `���0\o V��;  sw1�ś���܊�}����jJ'q]���G�q��2��MN     ���z; �� X��#��|�����/?W:�'�R�{Gq��E�}*�     ���� \o V��;  5k�x��q�98��~��x�ś�������YL۾t
      s�S����  ��� X�����~r�x�Z����篗N�r����(>�?�Ѵ-�     ���0\o ց�;  Ku>�Ư?:�o]��y�x�ֵ�I+�O�.�     T.�.r�z; �� (�l0�_}�(^y�F��/��D)�|w.bf�     P=���ub� @Q'�8���7��{�=o��\4MS:�J���ώq��"�.��     `	>��>.� ��� X	��Y�{�$n���^}>���󱻳U:�
�q��.b�d)��     �I�tP: �� �Rfm�ŝ����K��w^�/޺V:k-�����E�^NJ�      P@�g�;� ��� ��ԧO��d��v�[/݌��|���#�יu}<<�gǗ1�v�s      ((�� �!�   V�d�ŝ���{x/޺�y�V������jJ�����q<8���q�\�     ��r7��g�3  ���;  k#�Ǘ�x|9���������x3^}�F\��.��t��Y<z<���aL۾t      +#�� �-w  �R�9N.�qr1���[7v��n�k߸/޺V�nq��6����a'm�      VP��#RW: �J� ��`��`�Ɲ����ݎ�n]���/ݺ���+��L·�8�����0c�v      �FΑf��  Wf� @ufm�Gq�x�[M��ܵ?�޿��^�lo��j�����q�\L��rm�J'     �&�l���  Wf� @������$_N"�<""�v�����x��nܺ��]߉[��bwg��������4����p�J;      W�S�٨t �31p `#��>N�>N/'_��ww��k����{��qmg;���_��?��lE�4O��ק�I�i�Y�I�i��Y�)��      *M��� �z3p ���v)κ��g��&���h�>��?�눈�s�)Gץ�R�l�     �"�>r;.] ��� ��RΑ�ї.     `ӥ�eD�� ����         \]���ݤt �\�        ��ϯ� ���        `M�n��Jg  ̍�;        ��J�A� ��2p        XC�G��t �\�        ���z; P%w        �5��Èܗ�  �;w        �u�S�٨t �B�        ��4DD*� ��         k"�.r;.� �0�         k"O�Kg  ,��;        ���,r7)� �P�         k M.K'  ,��;        ����8"��3  ��        `��H�A� ��0p        Xai6��}� ��0p        XU9E�KW  ,��;        ��J�AD��  Kc�        ��r�"���  Ke�        ���t�t �R�        ����"w��  Kg�        �b��t @�         +$���Ԗ�  (��        `e�HS����e�        �"�l���  ��        ���"O��+  �2p        Xi:��T: �(w        ��r�"���  ��        ����ȥ3  �3p        ((���ݤt �J0p        ((M.K'  �w        �Br;�Hm� ��a� ��a�β9� 
����$�2�}POR�' �*�l��{      (�ї��  �"p        (��KD��  �"p        x���k�
 ���        <Y_^"�W�  8�;        �e�#�k� �C�        <Q�}���� pHw        �'ɶF��z �a	�        ��� �_�        <An׈�U�  84�;        ��e��z ��	�        �/�٪g  ��        ���G���  � p        x���DD�� p
w        �ɾGn��  �!p        x�~�Y= �4�         �m�hK� �S�        <��{;  !p        ��ܮ}�� p:w        �����K� �S�        �Q_/٪g  ���        �^�G.��+  NK�        p'}y��^= ��         ��[�v�^ pjw        �;�˷���  �&p        ��l[�~�� pzw        �/z{o ��         _��-���3  � p        �����T�  ��        ��r�F��z �0�         ��}�� pOw        �O��kD��  C�        |T���R� `8w        ��˷��� pow        �ȾGn��  C�        |@�}��  0,�;        �;�F��z ���         ����  �$p        x��n}�� 04�;        ���v �'�        �A_/٪g  O�        �;���k�
 �)�        ~���٫g  LA�        �+�#�K�
 �i�        ~�//� �Y�         ?�}�ܮ�3  �"p        ��\^""�g  LE�        �ٶ��V= `:w        ���˷�	  S�        �K�KD[�g  LI�        �/}y��  0-�;        �_r�F��z ���         ��� �	�        "����l�3  �&p        Ȍ\_�W  LO�        L���٫g  LO�        �-{�z�^ @�       ����%"�� ��        �V�=r�V�  �/w        `Z��DDV�  �/w        `Jٶ��V= ��        S��K�  �C�        L'�і�  ���        ���v �c�        S�}�hk�  ~B�        L�{; �q	�       �i�~��[�  ~A�        L�{; ��	�       �)�v��{�  ~C�        L �� ���        ^�׈l�3  ��;        0����V�  ��        ���z�� pw        `\���� NC�        ���٫g  �Nw        `L�#�K�
  >@�        ���� �L�        �x�G���  |��        N_^�{; ���       ����yo 8#�;        0���DDV�  ��        �0��ۭz  �$p        ����v �3�        CȾG��� �L�        �߾UO  ���        ��e�"�R= �/�        ����  #�        ���޾V�  ��        ��yo ��        8-��  c�        �� `,w        ��r_�� F�        �R__�'  pgw        �t�� �I�        ���v �1	�       �S�� 0.�;        p*�� �%p        N#��{; ���        �i��{; ���        �)�D��z  $p        N����  x0�;        px��m�� ��	�       ����K�  �@�        Z6��  ��        ����  ��        ��m�� 0�;        pX�� �"p        ��}�� �	�       �C�� 0�;        p8�� �$p        '���	  �        ��m��o�3  ( p        �{; ���        �ad߽� LL�        ��v ��	�       �c�-r�� 03�;        p}}���� @!�;        P/{�v�^ @1�;        P�{;  w        �Z���{;  w        �X_/ѫg  p w        �Nf�v�^ �A�       �2}�D��v  ��       �"�zo �w        �Dn��l�3  8�;        P����  8�;        �t��"�^= ���        O� ���        O��ѷ�  ��        x���TO  ��        ��d�"�Z= ���        O��k�  L�        <Go���z  &p        ��{o ��        ��e�ܮ�+  88�;        �p}�DDV�  ���        �ceFn��  ���        x��]"�W�  ��        �e�� ���        ��-"[�  NB�        <L�� ��       ���}��[�  ND�        <D__�'  p2w        ���m�� ���       ����R= ��        ��=r�V�  ���        �]��Y= ��        w��� �4�;        p7��"�U�  ��        ����R= ��        w��ѷ�  ���        ���  |��        ���{D[�g  prw        ��r}��  � �        ��d��n�+  ��        ���^""�g  0 �;        ��]�G  0�;        �i�-٪g  0�;        �i}}��  �@�        ��d�"�V= ���       �O��R= ���       ����ߪW  0�;        �a}�DDV�  `0w        ��2r�V�  `@w        �Cr["�U�  `@w        �C��Z= �A	�       �w˶E��z  ��        ��z  �        �=r�U�  ``w        �]�v���� ���        ���z��  ���        ��Dd�� ���        �u��  <��        ���"�R� �	�       ���۵z  ��        ���ۥz  ��        �����z  ��        �Խ� �Dw        ৲�m�� �D�        �O�� ���        ?ʌ�n�+  ���        �A��3  ���        �A_/�  ���        �N�-�o�3  ���        �Nn��	  LJ�        �#3r�U�  `Rw        �o��"�W�  `Rw        �o}�VO  `bw         ""��m�� ���        @DD��v  �	�       ��H�;  ��        @�Dd�� ���        @t��  ��        f�[D[�W  ��        f� ���       ��R� �A�       `b��٪g  @D�       `j�]�'  ���        0���R�  �&p       �I�v����  �       ���v��   ��       ����}��  ��       ��r�UO  ��       `B�]�'  ��        0��׈l�3  �w        ���v  �J�        3Ɍܗ�  �Sw        �H��3  ��        0��]�'  �/	�       `�E��z  ���        &��[�  �-�;        L"�k�  �-�;        L ����  �[w        ���v  �@�        �}��   $p      ��*h    IDAT ���Fd��  $p       ���~��   �"p       ���� ���       ��r_#�W�  �w�       ��r�� �y�       `T���R�  �M�        �z��{�  x7�;        *�[�  ��;        �(�w  8�;        ��=�g  ���       `@}�UO  ��       �h�G��z  |��        ��Y=  >L�        ��۵z  |��        F�=�m�+  �S�        0�ܗ���  �)w        �[�  �$p       �Qd
� 85�;        �-n��  �iw        D��	  �%w        BF�k�  ��;         �%"z�  ��;        �-p �s�       ��� �!�       ��r�"�W�  �/�       ���~��   w!p       ���}��   w!p       �˶Fd��  w!p       ��� �H�        pbw  F"p       ���-���+  �n�        pR}�UO  ���       �I�VO  ���       �eF4�;  c�       �	e[""�g  �]	�       ��r_�'  ��	�       ��r_�'  ��	�       �d�m٪g  ��	�       �dr_�'  �C�       �d�  �J�        g�=�o�+  �!�        p"�� ��        ND� ���        p���#  �a�        p�����3  �a�        p�/�  ��        p���	  �Pw        8�̈�U�  ���       �	���g�  x(�;        �@�K�  x8�;        ��ۃ;  �M�        G�=���+  ���        pp�/�  �)�        pp���  �)�        pp�<� 0�;        X�-"{�  x
�;        X��z  <��        ,w�;  ��       �ae�w  &"p       ��ʶGDV�  ���       �A��v  &#p       ��j[�  x*�;        �w  f#p       �ʶEd��  O%p       �#j[�  x:�;        P��z  <��        (=� 0!�;        L�="[�  x:�;        ��v  &%p       ��ɶVO  �w        8���  �I�        G�="[�
  (!p       ��� ���        p ��  �K�        �m��   e�        p���  PF�        �m����  e�        pm�^   ��        p��  �M�        �� ���        � 3���+  ���         ��v  �       �d� ��        �@�  w        8�   p       �z�#�U�  �rw        (�  ��       ���  ��       �Z߫  �!�       ��w  x#p       �J�#�U�  �C�       @��{�  8�;        Tjw  �?�;        ��  ��       @!�;  �C�        ���  �O�        Uz��^�  C�        E�{o ��       @�;  |O�        U��  �M�        E<� ���   ���;�m]ɡ(Z�|���_���C'�-�,i-���`�     PbC�  _�       ��v�cl�g  @+w        ��a�  ��       @��.p ���        P��Q}  �#p       �� �'�;        T�,� �ww        ȶ�?  ���        �mw��  ���        �	� �!�;        $���T�   -	�        �w  xH�        ɶM�  ��        ����  �%�;        d��  �A�        ���G�	  Ж�        2	� �)�;        $���T�   m	�        �f�  ��       @��~�>  ��       @�M�  ��        ��Q}  �%p       �4�w  xA�        I���v  xE�        Y�� �Kw        �r� �+w        H�m�'  @kw        ȲYp �W�        ��.p �W�        �d�>�O  ���        ��.p �W�        �e�W_   �	�        �vcl�W  @kw        H�Yo �]w        � p �]w        � p �]w        Ȱm�  @{w        H�Yp �]w        � p �]w        � p �]w        Ȱm�  @{w        H�Yp �]w        �`�  v	�        �w  �%p       �� `��        2lw  �#p       ��mÂ;  ��       �Ѭ� �[�        p4�;  �E�        ۆ�  �!p       ��Yp ���       �pw  x��        ��o ���       �p
w  x��        'p �w�       �h��  �!p          ��;           -�       �h�V}  LA�          @w           Z�       ����U�   S�          Ђ�          ��           � p          ��;           -�          hA�          @w        8X��>  � p          ��;           -�          hA�        G���   � p          ��;           -�          hA�          @w           Z�          Ђ�          ��        p��>   � p       ���� �-w           Z�       ��L� �;�        p8�;  �C�          @w        8�w  x��        �p �w�          hA�          @w        8ZD�  0�;           -�          hA�        ��'  ��        p�� �;�           � p          ��;        .�  �)�       �h�v  x��        �p �w�        �T  ��5       @#�  �K�        )�  �G�          @w        �� `��        R� `��        2Xp �]w           Z�       @
�  �G�        	"�  �G�          @w        �`�  v	�        ��  ��          hA�        B�  {��          hA�        "�/  ���        � ��  ��        �w  �%p       �w  �%p       �w  �#p       �� `��        R� `��        2Xp �]w        H� `��        2Xp �]w        H!p �=w        �`�  v	�        ��  ^�       @+�  ��        �� ��;        d	�  ���        Y;  �"p       �4w  xE�        I;  �$p       �,w  xI�        i�  ���        ��\  ^�c       �,a�  ^�       @���  /�1       @�  ���        ���  ^�       @�;  �$p       �4w  xE�        Y,� �Kw        H!� �W��        �w  xE�        Y"��  ��       @�� �3w        H%p �g�        �)$;  ���2        d� �S~�        �("�O  ���        �ɂ;  <�        �,� �Sw        �d�  ��[       �D!p ����        UT   m	�        �w  x�o        2�w  xF�        ��  ��        EHv  ��e        �d�  ��       @���  ��       @���  �#~�        �M�  �)       @���  �%�;        $�  �2        d� �C~�        �M�  �)       @���  �%�;        $�  �2        d� �C~�        �M�  �)       @���  �%�;        $�  �2        d�e�a�  ��       @�� �ww        ��  ��/        *� ��d        (w  ��/        *� ��d        � p ���       �@� ��d        � p ���       ��"� ����       ��w  ��/        
��  ~�K       �
��1��
  hE�        U�� �~�        PE�  _�!       @�;  |�        EB�  _�!       @�E�  ��        �Xp �/��       �H� �?d        �"p �/��       ���  ��C       �"���'  @+w        �Q}  �"p       �21FXq ���        P)$<  ��1        T� ����       �P,k�	  І�        *Yp ��       @�� ����       ��"� ����       �R��  @w        (!� ����       ��"� ����       �T�a�  �w        �k�  Ђ�        �Yp �1��        ��"� �1�        P/��  ��;        �E�  c�       �^�x  `�;        �� �C�        �bY�O  ��        P-�1FT_  ��        Ёw  �       @!�  �b        h ;  �       ��E�  w        h B�  ~�        Ёw  �       @� @�        �w  �       @��1��
  (%p       �.B� ���       @�Z}  ��       @!p ���        �E� �6�;        4a� ���       @� �8�;        t��y  �6?b        h"�  \��        ڈ1B� �u	�       �+�  \��        	�  \��        :�� ��	�       ��� paw        �$$=  \��0        tb� ��       @#w  �K�        �D��  ��O        ��� �E	�       ��Xn�'  @	�;        t�Xp ���        �L� �(�;        tw  �I�        �Xp ��        �Ͳ�1��
  H'p       ��B� ���       @G˭�  H'p       ��bY�O  �tw        �H� �	�       �!�  \��        :
�;  �#p       ��b�U�   ��        �Q�!� �Z��       ��X�/  �Tw        h*�[�	  �J�        ]-� ��;        4e� ���       @W� ��;        4w  .F�        ]���  �"�~       ���� �u�       ��Xn�'  @�;        t�Xp �:�        Иw  �D�        �Yp �B�        Иw  �D�        �E�2  ���        ��� �E�       ��X��   ��        ��� �E�       �9�  \��        ��� �E�       �����>  'p       ��b�e�>  'p       �	�r�>  'p       �Xp ��        0�  \��        f p ��        0�X��  �pw        �A,�  N̏        f�ܪ/  �C	�       `!p ���        0�e��   %p       �IXp ���        0	�;  g'p       �Y,��  pf~�        0�e��   #p       ���z�>  #p       ��,w  �K�        	�;  '&p       ��� 83�;        �dY�� ����       ��,k�  p�;        L&�[�	  p�;        �f� pNw        �L,�O  �C�       `2���'  �!�        0�e�  ��/        f�ު/  �_'p       �	�"p �|�        0�e��   ~��        &��  ��	�       `B�ܪO  �_'p       ��2F��W  ���       ���� p2w        �T��O  �_%p       �I�w  NF�        �Z�  ���        &�:ƈ�3  ���       `Z1�b� ���       ��b� pw        ��w  ND�        ��O�	  �k�        0�X-� pw        �Y,�  N��        f����   ~��        &�� �s�       ��b�U�   �B�        �[�  ���        &���. `~~�        pV� 8�;        ���;  �M�        '��  ��&p       �3�� �	�       �b��1��  ���       �;  ��    ����Ǯ��������)�EY6eS�eE�D�X��4
6.p�"�Vۥ��v*��VR��O��-�,���z-k%Q�1��P$[�g�9�{^�V?�H�{9��\   ��w  X.�;        4"��z  <�;        ��w  N�        �p� ���      ��Ml    IDAT @+2#:W� X.�;        4�w  �L�        -�]p `��        А�]p `��        А��  ,��        Z�!r `��        И��	  p*w        hL�� �B	�       �5�� �e�       @c�""�g  ��	�       �9��#  ���        Р���	  pbw        h�� �%�       @���z  ���        ��Y=  ND�        Mʈ~�  '"p       �Fe7TO  ��       @���TO  ��       @���'  ���       �U]�}�
  86�;        4�w  �D�        -� � w        hXvw  �C�        K� X�;        �,3�w  B�        ��~��   �"p       ��e���   �"p       ���c�  8�;        4.�!�B  ,�W�        ��P�   �J�        +���z  <��        V ��z  <��        V@� ��       `���D�  ̛�        V�w  �N�        +!p `��        �w  fN�        +����!  �˫U        X��7�  ��        �&�X�   K�        +�;  s&p       ��~����  �$p       �UɈ~�  �$p       ��I�;  3%p       ���~S=  I�        +�;  s%p       ���.�� 0?w        X!W� �#�;        �P���	  �w        X��  ̏�        �(���W  �7�       `�\q `n�        �R�� ��;        ��� ���       �Zu}D��+  �kw        X1W� ��;        �X�c�  ���        �lp� ���       ��e7Dd_=  "B�        ���X=  "B�        ��öz  D��        p� ���       ��e7Dd_=  �        @D���	   p        "r� PO�        �� �,�       ����Ⱦz  +'p        """W� �%p        """{�;  ��        @D� �'p        ����W�  `��        ��r�VO  `��        �ײ�TO  `��        ��r� PG�        �^v�X� ���        ���;  U�        �7d���  �J	�       �o�a���� �
	�       �oɈ~� �
	�       ���a[= ��        ߑ��z  +$p        �#�1"�E  \,�@       �Gr� ��&p        )�m�  VF�        <��  \4�;        �h]�}�
  VD�        <V��	  ���        x,�;  I�        <V�����  ���        x�̈~S� ���        O��� ��!p        �(�m�  VB�        <QvCD��3  X�;        �T�� p�        �S尩�  �
�       ���~Y= ��	�       ��ˌ���  4N�        K��	  4N�        K���	  4N�        K�cD��3  h��        8�\q ���       �c�a[= ��	�       �c�~Y= �F	�       ��ˌ�7�+  h��        8��  ��;        p"ݰW= �F	�       �����n�^ @��        ��尭�  @��        ��	� 8w        �Ĳ#R~ ���
����       �!#�M�@+@c� 4%#��       k�öz)p�)w �2M�m       E�s��J �6 ڒ�m       &��~S�V�w �"�1�g      �r��i% h� m�:�6      �$p�Z��1l 4eJ�      .RvCD7Vπ��t� �Ń��t�m       �w(��� �,� h��Wo       X�;ԙb��)l ���n      \��ǈt��h% h� mI�6      �
��C� h� ��l      (��^�X��.�7 �YД�&�6      �9�!G�Z	 ��@S��<�       Jd䰩듓� 4E@[�i��       �V9�UO���B+@S� �%c[=      `�����4\�̱z �%�; ��      T�.��T�����x�CW�h������      �BݸW=V�ͧ��; ��      �Pۈ���*w�P/@3� ��w      �J�E�c�
X�m�� �w Z��       źa�z�ʃ]�K@3� 4dʈp       �X�Z[�HC�q��f�h�[��cDd�      ���.����E9�����f�hƯ���7k       3����E針�p 4C�@3��]�      ��nث� ��;4 4C�@3�m'�F      ��������
]i& h���f���       s��+�p:� �Ќ�G.�      �I~�a�e�w ��1�Wo       ���"��z��A�  8+w ���]��       �7�W=��;�; ��Ў�	�      f��p�v�� �w ڱs�      `v�>��W@�v]�; ��Ў��       3��+�p�r7	�h���f�ެ      �P7��\e�WO ��"p�.�      �S�G���ЬGh������      `�\q�s�[�h���v��      0[9
�Ἰ�@K� �ç�      �+��~S��4E�Wo ��"p��L�      f�\q��0M��� 4C�@;��      �X�{��3�Ew �!p�%w      �9�.��T���dN�� ��hF
�      f���'@�:�h�������       <Y{��3�)S�a� 8+w 2=W�       ��Ȍ��+�)��]��  gE�@K�       ��^�hKƥ��W# ��; -�R=       ���a��%8C��_��a� 8^%Є[��W���      �qd���;���W�Vo �� p�	��x�z       Ǘ�����=�V� ΂��&L)p      X��7�WπfS�� �	w �0��I      X���'@3�~�� �	w �0M�M      ���W=�1ew�z ��; M�B�      �4��X=���j' h���&tޤ      ,�+�p6�]\��  gA�@��w      �%����	І����; ��	�      �(��~[��o
� M�Ј��       ��+��즌�� �,�h��      `�r�~y�8�)���  g��B ����^�      ����a�z,ZNӵ� p� ��w      �E�Q��$��� �,�h��       K��&"���\S
�h���F��      �t9�WO�Ś2� 4A�����˥��       �	���2�͍�?<�� �J����_\q�      �]�o�W�bݿ�ߨ�  �J�����\��       ��p�No�$p`�� ,^�\p      hD{!k��麝����J���<r�      ����z,Үs$����x����      �!9TO�E�v;GX<�; ��w      ��d?Ftc�X�k� �Y	�h���       8[9�UO����X<�; ؽ\�       ��Ս���3`Yv�#� ,������	       ���"�m�
X��� �Y	�X�.nVO       ���xP=�e�]��  �J���M�;      @�r�Dd_=�w �O���]�����w       p>rܯ� ˑ�SV� �g!p`�r|p�z       ���I�7?��׫G ����l�N�      в����+`1v��[� �Y�X�)�       ��6���q=|8h) X4�; K�M      @�r�Fd_=!� ,����˗�       p�2rt��c7MZ
 M���yS      �
���%�x�z <�; K'p      X�����W��ej) X6�; ����To       �b�+��T��; �&p`��W/       �b䰍Ⱦz��4ݬ�  �B��b���݋��w       pqrsP=f-C���	�X��>��{��;       �8ݸ~TO��B���P= NK��b�}���       \��"�m�
�����U= NK��b�v��      `�r<�� �6<��Wo ����XSī�       �x9l"��z��ԇ�� ,����ʈW�7       P�s�kw �K��rM��      �J���'x�)oUO ���
���x�z       E2��܁��I��b	�X��w      ��ƃ�	0K��^��  �%p`��|��6"nT�       �P�G{�+`v2��� �� ,�?歈��       �JW�Ủ��Xw )��]�      �z9l"��z�Kƕ�����3 �4� ,�Qt�Uo       `��+��mG�� ,������	       ""r܋H)��.�� �4��`�2�v�       �"#GW��M�
 J��R��      �׺q?"�z�G���' �i�X���       ������+`6r�� ,���Ź��Gۈx�z       󒛃�	0��j� 8�; �����      ��d�����0SN�To ���8]���	       �T�;DDDF܌���O| �8w �{�z       ��^D��3`��n��j� 8)�; ����]�      ����q�z��Ç�~X� NJ����"]p      ౺�ADd�(�������89�7_       <^v��^�
(7��� pRw '#^��       ����z���� pRw �ֿ���)�Z�       �-�1��g@�I��	�X����7�7       ���R��5�nWO ����(�._��       �2��}�(�7�|�Ѷz ����eI�;       ��;+��c��U� ����(ݴ�      pl9�G�L���ؾQ� N�+7 e�\p      �2#ǃ�Pf�t��E��,w�'       �,�� �R�U�$p`Q�j`1��ٯ^����;       X��"ǽ�Pb��� pw #��Wo       `��ͥ���p�r��7 �I�X�.�7�7       �P]9���M߯^  '!p`9��S=      �����	p�2^����J� 8.�; �1E�Y�      ���n���3��僣7�7 �q	�X��V       `ٺ�+��Q?��z ���E�����U�       `�r�Dtc��P9�~R� �K��"|~���W�       `�\qg}��� p\w !NoVo       �9n#ҍ5�#c�S� �K��"Lw       �HFn�G���"o���; �8� ,BF��z       ��ƃ��O����A��z �Wh ,�.�      p�2#GW�Y�i�{�z ������+�^��      @[��ADd��(?�  �!p`���x�G���      @c����W������ �8� �^��f�       ��m.UO�1M��� �8� �^F��z       ����a�z����a� 8�; �7e�U�      �v�+���ҵ�W�U� ���0S�]=      �ve?F���p�2�}G�=�; �v烏��O�w       жn{X=���92��	�����oF�X�      ��}y�}S=�U��� ̞��Y�.��z       ���;����O�7 ������Wc      p1�߸�N���� �i� ���;       �۸�N�2�����+�; �I� �[
�      �89��N˦n�oW� �'�0[7�э��Y�      �u�6��'�9z��  �&p`��ީ�       ��䰍���p.��V� �D��lMS��0       %��+�4j��TO �'�0_]�]=      �u�a�w�4���� �$w �k7�S=      ���6��Ӟ��u���V� ���0Kw>�hoU�       `�r܋��p�r�?rt���0K?�y;"6�;       X7W�i�.�Wo ���0K�����       ��+�4'��w fK��,M9	�      �W�i��v� x�; �4E
�      ���"���gg�~�~�Y�`~��WcF��0       3��m�G���8��o�N� x�; �s�ߊ���       �W�iδ��� �Q� �Ov�VO       �o��6��G���M�;� �Q� �N�$p      `vr��;��Q� x�; 3$p      `�2rsP=�H�U�  E��������       �R7D���˜^������� �m^i0+/u�y3".U�       �Gʌ���6M�q;�[= �M����v�UO       �'�6�Wπg6u��z |�P=  ��.�_e�fo;�q�7����f�c3�1�]�]F�_�	:���h7��n���ރ�q��Q|�Ńxp�+�       ˖�mc��慎�3�I�������|/b����}W6q�`�����	��w1�}l#"�_��{���/��>��~q?&�      ��q/�ާ�Q�8�)�w�7 ��9��l���=�̏#���]f\���.�ǥ�1�^�<<��ǟ݋�|�E|q����"      @��w]qg鎆�ϟ�����g�C �+.�0}���n7��Wn����A\;��R���.�_ُ�W��ӻ�>����޹��      ���q����cZ,V��ßE��� _�0G��=_-�^_��/\ދ����p�?���w�?������c�;      ���0vw?���v���C�����������}/^=��W�#g�3�^�׿x��7���{�-       ���^D7F�TO���x�z �!�; 3�?�^�źvy/n=)�����H���x�ֵ��O�Ư�Y��I      �}y����3�Tr�ީ�  h&wRX���������;�{�!^�q9������������I|z��      ໎>�ǈ���3�4���ϟ�����g�C  "b��RX�a߫���ˌx��A��ʵE������|5n�p�#�      ��t���	pZ�.V= �"p`.~^=��5]ܹu5^~�Ң���ǝ[Wc��      ~/�MD����r��6 �e 31�I��ϕ�����>VO9�1�x�Z���      �F��\=N'���	 ��; ��|��6"|�U�^~�R�v���^v}?�y5���W=      �������Y���w�7 �W�*� X�O.���7�ˌ�/����    IDAT]��TO97��޸/?�z
      0���Ch�޸�'���{��5�����u��޽}������1v������461c443ʌG�0�W#ED��`��H�m����m"�r��͈DJ�&b2�}�Z�V�����E�>�aw�CU=���Hv�v��W�vתU���� ,w @�X�NW����_���S�ų7�+ۑR�      �6W�YJ)�e��S�3  ������WȰߍ|���wk���+��=���      �۵ౕ��ӵ  ����J�� ���A/~�����K��[#w       RӍ�ݨ��%E�p� �0p���_��("������n��^���z����5��^5r     �u�[��,�Rʇj7 @��; �u���j7��v7���.D�xs&"��A�te�v      PQj��z���<R������� � ԕ���������>�b��]����l��       *j����\:��3� ����J����������u��!�{f3.�kg       �4W�Y*%�Gj7 ��; ռ���\����������{����F�v      PI3�3-�E)�'j7 �WN T3o��"<�m)������EJ���nz��)      @���߬]�$E�h�|�[���f�@5%��x|�n�����v��xT�&����      �����"��X,������� `�Y�PM*�˦Ӥ���/D��%���;�ޫ;�3      �R:��(��� �7�4 ������b����<��^݉��'�=�[��za�v      PA�o���RhJ��� �7w �z�߹/�/oǅ�A팥�¥���jg       �.E3��g_N�õ Xo� TQJ��xt]?5)E|�s���x      �&����X,��K������ `}YVPG)/�N��z�x�UWNS��ċ��kg       ���2h:���� ��2p��=s�;"ŏ����5)��>��&�NY9�l��֠v      p�R���B[.�3� X_� ��~���N���KW�c�߭���^�����c      �n��'>��J���	 �/�* �]i��xw�w7��ΰv�J�v�x�7�      `ݤN/Rw�v<TJ�W>�͝� �'w �_I/�N����x��V팵pqk�<~      ����T;�^�n�~�v ����s�̵�\�(�y��Ӥx�s��4�H9//^ގ&��      �JӉ�sŝŕ">^���d����G�������^����?E��m�y�     `�_q7�ba}�v  �ɫ# �W�O�N��v7�qygX;c-]�݈a�[;      8O��4p���Oĵk.�p 8W9��vo�Ӥx��N팵�R�K�������j�   �NJ>�m9�M��"JDD��˓z�Ž��;K���a|�?x�_o�����SDJ��ٻ�����1   N�ߌv:�(m�x��s�����[���b����|��/�(����{��v���R��F/.l���v
  �
*�������˽?%Gyӯ���C�gX|ʚ�C�tw�D�;�O�� ��?����E���  �4�hۑ'�k��[���υ�; ����s�D��ka�iw��v��3��.mŝ���C�   <T���������w�~o��hW�W[����*��}��ߖ���?�0|词�  �I�mDL�yV;ޠI�g#��jw �^�87)�_���[u�ﹲS;��^'.�n�����)   �<0\�m��F����s����������:�O�����9�u��:��1|��b<  ��i�;��7jg��R>QRDr��sc��9))����+;�뺢�H���7_�D��?   ������<^�w}�}���Si���}�O�[��m"��������t\�  VV��#u�Q��)pOJq��+���^�7��n`}�p.�{��~��x�vo��ыg��3x�n��+6�?��N  x'����x�>�7jwy�ww�J��!�[G��d��=�7wG���  �PlG��;<�ݼ�OD�p~�8'��x��"^��];���za3��Lb�~   ��ܿ�o��윏r��Z۾�>=p���|:�-  ��JM7Ro#��1,G��g"��jw �>�89�/�T��]�݈�����Ӥ�za#��Q�  `������!�Kr,��O�����0���{��1��;  P_3؎v6	OAcQ��()"yC�saj��{�z��g�ݏ���)�v������K�E�s���7\q  �^)'����e�y�v�;k���{7R�d����   �)OGQ�^���4i������jw ��m��]�z�#aܾP^��eܾ�&���a���?  ����;d���}Cv��D���\~O���7���vN����  �hz��NǾgga�����0p�\�p�Rz�v�m�qigX;�Gtew#�nF�=�  xL%_co�Ǻ�����x|��CN~u"E�&R�w����<  ��H)��N�ɭ�%%��F�S����V �\*�CV��=W�k'���&.��ۇ�S  �E��7��K;s��E�(m�y{�W'����7�߽I  <��F���v
D��hDI�� ΜwR8SW�}����߆�9���0�{u�v�i:�����(�&   "�/���(�ɐ=�"J�]��to螚�� ���m  <\ig����3 ""�4�������w�; X}.�p�>���I)�{f�vO��m��� n�N  �[�Q��ɐ�evXn%"ώ��<��y`���Gj�F�  �=�Ӌ�݈2��g꛷�OG��; g���3դx����pyw�nS;�'t�¦�;  ����'��{�فՖ���ߟG�{��=p����ݐ  ���w�=8�Op�����"⿮����n( g��_w�M{ߍ�K�S�]�R|�{.E�c������q  �����v�������N��w�яH�� �u���Ljg�������K�^��.`�����y6�$���Ջ��+��;  ,���٧'���xT%�����:�:w/��]y ������F��v
k-�\�h?���.`��pfJ�WRy�g�Ӥ���Q;�Spqk�ib޺�  ˠ��7�� 8M��2o#擓���W����wW� `u��`;��v��\��Sa��3p��4�|ƾ���6]o_)E<�=��n�N  ޢDi��>�(>�
��������ԉ���Gө�  <��ۈ��#��>SO)�r� V�gUp&����Ws��aY]Q����}��4�䯊ɴ�����Q;  ���F�O#�YD�.u"u�'�� `�vy�_;�5VJ�E�u�ƿ�Wwj� ��\p�L��J��ڞ��iܾb��Nlo����U  8w�=���,��F�F��<.u���w�  �$�_���'�SXS)�^�g~."���- �.w �Fi>QjW��n���;������Cw  8%�#ڙA;��Je���4�{��S��ܯ  �E�v�����SMI�w ΐ�; ��G��u����t�uwyw���+��� �v� r�  ���O.�_i���.8_y%ϣ��ǿnzo���  ��D�oE��.am��k �ڜ� �Խּ�rD���Xg)E\�٨���4)v7��3  `%�v�� ��h�����Ӹ "Ϣ�ƑoF{��h�7"OGQZO� �ښ�VD���`m������׮ `u����K�sW��K;����*{fg�FG�3  `����J�Q�vQr�"�%Q"����C#"R�ӿݽ1� �s�R4Ýȇ�j���J�s�LD�O�K XM� ��R�/�nXwWv]o_u;��v����8  �nJ;;�Ϗ"��� ���(�I����שs<v�#u{��� �:H�aD��Nk���R*�w Έ�; ��k��?+�W�c�]�İ�b֪K)bw�7^��N ��S��+��#W��Ci���Qf�h"u]w ���w#��#�s�9_%�/D������kj �bR�s��������[��	  �0J;�<E;���w#ފ2;4n����{�܎v�Z����GQZO�  �Ӗ�n���SC�z��� �&�8U%�����A7��������~t�m��x  �Q��Σ�O����� x�<�2�E�D����{w�ۏ�T�  �^3؎v>�A�]��~)"�m� V�� �����g#�õ;�����8G)E�� �:)\~�����(��q;�2)9��0���㿗{�  <��D�߮]�z�D�  V��; �&���זj��&.;����~�  8[�=Bފ���!dB,�>�t��h�7�L���  �R3��o�[��g>��/Ԯ `�tk �:R�_�H�z��D�?�����GJ��. ��S�<�le~�g�s 8/�4r;�8���"�����H�g ��h�;��7jg�FRJ�No���k� �Z\��T����lF�O��Xg�v6j'PA�I�5t� ��W�<��A���ȣ�(��v�u�gQ�^�<�;~���N��4"|�  &u���~n������ ��q��S1ߜ&Jڪݱ�����;�3�dws��?  ,��΢�'Qf�����`Q�6�le6�H����a�n�v  ,�f���("r��D)铵 X=.�p:J�B�uvigX;��v6�0 ��Q�i�ɝ�k���(ӑq; ��d�oܿ����?  ��t"ܦ���T�s����Gjw �Z\p��}�;�t��E��Ӥ��5��AE�~'z�&f�+  ,��N��&Q�G�� ��7_v��/�wz��  ������0"�k��&J�."�}� V�� <�go�/���XW���4�v�mm��-  ���y䣃�K�7�Ǉ�� ���F��"��]v �H�vkG�FRI��n `��p
�j��K;��	,��~�  �?j�E�E��p�N.���~����GQ\� `ͤn?R�ϒ9'M|����/�� `u��t�_o"�/��XW�nl��3X �C� ��mG�F� ,�<�2=�<�;�OG%׮ �s�v�<��"�ݍ���; X^� �T������jw���[��	,�A����v  ���#OG�CA�v �E�E9z=ڃ�F;�evh� �jk:�[�+X95� �+( �Jj�j7���<`�w  �T�2�D>���kQ�^�ȳ�Q �d�i���h^�|x+�|�v  �����x*8g/����8�� �>_;`]m�1�ujg�@6�  ��2? �n �*z����N���  X%)��n��AJW��L|�v ���� xbW�}�Ǣ����XW]o�M\p ഔvevx<f/�v ������Qf㈦Mo#Ro�܋ `��n?Rwxr� �N��+��� `�yG�'֤����w�d�ߍ&��  ,���L�ю�#����}�� ��<�|t����'�  ���n��q�R�O�n `5x��+)~�vú�tc����`��t��  <�e~������ND�Վ�R��''_+�"O�D���Q  ��Ri�U��U��/~���jg ���x"W^���%~�vǺ��z;a� ��(�,���Uڛ����(m��8�h/��(�CO; `�4�͈��9S���/׎ `���D:���nXg�y�a�R  <Dɑ��hG{���Qfc�< xR�4���ɇ�nGi���  ��h���#Xq%���n `���DJI�V�a]���:�3XP�  �I�O#ފ��(G�G�y�$ X!%��0����Ȧ#  `��N?Ro�v+,E|��Ǿ�S���f��c�������jg�W;����FJ�+  �.����^�|x#�|�v ��<�r�����[Q殺 ����ND2㌤ƅ�/�� `�y��ckr�V�a��l�k'��R��\q XO%�|��f���k� k��kr><��^���f  ,����᬴�_�� �r3p�	�/�.XWMJ�5p��w6�uj'  p�J�G�ܹw-6ڣ�I �]y������N�<�]  �z��8��OǇ�n� �3p�<��~2"~�vǺ���iR�ܠo� ���(���ȣ�(�qDɵ� ���Qf�ȣ�hG�Qf��;  u5�݈��gN_��x�ʳ�P���e��cɑ��nXg;�>Aϻ���  8+%G��N���t� �Q�E��v� ��RӍ�߬���J�/�N `y��J��mox��n�s� `Ք�4��h�������N �Vy���f��� p���vD��E��gk ���xdW����"�}�;�U���F�en���� `5�e:>��~#�|R� 8+�Q�Û�_�����k �.R�f�S���Ry��O_�p� ���; �,5�˵���f�vK�iRt;^� ,���"O�D{���k� �NJ������;��   �^�#u��3XA%ů�n `9Y>�h^�ލ_���ζ���	,�^��< ��RJ��a������(�qD��
 �+G������V���v  +��)�-E��� XN^� �H�\}���l�u�9��N`�����	  <���'��_�<��g�� �S�ȇ7�߈2�DD�� �*j:�[�+X5)����W�v ����G�4����Ӥ��yt}� X�2�D;�y��Z; �h�i�ɭh�"OG��  NW�ߌh<Y�ӕ�ޫ� X>�O ��?���(�˵;��Ơ)ծ`��\p X<�D���Gi�[�v ��J�����w��y�"  VF�f�[;��">_���c���j���#b�v�:���<����2 `Q�<�<���k���D��v �r��8�h/���(��A  ����E�m��`�4��~����� `�X>��R|�vº�tk'�dz�  Օ�4��ȣ�(�qD��I ��j�"ތv�e6�] ��k;��95�i�# X.�O ���\�.��O��Xw.��:�T; `M�(��hG��oD�� �(�"OnE{�Z��8"J�"  �QJ�wkW�B�H��� �r1p�Mc�jD�kw��^��^חl��  ����Q�{�'�#�v ��J����k����b� ��I�A��v�"�O<���S;��a��;K��j'��-��y�N�w �3W�<����ԣ�#J[;	 ��F�D{����=�. `�4�݈d^�i(Mt�֮ `yx�C]��_�`D�H�u7�wk'��w �3S��ȇ�"������** �����}/��ND��<  Aj��o׮`E�h�P���a���u�W#�B�����;O�i�� �T�ev�h/��(�I�" �ǔ���ǯg&���y�   \�oFt��3X)Ň/���T���`��C��J�r�
\p��u/�  NEɑ�^���ȓ��` ��;��^�E>���� `�5��p�S�)�ޫ�# XVO ����/_���ݱ&�]_�y2M�& ��(yyr;ڃעLG�k' ��2�D�G;����� `����U;�U���k' �,� x[9�Wk71�wj'��:��; ��(�,��ȣ�(�È(��  �^{y|#��Cw  ޢlE4�>��I)>z������3p�-���?ۊ�_��A�F�<9� Ͻa�x?�|R; ��vj� ��H�/Ԏ`�uJ��v �����(��_����D�y
�� ����Q����  2t �MR���Y;�%�D��j7 ���x;_��1w��y; �;)Qf�ю�"ތ0� x{��  <��D�N��Y*?y���3 Xl� ���k�~)Ry�v)El��4,� ު�(�q�{�'�#�v �r�7t���ծ ����^�]�rKm���� ,6w ޠ��W#�ǭ��׍d��SH� ����Gю^�|t'����  �S{y�o� ��R���Q;�eV�k' ���x@I%�wjWplc�z;O��R; ���F�܉�`/�� ���E  ��� `�5Ý�dzƓI)~��O��kw ���� �.��]    IDAT���>�������;Oɾ Xc%Ϗ��(�qD� ����{>�e� �NR�`�vK�i�_�� ��2p������nྭ��;OǾ XG%�#ފ|o��U �y(�����vDnk�  pRo�;������� ,.w ""�k߹�Z��c)E{�<�R�� ��q|����}>�� ����0��^�ɝ��):  ���F$4�@���?�P� �W DDD/�#b�v��n4M�����o �Aig\l?�� @DD�(�q�{���Q ��R�`�vK*w���n `1�)�߭��}��yz%�� X]%Ϗ���}� V�2=�v�Z��(��U  +)�6":��,�r-�# o� ����GK��>-����;O�a, `��b�a; �r(9�����E�y ����N���R�K�?=��� ,�* ���?���m�yz� �*q� `�6��V�#��  VMj��[�3XF����	 ,w�5��W�|PJ���ܗRİg���+� ��{�v� VG>~*O;���ծ ��4���N�v��W����d�v ���`ͽ���Ո�R����n4M��  U� ���(�x?��(y^� �S�^�4K�����jg �X�� Xs����n��6��s:rv� X>��� ��2�D�G�܉(�v  O��Dlծ`����f� ��;��r�/(��x��h���Sb� ,�{�����  k�D����E��"�{[  ˪�oEt��3X*���}����+ X� k�I��""����6��	���� X���.� Qr��ף��# �2�/�i�*�ԛu�/�� `qx����ʟ"�Wjw�FMJ��w���WJD.� ��m���v  ���!��(y^� ���t"�jW�DR�ߨ� ��0pXSwv��"�j��hs؍�>��͹v ��+9��A���(�q�  ];�<ڋ<�Q�� �L��VD�_;����+���Վ `1���߫�[mz�X��v `����E�D�,  <�2;�v�y:
�% �G3܍W�x$���# X� k�W�����X��jsЭ���p� X�D���/�O"��  �P�Q�^�v�e>�] �#HM7�`�vK���R�u�F ��Q.���H/$�9-�	w ��r��f9z=�� pJ�<��h�7��y�  �E�ߊ��kg�R��.z��; ���`ͼ���_���[�{��u}i�t�� @Eev��^������ `U��ȣ�ȓ;>P	 ����n��ǣI�S� ���� ��Q^-����6��	��\���W�Gю�� 8We6>~r�t\; ��HM7��N��AJ�|�c����3pX7)�~����W;��; p�J;�v|#��͈<�� �:*9�ѝhG�QZ�I Q�oFt�3Xt)�۝��kg P��;�y�7��R�O����m]p����G2 g��y��[����v  D�Y��ݧ
y� `�t6.D$�5�Y��[� �˫�5RJ����&������� g�ް}�e>��  oQf�ю���k�  ��D3ة]��K)}��g��C�; ���`M<�ϯF�k�;x{[�^�T��U2�� g���G�G���  ,��#OnG;ڏ��j�  p"�6"u��3Xl���ߩ@=� k�D���;��5t���5�� �i*�/`N"�� �G�g����'�#���  A3܍H�k<\I�7#���`M� ���u�4������9m3��SRf�h���  Xz�>�9;�� @j�G��)��\ze��� �a���M����[����R��[;��fWU��S�Y���'�"J[;  NGɑ'���Gig�k  �Z�#u7jg������� �a��J�o�n��6�h�T;�RJļu] x2%�#ފ<ޏh��s  �l�Y��' T�w"R�v�D������� �?w��«��@�x�v�5��N`�� O��ȓ;�G�Q��5  p.��������  u�&���,�T����Wkg p��V\[�?�����;�mf� <�e:�v�e6��R;  �Wi��btx+"��k  �N��#�6kg��R�|�v ���`�]��?ߍ(_���;3p紹� <�2�D{���ND� ��V��k��q� ���v"R�v�郗>�?];��e��º���#b�v�1�F�q`��e� ���΢߈<�Q\� ��r�;юoD���1  �#�h6.֮`A����n �|���k݉H�_;�w�z;ga67p �^��ȇ�"��#�i�  X\�4�h?��AD��5  k!uz��۵3XD)�x�c�ܩ���1pXQϦ��G�������l�k'���殰 oRr䣃ȣ�(�I�  X%�� ��~ 8�`+����Y�iw�_�]��1pXU����	���\p�l�����a���(S�' ���y��ȓ��� �V���B���fMi�V���� �
���_��H�3�;xg��^t�T;�4��! Q�Y�F8  pj�?<�H  g��D3ܩ]��I�᫟������0pXAMi\o_���s�Jq� �^n#ގ<ޏh��k  `��6��ȇ�|� ���F��v&���k7 p>�V�s_����j����F�v+h��(�v PG�|tprQ�v  ��2�D;ڋ2�� �4�݈d��}%�K/~��f� ΞW  +���DĠv�Ӥ�����s� �S�E{�ez�H ��(9��v�㛮� ���D3�X���".N��Wjw p��V����?#������m{�R�
V�t�i �NJ�G;���fD�A7  ��=r� ���n?R��n�K9�^���g��BG�������mo�k'���3�6 X%G�܉<ڏh�j�   '����-�� NY3؉h��3XM�ЕO��O�� �l����כ������lo�j'���sw Xuevxrr�v  ��2��� p�R�fx!"<&�c��|�v g��`E<�7W?�">P��w��4����r��l�: ���N��G��v  �k�  �.uz��[�3X�.�|�b� Ύ�;��(�Ok'�h�\o�Mf��	 �i�m��[��7"�v  ������G�Oj�  ��f�����`���گ�� ��������?�~�v�fwsP;��sq� VJ�2�  �2+'Xu� ���/D$�7"R��k7 pv|�XM4߬���I)b�w��d��N  NIi�юnD>�F0  ��\s 8%M'��n�
A�>p���� �w�%����GJ�gkw�h6��v|��l���+9�����yV�  8Mw��OnG�R� `i��0Ro�v��I��v g��`��N��""�����n�k'�f��	 �S(��hG{Q懵S  �3t�;�� ����nDӭ�Ae��/\��?~�v ���`�]���"�K�;xt;��� ��J;�v�r�1��  �Ci#�oD>:��� [J�/�{��-E�s���� �>w�%�I��D�����u����9g�p�; ,��#O�D�G�Y�  ��2=�vt#J�� ��J�^��v�*kR����jw p����3׾s!"���<��M�OqvJ���]p�eQf�ю���ƵS  ���,��F���  W�ߊ��Y�ZK���̗kg p���T?�߈��;xt����sv�fmO2��W�<��ȓ�%��  F�|t'��-�+  <��ƅ�ԩ�AE)�7j7 p�����_��A����<��"��������G�B+%��A��~D;�]  ,�2�D;ڏ2�} �#KM4C��Z�>t�S���3 8=� K����W#��<��a?�&��`����	 �C��Q���(Ӄ���  �]�6��ȓ;�{ �G���H���T�6�?�� ��1pX6ׯ79�?��������N`�M�`��6���ȇ7#���  ��)�q��Q��7 <�f��x���ʿr�S��� �w�%���\�|��@�υ�A�V�x2��  �S"D;ڋh�j�   �,�"���LǵK  �@�f�B�ĭ��R/���� �t�j�lJ���	<��A/�]_r9;9���]��EP�����AD��9  �J(���D>�Qr� ������%w�Sʿ󾗯kg ���� �ȕk���ӵ;x<�]o�lMf�(�s PW9�ڞ��ٓU  ��W�hG�QZ�s  ���ۈ�ݨ�A)]����v� ���;���g�x|����	���Ѽv ��2?�v�wr�  ��6��F�#�  ��f��tkgPA�� xz� K�W������<�a��^�v+��� �(9��v�Û��]  ��ez��fDɵc  SJ�l\��T�����+����kG �t��D��'�;��sqkP;�5p85p��Vf��W�g��S  �u�E;ڏ2��. XH��F3ة�AmJ��v O��`	���>�J\��������N`ŕq4u1 �K��h�7"On��  �W�ȇ7"�. XH���;���9kJ�������� <9w�%�F�������ub�߭������K�� k�D��"��#Z� ��R�юo� . ��h���S;���D���3 xrƒ ��o�?J�z��ŭA����Ѽv ���΢݈r�zD�`  ���i���(s� x��D�q1"R��U�ڋ���Y��'c���R��ED8��.�s�� pfJ�|ty��g�k   �]ɑoD��	� �/uz�۵38G)ť�Y��� <w������(��<�^��́�%p�&� p&��������v
  �c+�q��%�N XM+��P�:i"�Q��'c������K��휃R"�w 8U%G>���fDik�   <�v�h?J�T  wu6.D�N��KJ?|�S��� <>w��������߬�����=���8��#���Rf����I�  ��Q������{�=�����|�{fzf�\�93����J\,[ #C�1ج�����肍��H8B�J>��#�Vk�S�8IU*��W�*c�C�r�J*N�S`�d�����t�t��������sfz�ӗ��/xVmU������ݏ<�. ������t	W%��J� ��;��jZ�xDtJw���;�X]vx��w:py	 &��W���)]  0a9���h�GϾ `���R����\�TUo�y�co,���1p�B�=����Kwp>ۮ�sEzg� pQy�j;  ��u�n�f\: ��ji-R�o��!WMt ��`
���C�T����Z_.���p� .��W����  �Gs��!_ ���V6"R�tW ����o���� �?w�)s��O�*"}O��gu�� s�F�&Fcc< 8W� �������ȥc  �IUTݭ�H�K�d)b)uW�f��;��i7�c���r���rz�z; <0W�  ~G����� Xh�Չj�Z��@��}������ �w�)r��<�PD����OJ[k�\�Ӂ�; <W�  ^@=���n�ڿ7 �+-�FjwKgp�ҵN���� �w�)�j��5ͨ����}�r5��>5uԽW�  ^L����G�K�  S�lDT��\�T���ȣwVJw ��� �����s��/���m�����h���t L�<�G}z7�>+�  0�r4��h��K�  \����n�9ݼ˷����-]���0%R�>��Ϭ*��\3p�j��Ƒ�� /��W�G�j;  ��ʣ^Խo� R��Q�\+��e��co�U:��f�0~�S7#���3lcm)ZU*���蝍J' ��r�  ���aԧw#�� X<�Ӎ�q�p�U)}���|G� ^��;����"b�t�w�?p�:'}?,��h�{���  LB���DJ�  \�jy#��������� �4w��n����H�-���-uZ����-W�ir�������a�  �9�D�?���t ��J)��f��ͳ�7�r�[KW ��|V������������	,���8��Kg �t�ύ-\m  �4yxM�0¿K $U��F�̫���n ���t��O>�W���پf��չ�w� ""�x�����A�  ���ǃ�{�M]: �ʤ�r����\�TUo�y�co,��3p(�i�߈�������R,�}�ruN���	 PV������Gd�
  �+ӌ��ݍ<v� X��zDk�t�"WMn�p�
 ^�E@!�����G�w���b���������; �+�ύ)F��)   �)7�����. �2��fDj����T�m۝W�� �K��T��>�gZ�U�ƪ'��:'�a�\� J�ќ݋�w7���  Xp9�ٽhǥC  �F���nED*]����i�_��/eX	P��w=�D��^����^_���W�����v On�Q��Gv  `��Q/��A�� ,���D��Q:�K�"ߵ7=~�t �g�P@�T?�yׯuK'�`N�� ,�fx��݈�w   �T�Ϣ��G4u� �K�:�H;����u���� ������;?�G#�7���b�V:���*����ǥ3 �j4uԽ��g�"�%@  ��֌����p2 0������S:�	K��K;��o�t ������H-���]��R:�s2�� �!��Q�ލ���S   �_���wy|V� ���hu�"���\Iig����� �.ߴ W�ֻ>��#�7���bڭ*�֖Kg�`���� �s�����("��5   <�&��A4g'�C  .WՊje�t�R�y�k� S���ܹS�\�x�.������T:�s�3p`~�� ��g"��S   ��<<�fp�t
 ��I�H��Jg0A)�C�K�{Kw �,w�+����zOD���\LJ���*��F1�]�`���8��aD�]  0/�u�0"� �ZZ�Զ�+U|�w��`�p~�N��z��X]��N�t���v �Pn�Q��#�z�S   ��YԽ���.] pi��͈�S:�	I)>�6�_� w�+�{X����;�������0_��i4�w#�Q�   .S3z����� ��J)��fD2ÛU�?��[*���|�\�G���D�����;����7Wk8nb0�� ���M4���g�"�k�  B���D;� ̧T��Z�*����*�z������ ������z���_Y������-��:N ����aԧw#��S   �rM4���# �)��"-_+����*�h<z�]�`��\���'�#ҏ����ZU�����,�{=W� �u9��q4���\��  ����0����!  ��ZZ�Զ+�)������� Xd� �������\����hU�t�ir��G�3 ��r3��t?�W:  �)��'��Kg  \�je3���`r��bo�U�`Q�\�{O�"��WJw07�uK'�������\: �%��ќ�G4�  ���M�0"��' 0gR�Vw+"��ͺ*�/�q�u�]�`Q�&�$���fD�����u�be�C�\��ްt <��D�?�fpM�   �T��D8� ̛���VDxK����C���a�p	v������77]o��{� ̘<F}z7�xP:  �YP���GdH �%��"-���ࢪ����{O��Ed�pr���3v.�,�ccu�t�w6�Q�G fE���$��~D�K�   0K�ѳK7��%  U-�E�8�7��P� �+�`�n�}�OD�7��`2v�VK'���N]o`6�f��~��I�   fU����G�G�K  &�Zو�:�3��*�ޝ���Jg ,w�I��ǭ*�GKg0�v[k˥3XP��g� �e�� �����   ��M4���c�? �y���݊Hfz���Zq��j�������_���.��d�l�FJ�+XD��QGu� x	9��q4�ÈhJ�   07�h��ǃ�!  �S���nG���J������� ���`Bv��X���Z�&�U��qm�t����v �Wn�Q��G�J%B�8    IDAT�   0�r4��ȣ~� ��I�NT+�3�����n X$� �R|0"*��d���FUyz�2�z^��tʣ~4��ͨt
   s�� s%u����Jgp^)����~�w�+b�07����#��Kw0UJq�Z�t�w6��.� ϗs4��hGє�  `A4��h�NJg  LL�|-R���gV��q���
����V������ؾ����H�8<9+�  ϓ�qԽ��cW�   �zyxb� ̕je3����|��ƛ��*��� .h�=�xC���;���"v6]o���Sw �G��9ݏhF�S   X`yx��t �d���VD2ݛE�����V��y�[����\����r,w�礌��(F�t D�M�(��QD�n  ��<�E�?��\: ��VTݭ�H�Kx@�J_�}�U�_�`��\�λ>��H��L�Ζ��sx�z; ��zu�n�q�t
   <O������ZKQ�l���R���#��Y)�0���k��RN?]:���X]���N��ᩁ; e�a/��~D3.�   /(�Q�#��; 0�R���Z:��Rz��J��� �����n��}_D���Lέm4R��`�qS:�E�s4��hΎ�<   �^}u��� ��ʵ��r�P���;��o�t��2p8���'�s�/����Ni��PJ�GQ�>y<(�   ��� s"E��Q�K�� R�����/�0���#����Jg09��SR��'� \�<�G�ۏ�u�   xpF� ��HUTݭ�d�7SR�?���ǶKg �#߈ ����^�">P���q��Ҏzg1��� ,���8��QD   0��aԽ����X�ٖ���#�H�S�O)���Z�� �����T��X)����Ni�� X �G}�y�+�   �ь��� 3/���Z�(����⽻o�Э� ������{�[#�w��`r\o��q�Ľ��t "�Ϣ��G4��)   0YF� ��H�n����ܷt�^j�t��1p�_��i�?_:��r���N�"�� ̿��I4}?�  0ǌ��9Q-�GjwKgp�r|����<R:`��ܧ��[��_S���q��i�oP:�y���{��'�K   ��� s��nD��Jgp?R��r��� ����>�r����?V���r���zg�ǥ3 �c�F}z7��N  ��c� ̅��VDj��>��}�m�=�; 慁;�}������;��ۙ'��py�M� "ץS   ��� � UQ�n����K)u����; �o>�������F��P��ɺ��V:��s���Y� �Q����9;��\�   �1r �@��Qu�""�N�e���Ν�?��� ����eT)�|Dx���Z[���v��q�,ƵU ��\��>}&��[B    "�����: 0�R{)�������8w\q� w��pk�w�o)���q����w�z; �G�hz�.�   ӥF�?0r fZ�t#uVKg�2������}��Kw �:w��ʽ���U���L֍�n,w䧬q��q���I����E���   ����^r#w `vU+��+�3xi��T�t��3pxô�x����LN�J���if�ۿ7p(���MԽ�ȣ^�   �~�Y�=#w `�U�͈�R�^R���o��;KW �2w�p��O�*"�p�&kgs5:m_}���q�t s ף�O�F���)   0;�h�Ga� ̮��VD�.�K�Z?���$�9Y���v�~."���#�V;���ǽa��M� f\����G�t
   ̜<<7r �Q��������U����|��Jw �*�p _��;��c��L֭�kQU�t�]������8��Ks   py<x��k �ٔ�vT�툰��Z)}x��.�0�����?n59�|�&k�ӊ��+�3 ��&����3 �U���wy�+]   s!����Kg  �[ju��n���E�7[���Kw �"w�/����O"�Jw0Y]_��e����~d�v8�\��>�Q{P
   &)�z�OKg  �[j�DZ�V:�������ï*�0k��s�;�ܭ"�F�&ku��k˥3 r�ؿ7(��ʣ~4���\�N  �����Ezc 0����H��������~�t��1pxN���ۥ;���o��N���8<=�qݔ� `��hG��"�+@   �25gǑǎ�  ��Zو�^)��I�=7���?P:`��D�����]����Z[���N��������	 ̒�D}�y��   �J�?�<��  8����Z*���j5���� �����;�鉈H�S��*��}��v�C8����t 3"�èO�F4�;   �j�h���k� �*E��Q�K��ER��t���S�; f��;��vww�)�P�������r�U:""����p�M� "ץS   `A5��"7��!  瓪hu�#�i�ɹ�h��� ��b�B���'^�>R���괫��\-�Q79O�x99��Q4���ȥc   `������ 3�jE����)���~���-�0|����ߍ���L��7֣�R�����{��CE ^Bn��D�K�    �����)] p.�Չ���S%ŝ���\mx����}�o�H�Q���Z�vbkm�tDDD��;�� `��z��݈zX:   �b�8��ax� 0�R{)����|���+;�?R�`���{�)�t��ҳ��aZ���h� /,�Ͼ�<{�9   L�zM��t ���N7���|�����<�#�Kw L3w`!���㵥;����.�Kg��p���O��F��   `��� ��q� �s���"-����wm�++?^:`����>�U郥;��v��[[��3�w��G�?�� `��M�0�ٽ�%   �ȣ^4���  �V-_������R������[:`Z��j������L���k�n�Zcz�����MԽ���A�   ���=� 3��nD�Lf�A�Xʭ�S�`ZY����o/��du��q}}�t������ްt S$ף�O�F4��)   �4��ȵ���Y���݊h-�!"R��v���?,�0�܁�q���ZN�o��`�^qc=R*]��i���y4������)   ���h���q� ��Iύܫv�"���g��{�8 �"���H+g="^Q���ھ�k+���;F�&O���g5g'�#"�N   &%7��"rS� �|R��vDj�.YxUJ_��ʯ��� ���X��>�5)�Kw0Y�V__+����q?�# 9G�;�<<)]   \�\G��P; 0êVTݭ0!,/��C;����� �ķ� r���dD8�=g��햯2�G��ؿ�z;����8��݈��t
   p��a4���  �Z��V�""�NYh)��fy�'Kw L����n�ňxo�&k�ۉW�X/����� �N�Y����"r]:   �
�8""R{�p �����Վ<�[wQ)�a�˾���ͯ}�t
�4p��k;{O�N9�T�&�J)^y�Z�x��#>w�+�@Ayԏ�w���)   ��Ó�#o� fWj�D��Y:cѵrg��KG Lw`��T},Gl��`�v�Vc��%$L���A��� ��9;�fp�t
   P@38�\�Jg  �[�D��Q:c����[?�]�; ���;0�v���?���t���Ԏݭ���<9G<}�z;�b���"OJ�    E�h��M]: ����j�����I��>�u?`,<w`.���_��|�t��ʛ�R�
x���AG~� X8���wy�/]   L�\G�?|�*
 �����#-���XX)�Wvn=^��4w`.����L�*��d�����J�t<��� �)7�{���t
   0M�Q4���  R-_����XX)������#�; J2p���'�`�齥;��N����{B��sp2�3��J���G4��)   ���A4g'�3  .�Zٌ�^)���R�V���� %����;�&�"�U:��z���hU�t<��� �'����"rS:   �byxy�/� p!Uw3��\:c!�������� ��s���ΏF�ז�`�6V�bs�LL���3��Hsv��+�s�   `4�����t ��hu�"�N�E�r��swl<�����;���W�>\���jU)^q�Z��9G|��t W"G�?�<�jq   �A�h��� ̶����m�^BJo�~��Jg �`�̉�R����n�&����u��q�`A�&��A�W�   ��{�p �LKճ#��*]�p������m�� �j��\�y�'�7R~S�&�Zw)n\[)�/���^� .Yn�Q�ލ���S   �Y֌���  ��TEk�����K����/]p�|� 3���<u3�濍���-LN�J񚇶�U��)�%O���K� �,����"�+�  �	h�)Ej-�. 8�TEj/G�j�R�˯���~���ߗ.�*.�3oT�����;��WܼKm_SL����0��xM߸   ��|v/���t ��������d�qURJ����xD�	,�2�L��{�m)�ݥ;��͵��^_.�/���,�q� .I�����#   �eh�G��� ̶T���n�_���7�x�G��� W�70��SO��*=Q���j��xō����r�����3 �$��8����   �\k�}�>{� �m��yv�n�x�~�ڛ�Q:�*�vfָ��D�xm�&�7ף����tz��Q]:�����#�z�C   �EЌ����  ����D���t�bHi��j��� W�U: �<n����9����\�Z_���k�3��M���q4�� ̗�<��r}V�   X$��c*��T8 �bRՊ��D���*�*�q��������v���d
̜�x�/,�����\鴪xō���>wԋqݔ� `��:��~D=,]   ,�<<�<��  ���^���.�_�VT��wl?���C�9����Z�x}�&�;ע���t����a�t ��QԽ�͸t
   ����qd�> ́�^yn�ΥK���o��� ��#S�L��{�kSJ�kDtJ�09ׯ�īv��΀��gN�;����a4�È�f   `
T�h�ވH~� f_���Θ{9�3æ������.�p��fǣw�)�/�q�\鴫x��z�xQ�a�����E����q;   05�� 07R���F錹�R�\��?]���3cww�F�7��`rR�x��F�*I�^�=8��KW 0	���s?�`   �K����  ����i�Z����?�͏K���`�̄��|����L���j�w�gz��FqxzV:����#OJ�    ��|v/�ؿI �ZZ3r�t�ʭ��bo�U�`�܁���v�_����)L��J'nm��΀���}�r f^�Q�#�z�K    ^V38�h��  a�~R���G_��Kg L��;0�n��~0����;��V��ջ�R�xqǽa��G�3 ���D�?��]>   fDn��F�\� `"�ܯ@��k7����Kg L��;0�n���刏��`�^�s-�ھ��^9��0�ru� ��.   x0�(��q�
 ��1r�\)�ͦ���Kw L�u!0��ܩZ��#b�t
�sc��k˥3�%=s܏�p\:�s��8�ӻ�7q    �)���b 懑��J)��ƛ?��� �b�L���������L��R;��V:^Ҹn���^� �)ףhz��.�   p!��$r�~ `~�_��������! ��* �Bn���_���/#�S��ɨR��<�Km_=L�O���� �(��hz�єN   ��<F��F�T: `"Rk�������S�O���kۣ����_-�pQ.���Ν�ʭ���)L��7ף��.�/�?���~� �!���¸   �+����t	 �ĸ�~yRj��[~�u�; .���:;���_���t����7���΀���'��F 0s��z  �yU�9;-] 0Q��Z�����'�J��'Kg \T�t ����'����X*��dt�U���fT�Wg2�N��sG��̚��$��^�   ��U#�:�*o� �Gj?7��eC�MJ�t_��?���_�?J� ����ɩn�/G��3�DJ��ڈv��ӭir|f��t �9�y��   X��(��Kg  LT��i�Z��Su>����� 8/�C`j����_N�t�����X]�΀���Q/F�t �-G�?�<�jn   `��&��aDΥK  &�ZZ3r�����r��\���j� �����O�6W鿊���-L���r<|�1~��٨��z�^�9 `F������t	   ���MDΑ�˥K  &*��"R����S�GJ_���?�/{�����t
��r�(�Ν*W�#�zN,wZ��O�2>��k7 �!7Q�"��%    ��Q/�_: `⪥��V6Kg̓�T�/�z��J� <(w������#�)��dT)�#�6�U��)�N��8:5��	���w�j   @D4�����t �ĥN��}�R�׌�ʏ�� xPև@Q��>�����ˈX)��d|٭��Z�ZL�_����b0�N��|~����   �wT�h�ވH~� �O�E�7�_T�yT�?��?����t��r�(��;��?
���qs�k�����Qϸ`4uԧw��   �X3�fp\� �R���s��=�wQ)�N^j�b��J� �/w���[��)}}�&cu�__/���lT�gz�3 x�G�ۏ�u�   �����ȣ~� �K�:+Qu��'"�7^?�=?T:�~����y��oLM�_"�S���k����WlG��)f�o|�(����3 x	�E�?��M�   �)WE�v=R�. p)��,��aD��)�-�ɸi�p�O�ߔNx9���������rj���s!��W�^3ngf���L9�v   ��D�?��_ �|J�娺����Xo���� ���r���?_]��ɸ��׺K�3ྌ�&>�Z:�����hz��    �Esv�t ��I�%#�	HU�7������ x9>�+����o�����h�n��6V��5�7Kg�}�wO���Y� ^��K   \L����R: ���zM�0"K:�����W��GJ� �܁+��zj5���q�\X��ջ�3����� S,���    ��#7��  �&���Z�
���K)=�Zk�L����S�2�n�3��+Kwpq�*�#�6�Uy��nr|��f�Vyԏf`�   pqM4����, �<{v��痪���x�c�Z������ĭ�'�5"�W���x��Ft�ڥ3�}��I��^O0���i4���    �E3p� �o��1r��V�:�x�-X+�B|����������?�������X]*���^���3 x��4�[   &-�z�G�m �o�3rOf��Rz͸Z��� /�';p�:���GīKwpq�k�qk{�tܷ���[�3��F��    ��9;�h��  �*�:Qu���-U��~���t��\�[������[���[Yjǫw��΀��'17�3 �"��    W 7Q�#"�. �TF��J���{�7��n��/��4����ݜ�S�;��v��GnmDU��)p�������W�Msvb�   pU�Q4g'�+  .�����*^��X��; ��Os�������V�.&��/�݈�N�t
ܷ���[�3��6��I�T   �R�F���  �t�Չj�zD�qyP��~h�͏S���3p.��>���'Jwpq]_��n�t<�O}�^��M� ��q;   @9��(��Kg  \�T��Z�6rp��j��x��\: "§80q��z��#��&"�J�p1��V���k�3�����Ӈ�� |�fpytZ:   `����8��JD��1  �*�*R{9�x�t��Hig�Y������t
���d=z�M�_D�z�.fu���y�t���z    IDAT<��Q���:0�4yv���#   ���a4g�  ���K��#���HU���?��ו� ��L���ΏE�o(���tZU<rk#�̐�#~��{Q7�����    �%O"���3  �D��Qu��L�����fi���;��-�b��L��w��#�c�;��*�x��Ftھ"�-O��w6*��s��   �S38��M� �+�Z��V��D��k�/�>T�Xl���|���?��Ɲ��[��W�n���R�x ��Q����� �9��(�_:   ��#�:Rg�t ��HU+R�y4(�23RT߸������??]�XLK&"���\D|U�.���jl�/�΀�49~��{�s� ">�ݸ   `������  %����nGD*�2R�T��{{�(E������"�_(���l�-������>u�$�Fu� ����^�    �C38�܌Kg  \��^���F����?�}��)�,&���������&�����]����.��+ڊ���l9:=����� �q;   �L�:�Z�� �"��A4���������������O���)�bq���&�1��gZ�U�#�6�ۙ9�q�z�t a�   0��Q4g�� X,����F�ِ����"�ؚWʇpn�����Gķ�����������u����3�b\7�3 ^svb�   0���4�xX: �J�N7�e#���R���>P�X,���r��xmn���J�p~��ڈ͵����>wԏO�uQ����$���1   ��K�h�݈H�" ���F>�W:c��<h��?x�?���]:X�:ܣwڹ�%��g�C�׌ۙI��Q|fߘ�4�v   �9��hǥ+  �\��ii�t��Ki�j-��x�N�t
�܁����c�Kwp~[k˱��Z:ظn��~�8r.]�،�   �O"���3  �\���cG��u�;�GJg �!� f��;������#�U���Y[�ė?��7 3�7>s���� ͸   `�UQ�]�T9�	 ,��y<(�1�r�0��|����V��o.��m{�͈�+a�>�:�*��a��L��Aϸ��fxj�   0ךh�G�U� �⩺����S-E,E��y��J�`����S՟��GJwp>�*�knoF�壟�s��gOKg ,�fx��^�    .[3��̿� �(E���Z*2�R�}���(��7+G���=�ݑ�Jwp>)E�zw#�K^'�����ͧ�#;PL���   H�D{�* ���s#���楤����o~�[Jw ���xY��>��H��;8�����ƪ�K�=9G���cT7�S V��9;.�   �kGٿ� (U��nG�V�i�j��_�y�}�C��d���G�s�~%"6J�p>77����-����N�?*����x���   `!�ڿ ��jE���L,_L���z���*��'���Kڽ���H�Kwp>�K��uJ2��{�x��W:`a��0��QD��)    �ǃȣ~� �"RՎ��f�/.�Z߿����x�`������}����yDx���.��+ڊ��Q������~� ƵW����Q4����9   @���HU�t @y|M�0�za9ǧ���~��[����"�m�=��%��gR�U�knm�3�r��w�=6n(ĸ   ��k�� Xh����f錩�R�������;��b���N?��������yh3:m�̦߾{��Q�����q4}�v    �H3���t @1��i�Z��UU���������~���;?��"ҟ-���K)��nmDw�+"�M'gq��_:`!�f����l�   ����y�egy���s�]��Y�Ui�R��W��Y�L��a��,a���V�m���{:c��nT	am6H�3��тl�D0ƍ��``P-��\n.w?�3��T��*U��y����`��D��y�x<o��3�  �ޕ�d���ye�ŽS?���! 6��fz��;$�݁�ٶePC�R�`]j͎:�; zS�n�b�       �\�Q��c�   D��Ii9vF>��:���� 6�4v ��=W�M�]�Sp���55�)Qt�v'���%e�/�`�yPVg�      g���.+0�  z�))��;-nF~f�C��_�P}�}_��������MMM��L/�݁s7:P���@�`]ܥ�/��� l8�j�R��.     @��v��@  @�2S�?&���PR��#/{��3 t7�H�&߰�j�~?v��@_Q�N�� ��+Zk�cg @�qx��g0      �MhT�X
  z�%J*�b���l�P(��fg9 `�x� ����2�)i,v�M��j�����N��D���K�� Ѓ\Y}I
l�     �z��AV�  �%�,-�;��)�c��������B� ݉�C@�s+��.�]�sSH�Q!�Q���h���j� �I�^��f�      t1o��  =�
%%}ñ3�)I�>����0v���w��M�N��Lo�݁s��i�̈�˅�)���:A�T��N����N=v      6�ZJ�ɸm  �.K��\�ڱSrŤ��=t�~�v蟹Z�9a�/�æg��cn���8w�Li��;X�\��U��B� �9��"o�bg      `���X�]  ]R�*�3r'1ە����@�a�;У���JwI6��fۖAmꋝ�ۃ�W�Z��2 l4o����      �lBG��o.  �]V,˳��Y�\1K~�rŋ�Q������{���Q���n?��fr���N{�{[�ii�; z���
M6i     ���)0�  z�)��J���3�yq����e+��ƀ;Ѓ�g�^'�Wbw�܌��m�`�`ݪkM]\�� =�;M��     ��5��#   �DI���<�i*���o�3 t�
=frv�.�}FR9v��@_Qۧ�ef�S�u��::tlY�K ��x�V�/I�     ��3�L��b�   De��҂�ӈ��+f��|�����|9v����K���h��K����W*��>=�$a�ݩ�:��,0\	 �CG��()�N     @���<tbg   Dg���<;#w�$y������� �pz��R��^�g��&�|fD���5�S��G��jg�S ���L��(9��      �H�P��  ��4 +Tbg䋩b���u�o�c� �7&&�1yݾkM���8{��v��\Lc� ����՚�� �[<(�-��      �h���\�]  �IeXJ��3r�L��F�0v�|cj�[fo�(��4�g�L�ljXC�R�`ݾ7��ŕF� �-��j��s4      "�ڲBY�0�   z�))�坦���Q��v^uom���b� �'6����-i"�����)8{۶jd��xн�W:Y��� ����R��      ��
���  ���J*��,vI���ҏ��~�h� �Ā;��M���ʹ;v���X�&�+�3�u[�����+�3 ������bg       ���Bs5v  @.XZT�7;#W�첤o�C�; �������]m�G�a��1:X��C�3�u�5;:x�*g! l��\��k�3      ��emY�$KM   ��(ɥ��af?ҷ�꣍���J� �§H`�y㾱B���c���V��>="�6"t�V'���%e��v �Hު�[l�     @>y����/^�  HV(K�s�$I&���/��q���c� ��:�T����uY����R��vt�,������) �S��Ph.��       ��g
͕�   ���KI!vF~���P����s}�S ���&4yݾߐ���8;�b��gF�&L��;�K_V���b �H�����      ���vM��bg   �%J*�b|�Qfz�J��G�; �G; ��5}�M?*�-���[��
i��gFU.�8F������V��3 ��x�(�%y�      �x����/�4  ��Y��;��)���?ٿ�%_���۱S �� `���?�H��n��K̴cfX}%��ѽ�/�4�\�� �ŃBmQ��      8{�)�VcW   ��d���9�[�����]�@|����?`�����3�.�R�E��^��MYX�� ��]YmQ�,v	      pμ�&�Z�3   r#)Ji)vFn�i�B�1i��V��� 6��=7���bw��\41���r�`ݖk-}��r� �1���$�v�      `�B�*���   �	SZ�,��������� ��lS�ݼ��N�]`fl@�#����՚m<��w� ��B�*e��      �3t��x�	   I2��%y��$?,��rً����) �`�;�����}B�p�<��>M���� ֭��t���� ��BsE��-      l�Z�g��   �aiQIy(vFn�TR�����<�@�]n���K������/��	~E�jw��YR'�S ��x�.o���       ΫP���b  e�~Y�;#7�l{Z��@i�  �79���&��$�݂��_.j�̈���U�NYp�?RU���N��❖B�;      � N�[��   ?,-�;-�Y>(I2�������_b� �XLZ]j��dZY�k�fb�੕��vmU!��t�\�V��h�N���Y[��(�/�      �y%�㲴;   7<t��{��[6o<�����v� �iK���%����WL]���vt/w��+��F�P__Z     `���   �$YRPR���'�A�O�������0q	t���z������SKӎ�#*xԢ{=trEյf� �-��j��g�K      ��3��j�
  �\�BYV���f���l�=�; l�4v �s3��?%�G��\3�v̌j��;X���_n�� ����KRh�      6N֖J��  �GX�$��,�z�%���w��_������- .<d�.23��IS��
�[��.��`��vt�պNT�3 ��Ɗ�qs      zO�W%��   9bJ�F$c��O\韌���c� ��x�]�-�%]�OmۖA��cg 붰���y���Zk�v-v      �g
-�O   �&I��Ǯ�3mI��I]y=�G�M����.19;�V3�z�<���~M���� ֭���wO��� ���톼�;      �+k�
%Y�(  �#,)H�Ў��vq��������b� �p�Tt��7|��}L�����`YO�� �m��ҡc���	 ̳�B})v      �����*�,v
  @nX�$�N�C�$/�u��j�����- .�$v ��6��}c�ɧ$q�J�V��t��н�m:�p; l4����y       ���Qh�Ů   �SR#���$(���+�~I� O; ���m��\��.�����1="c��T�����U��`cy85�Ζ      �4�Z�g��   �bIAI���0ӄ��S�=W����Kc xrS{��W�~#v�\��j�̨
)�Нꭎ]Vn�����KR�%      �D<�()U$�e
  ��N-��=�$�L��%�bc��w�np~1�����M�w����in�D�ό�\�o�S������:��`��Ɗ�i��       �˃d�,-�.  �+��7E?̒�ŕ�/�r}�}��np��rȡ�׽w4�R���Tb�3��+1܎����?��6�� ��BkMޮ��       rϛ��Љ�  �3��2"�?�/���щ��e[� �O8 w�J��G$�]�'f&m�V�;X��#����`�y�)o���       ��+4�cG   �%%}C�3�dƓ�'�9fb�M���@�L_7�f���O��!��cg ���N���Y� �9���K�<v
      �=<�Y"KY>  �X���9����ʎ������) �9܁�x����R�l����M�Tbg �ׁ�U5Z����P[���      ��򬭤�'9  �
%y�!�l�bI���W}�����[ <3|�rb�u�M<|JR)v�ؖኦF�cg ����Ѫ�MN���se�%�9`      �OP֨Ǝ   �K��ĮȓTI��&w��L� ��@N�J�?����xb�e]<1;X������F;v
 ��P�JY+v      �ݲ��]�]  �;V(Ɋ,�|���f��Ǥ9�c�.�0�����I��݁'6X)�ҩ������:x��v �%4W�F�      `S��C�  ��I����;#7,I^6~Mg.v��Kc �n��=ۂn�T�݂��+t��Q%��N��#��u�� �4����      �&�R�dž�!   9c�B�o��^�w��������np���D49�wP�n��709T*��|fD)���B�@\�����      ����&  <K
��`�<I-)�����.���1�Dd��,�Y�;�x�4ю�<&�}Bp:��p; ��A��$�c�       �Rh,Kbg   �NR��r��0ӄ�'u����- ���@$S�7��\o�݁�K̴cfX}�4v
p�ܥ�/k�ފ� =ʕ�%�b�       ����J�
  �\J+#�1�3�h|b�{bw 87LoLϾ��dv�$N�匙�cfD�}��)�9s��j��p; ���R֌�      l~�#K����   _�dI*�4b��Y����/�F��}ߌ���pL�`��{�$�H��n��]<1��
���>�@|��*��cg       =#4�O�$  �i��'+2��(OT(~x�oyV� g�w`���M����;�x۶j|�/vp�n���Ӑ�Vcg       ��3��J�
  �\J�Ò��3r��F�ʟھ{�1�0�l��={���_�݁Ǜ�hr�S��>�@|:
���      @O�vM��  �q̔�Į�3{�r���� ��s�2}�M?��_I*�n��F˺dr(vp�ܥ�/3� 1yP�-H
�K      ���Y[I�"�b�   �%��A
��)�a��D������k�[ <96�`���h ��"�?vN7T)������9{ds{u�; z�+�/I��      z[�(4�bW   �RR��]ȧI����mύ���1�l o�3�bw�t�墶O�X�.��v ȇ�X���      �o��36�  <����H�|1H���W�e(v
�'ƀ;p�M^��W%�J���TL�}zXI�t;�K��G�� �y�&o�bg       �>Wh,ǎ   �%KK�b�\1�g���ͱ; <1� .����Gd�I*�n���i�]��T*p��%��cU���> 1y��Ш��       p&2Kd)�g  �diI�nH��)�af?ַ�%��~9v��1�\ ���ѾV�}V�%�[�41��:���?t�,��j��p; �䡣P__�       ��Y[I�O2�]  ��L���z�\��~�o�U��8p�wc� x���^�����x��t����˅�)�9yd���d� �rW�W%�K       <����;   �,-Ɋ��3�Ŭli�S��w&v
�G1�\ �����~5vNw�԰�*���9iw��?��p; �@hT���      Ƚ�)o7bW   �RR��>��]��ʟ��l��)�0����?x��?#���ڶeP[��bg ��	:p��F�; z^h��۵�       Βg-%�ʩk�  �(3YZ���Kr���_/���{w� ����7}�����tY�<jz�_ӣ\������?��f;�� =�;-y�;      �9qɃ��,  �3Y�J���LI���]W������f���%��ͤVk�O�scw�QcC}�����G��[�@t:
���       ���uy�;   ���d�H>�'.�ȖW���.z��y2��=����x�pI�L�� �I�����-2� y�P���\       �+�FUr�܂��    IDAT�  �?fJ�FbW䎙�x���mW^���e������]&���x�@_Q�M�,v	p�ꭎYR;c� � 4�\�      t;�Zk�+   r�
%Y�;#w��9�-S7�� z�K �Юk�Wn��K������.�:�4��G�������0� ����v-v      ��!k�
eY  ���P��뒸��4�=�|�����|9v
Ћ�������{%���8��&�|�
������:p��p; �w���j�       �+4���  ��DIy(vE.��������@/bx&g��{�~-vNIӎ�#*x��{,�Z:x��,��* 䁇�B�;      ���
-nm  x"V�Hi9vF���--|jr����NzS��:M]w�N3���8%1ӎ�UJ��)�Y[\m�б��3� ����p;7j       ��7פ���   ȥ�oX��>��]��ʟ��l��%���q��ŁFv��]�S �I�Mk��;8k'�u=tr%v �1B�*e��       .��LI�;   ,�L�3}�؎��x���޻c� ���6�:L/e�U�cw������t��K5�_�� x��\�w�3       \hYSޮǮ   ȥ�4 %�����2~��_;���hj���s�?���)�c��a�����UYX�� x�4�-      �"4W$�3   r)�֩U�8�'��O&~� v	�p���ٛ/��������`Y3c�3���.}�ĊNT� �2�F5v      ����Ԑ;   �Ң��;#��l����Uo��lv�g�����|R�x�H���.����w����ZXi�N �ƕ՗��      � o��V�  �\JJ����3�)��
.����Y�Z
��E�; U����+�@��G�ZZk�N �!4��Ў�       �Ш��T  �ә)�cI��I��붼�mo��lf�����W��}��Ut�b��3�*���A�u���ǖ��`x �&��䭵�       �rI&+�b�   �%)tN���%�Kv^����{�;،�����^���L�GWH�Q�������?R��� �;������       r�[k��9   O�ʃbl�I�!)||�+~�c� �S��S�=W(�KI[b����L;f��W��	�_���;��hq� rǃB}I�63      �+4�cG   �%Yi vFn�4����&w��`�`�a�x
S�S�tU�^g&]:5��r1v
�jͶ�YR�b�  Ǖ՗$�b�       ȓЖ�j�+   r))HI!vF~��p�7�gb�=p^�<��=|�)|F��Dw�Ġ&�+�3���Ro�c��[� �BcY��%  F��
mI5I2�%%g��������5%�oX& �X������_�36��~�J��~;���6� ��)Q:8!{  �䝖B}!vF���y���|w�`�`px�?�����W%M�n�u3c�돝<��զ�{bY�l; 䒷�
�j�  �œ�[X6%K.���$�%�]Z���J�!IZ�aɃ�]V��jAi�^Ȫ#}�k���� ���?�T��N:�QV�'#&��+n�h�y93�4fҘLcrui�d#.3ٰ�c�o �+�)����   ȥP_�w�3�����y��+v
�0��i�\ajr�d�:vJ���%�,�A����ux~5v �Ix�V�-H� `ssi�d�.7�1�N(�{fvL�*�L��|���+�͝�� ��q���ƉN1Y{�y6i�)w�V���t��ɦ]���㱋 �-���
}�3   �ǃ�Փ�B��r�ɠ��nס�-@�c�8��}7�����n�����#2�Rȹ#k:�T�� x2���K��. `��VevD҃���a)��+U��!I/t��ֹV�T  ���+���&��R�m!hZ
�}���%]*�m�"� ��R��E%  ��֚��;#�<����<~��|��"���ӳ7����))������E��:�$���r�:����^�<�< @wH�2=(��ؑ�:li��=ܯ4yh�o~��� �l&w��`(�\li�d�\�,��]��̴M�+ ��e�~%}ñ3   rȕ�-H�;$��çn�l���1=
<l��oޚ��I�����J�T����XHb� O*�Ǘ�\c9" ��  ���q�C&�����w��3�yr�u���  ���\i�Y����g��]��v��s],�B�D ����o����   �㝖B}!vF�y��;w��Ǳ;�nŀ; Iss�ԿM�!�e�SzY1M�sۨ�E�� �:Y���˪59�
 y�YK��(�c�  zG��a�0�C�:`��{'�N�������� �yr��ŉ��;���.�.�|�d����T�� 8��ҁq1V  �xܤ}\W�gn��S�n�'1@��}�g�;cw���L;������W����Ѫ��,v
 �xP�6/9�k �qj����f�M3�F�?b  ��?�n�~N�G-�+�Y�@w���@�  ��	����b��Ss�ɠ��nס�-@�a�=o溽�n_��du$fҎ�UJ�S�'Ukvt�hU�,�N <%WV[��V� @�{�A��b�����j��  @���+M����9���g��/� �L����p5  ��BsU�Z����_�TW�z�K�eIppGO��y�h�W%����.���P_��I��[z�ز���S Ȼ�\���bg  �N��oX���ۿ��_m�������f�2  ����}���ҳ��?��Bx�����c� �����Ů   ��S[ܹY�����w����t��Ӧ���	�����m��h��I-�4���9�� �{�i*�cg  ��˾���%%�ݼ����?�&�� ��{�ܥ�`/�ܟ��?.�g�tI�. �UIߨ���.  �3y��Ш���
��y�w���;�n��;z��u�����$vG/��%�C�3�'ul����l�nࡣ�� )�N �K�����kf��e�/����Gbw  ����s���n��ܟ���0� ���%�K   r'�-HY+vF��7-�\s��;���'M���WX�E�`�^5�_���O!䐻���-�4b�  Ί+[[�B;v  &�U��%ٗ����N�>�� �f7��Ǌ޼*H?���+M�� ��+J�Fbg   �gm��|���~"k��-���N��R��]׾��<T�$=7vK��/�s눒�G�'�Ǘ�\�d) t�Ш���� ���ɒ2}݃��*��_��Wy  ��7���K�n~����ҳM^�� �AR�x�  ��w�� �W���K}~�͛�S`�=g����w����W�����6�B��}ȟv'�౪��N� �Y�v]�Q�� ��\���If_��|�oh�������  �,l{�\+�<d/���K���cw@WJ
J��Q  �3xP�zR{hΆ{�������;�<�Sz���W'������(��v]4�R��v�O�����%�;�� ��CGam^��N �o�<(ӗ/�kI��?�֯�N  �L�^3wi���d/q�J��� Ί���cg   �Nh�ɛ+�3�F��K�}��cw y�U�[fo�(5���-�[zQb���F�_.�Ng��֡c��d�@�pWV���n �&�ɒ��I��J��<��sGcG  ���kn�j��KB�%��?�L��] �O�d`�,�'  ����w�b�t�f�+����)@1���0{K:m'�v饱Sz��t�԰FʱS��YZk��W�� �MB�*��cg  �íᲯ*���랅��-��  ���^���������̮�gϕ�/��iIi�x�
  ���v]�Q���5��{I�|�ɻ�s8v�7��'L��?K>��W]41���J��qNT�:<�; p��R �N&%�&��f��o`��n�mN)  t�+�/�O^����J�Z�/`�;�^��Ȋ�  8S�6/�v쌮�!|i�o��7nm�n�wlz�o�w����4vK/�������iܥ�ͯj~�� �6:
k�y r�%}K�|�e��V�s��{+'�   6��W�8V���]����S�_!�;�9���	ɒ�!   �❖B}!vFw	�����bg y�M��F_���R��5�.��ҋFʺlz8vp�,��j��IQ �:��j�R��. ����%_0�}��/���?�	   g��z��r��=�ԤKb7�F�B���h�  ��	�%y�;��d
����w�?v��cS�ڳ��%����h����gF�$<f��v��G�j���) �u����� �%_P��QP��c�{b7   ?&^��j\+�W��jIC�� �BI*c�B9v  @�����d���jd!�f�����ش�����r��������6�B�u|ȏZ��CG���B� �:x��Ш�� ��f�w��Lw�Н�u�;	   ]`��t|�[�W~�\���w� 6K�LHƣ  �BcYޮ���.�'2���t���Nb�6����GB����J�^SH��6�r1��|_u����(��N �é���x��FrْI���n/�o�{0v   ����fB�W������4�	 �)+()sY  �i<([=)�e����W�'����W>�� �4ܱ�l�G�jk���ٱ[zMb�˷�h��;��պϯ��  ����ڼ:�K �X���>o�;O;|���v�*   lb�lw��J��J�OH��� �RҿE��  �BsU�bn�\��O/���=bz��t���w�\����E�Mkt�;�$�Kߛ_��r=v
 ����ó .�U�>oJ�6��o��9w<v   z��57l���:��Ƥ�R�^ �#)*c   ��l��Y쒮�����]�;�X�d�Mej�M���ӱ;zѶ-���{f�C\[�J�; �x��Ш�� �M�e�͒��mk~ۡ��5b7   g�x��+�ե���n�Y�gb7�ӱ��@�  �\��e:���;��w�C�pǦ1�����}M�x�^3>ԧK&�bg ��V'�б���N� �3ࡣ�6/n\��Ē��u���f����$�  ��2y��x��u&��W��� r)Q:�EJ��!   9�����,Ϲri�ڍ��=ߌ�l4����{�055�yIW�N�5��%m���4A�5�:tlY�,�N <��j|� ψ��f�l��}'M>Y���N   Η�k�pgG�k��j�_j�b�& �����,v  @�x���X��ѕ<��<;����}�5��)��bS���w���cw���RA���*Mx� �����{|E�YD	 �.ԫ�N=v t�5)�Kf����ٹ��A   ��6���J��s���f����	 ��QY�/v  @����ގ�ѕ<��-ܑ�V�c�'zS��z��^����=o��&�uјJ�$v
��K5YX�� 8�]Whp� �^�,�=f�gTX�������E   @,�^3���� ߣ�_)���M z�%J&$�]*  �#��T�/���^�λ��z�[cg �wt�m�p�D'˾.i[�^��i�����q�K�X��j3v
 �<��QX���m �<�*�]�양0����7��   8�ų\i�V~6��(�R����X�_I�  ���jR֊�ѥ,X��K'�z�_�.6��bn��7���~6vI��tjXc����q�,�бe�5�� 6we�y)tb� @.�4o��7%�>y��g���0   p�~d��������N纠ε&��n��ʸ�P��  ���j�3��k5�~�������)��ƀ;���u{]n{cw�����폝�Wout�hU�N�� 8OB�*��cg @�$'$}&M��:���t�,v   �����81��Zwͺ�W�4;	�&��l�   �
�%y�;�k���V��`���r<vp!�)
]i�u{(s���@cC}�tr(vz�J���-+; p�x��Ш�� ��XQ�ܑ�n9���[縧   �PfoI��|s����N惱� l>VTR��  �����3��{�o�����_lf���\sqr)��Iϋ��K��ڹuT�S���udaU�l; l�������@s5]vo�$�������Vc'   ����?�4k+?�{�z�<Tb7�,L��YR�  ���}���w��k�3��QUt��=7�[����%�b�+����&�SУܥ�ͯj~�_l`SqWV��B'v	 Đ��K�%�Z�O.~�\e   ��ȫo+zkO�ߛ�[�L�xfҒ����   ��"��#s������}�;��wt��7�ڂ�QR��W��i�QUJ|w�8:Y�Ǘ�Z�F �l8���X��/���,K���o?�   �S����MwJ�_0�/J~�x�
`���Y��!   ��v-vFwsoZֹ��]7~!v
p�������;Z*��.���-��L�13��J)v
zT�����U�;!v
 �<�v]���b =��[�}"K
[��� v   ���|퍻B��&){����{ t�D���dܚ   I
����b��3v4��/X�ܻ��O��kL��/$����䢉AM�E q,�Zz�����/� �ٜ�nnA� l^�Z�ܦ`�m���|w�    �����A鯺�M>�@w�B���h�  ��`��y����_r�+�/&6������%I���K&F*�h�`���c�5]\�� � \�ڂڱC �sYK�{�`��蓺u��	   ����������kC���ט��	@�%�1Y�;   ��~޸�O/���=�/&6	ܑ{�?�������pi,vK����cfD�,�C�Z\i�N \ ���9%�*��L���۷�]    ����M;�%����?�@NY�t`B��  8�w��O�:o[��7�� �>1!����oL�m�ݱSzE���m�*�I���v'�бe՚l����;M��b� 8_�I�-^�n^���;   @�L�v�ٝ�~I���E�{ ������   ����O�e�ם������)ܑk�{��ͥbw�41��6�J�;=����б�ڝ; p��LYm^r�� ��[Cf��>|�~���x�   xj���[��|����5f*�N�I�Y�#  @b�����/:y�{��x&pGnM��21}I⋾��cfD�����1��M=tbE�9�	 �YV[��V� X'��u:������w�v�������>gf�,�d&3	��e�E�Z��E�UB�~��o��V��ʖ���u�%��m?�E��@2@��E��~j]Z�X�Q ��9���}]�bo�@�Lf�u���/x�29ɼ��u��+
�5    Z�ș���%���A1k����*�c   b���!�WL�<o�맭[���I	M�Wv��g�#���[:�!C}��@��3Y���y� �2�9�ڜu ,Ԭ��>F��x����   �^֞��E
�Q:G
9� 6\��|W�u  @S`��Ҋ!�(ޖ�#q#1Z�hJ��n����k��)��u�U�� !D�d|V��U� �2�iM�T�� ��?���|��ى�>2k]   ���yɇW']�W�^�ú�Js�}�r>c  `�-�K/M?\��CXg ���;�����/�YRb��	r�sȠ����j=Ճ{fT�5�S  �-��)��% ���w�s�S7�k]   �3����S�Կ9J���{ ���[I��
  ������B��_S���/Y� �D+�ʡgo�m���I:κ�d�cTw��X��3�F��7 �	ByJ�Q�� �'Ⴂ����3}�˺!_�.    I:|�'rչ�פQov.<O|��=߳Z.���   ����5B����?�S���e�ʺMۮ��;�;:�sү�T.k��Q��葉YE~����e�ʴu <?�\����щ��m]    �3�!���8*��)Z� X&�+�[+9o]  `.T��e댶�oM�i�    IDAT��g���ɢup�pG��x�o8�&���p��~�]� ,��ݓ��;��A �)bh(�ĩz ��� J�����Go���)   ��r��O��噍J�;��k�= �����s��3   ����y�:���n/ޚ� �up pGSX�����j�H:ں�������� �4衽3�+׭S  +&*�/J��4�y9�JuU����c    `)�q��oSԫ��6#�����L�u  ��P�RlT�3�O�+
�_z�up pGS�t��R|�uG'����C���c�Uj��3�Z=�N ��P�Q����(w��P��ٛ��    ЖV�uŚ$T�षI�X� K�%J��%ǥ�  ��Ŵ�P*Xg�!b�����ɺx*�������~W.�&�>.�L�u�akԕ���l�����(�: ��b��P��� СbT�9w�sn���-;$�/�    :��[_,ޥ�3�bƺ��l�|�*�   siiRJ���'j���o���߭S��a�����]]=?����-��WY��\�u�\a��G&f'��R����u	�N�^9��WO�v�.�    �4x�����.)��)Y� X�;,�d�3   L��}���'���i���0�S��n�+E�κ�2ԧ��^����G
s*̔�S  �RQJk� :���s��yݐ�     �G�0�3ۯM1�yN�4� �3J���H  �t|�|b�o�l��l�CS�if֝{����o����z������3��i�C{g4W�[�  ��bm�:@�Qu'���?1~k��=    �
��������+��2I�u������3   L�FM�\��h_�]^�m�E��a�&�lܾ:��J:̺��e3^��F��[��MU��=�j=�N �iM�� �+J'��i�'�n�?h�    �h���#\��+Ʒ8�A� O����%Y�   S�|A
,�\.�PM�˿d]�2�abݦm��қ�;ڝwNG:���u
��l�����(�: `!�}/"�� ,������$�ţ7�K�9    �=;�[N�z�yR<κ�~$]Jz��+   L�FE�<e�Ѿ��o�������:�E�cŭ�x��D�����F44�c��6U��葉YEf��c��b�b���������;�X�    @;>c��»��ARb���|�*��^�   S�����쾆�={zǇ'�C��ƀ1V���k��s?�t�uK����F�3Іb���Uq��F �d�VR��Xg h'��ɹ����۳���s    �����'(T�/�s���$��x%}Ò�
  �\|?��b�;��]z��Xw���V���g}\r/��hw�]%�8Â�B�C{g45_�N ���p ���K���tm����/���U6C    �
+�s�D��;o8�	!�]�'ȩϺ�$EŐ�gs�!   f��(�˒��^.ι�z���^��k�l�Hlp�
�x����7$y�v�x��RW�?f,�z#�=�*W�� :[T:_�B�:@���sɧ'���uC�f    ���^���uo���V�Z� �|Ϡ\�  @�
�9�ڜuF�K�ӆ��K��:`�+�Wv�d�+�D�vw��*����@���Sݿ{Z�zj� 0*3���u���������_�C    hvѭ=s�Y!�?s.�ĺ�h�+�[+9� ��ҹq��}ٍ�����;�?�Agc�+bݦm����;�ݚ�12`��6S�����5�`� 05�r�:@�Qu��t^WLܜ��u    `�ϼ��r�=
�����LN>��:  ��VF���b�����7�[йpǲ=��SÿI�Z����l��[����ҙ���'{g"'��Št� En� � ��9��m���[�Z�     ��9W��wJz�VY� ����2=�   &bh(�OXgt�(������;й��������ѩ�[�N�Nig�I�:��n�`�g+zxbV̶ $)��� �c���::]Y��X�     ������]�;?��V�8d�t�(�[��Kb  ��w�+Ņ(wnq,�e�t&�x���m�vq�.��hw���iݚ^���=�%힜��  4�X+)T�O�Ԣ�S�ks}�z�����=    ��w��=39������:�����p�  �L1�+�
��!j�)���[/��u
:�X6ï�~|��ߓ��h˨�'���>�D����*�r� �Ͼ+ފ��u
������D����R�    ��������M1���1�9@��!�L�u  ���T�ҚuF��Q&-={��c[*V#�X���k��^`����t��C��x�����;���� �[T:_�B�:@�r���d|��/K.Z�     �@>�G�ͽ*�x�N��ږK�����  @'���By�:�sD��­���:��',��s�}�b�κ��>2�����!��=Ӛ+3� ��P�U�q����W�2����;�c     �k���/�
p.�ĺhG.�+߳�:  �@T:7!E.^)Az��إ�Zw�s0��%7���޹���ƺ����:��A���4DݿkZ�*�� ���iM�T�� �T\���+l��{�5    ��1���s��{�+$%�=@;�CrI�u  ���y��uF爮��~�p[�[�)��cɍ���o]Թ���9�Æ����?�z#���Ӫ��) �f�����H��\��}1Q�c��g�    h]���OIS] ;��|FI��/�  :IJ��%E뒎���ܯN��i��?�p��F6^s�sn̺��2ԧ��^���Z#��]S��^ <V(O+6�� �E��s�Ki�%S����    ���s�8&6*�Q�w���������   Xq�2�X/Ygt�({ql���d��X2������K�S�ӭ[�YOWF����8(�z��wO��p; ���zY��ak������2F}�8�غ    оF^~ٱ!M��69��u��|�\��  t�
��'D���[w��1"�%3z(��������͋	,^����]S���: �lB�t� ��#������/�F�����Ժ    �9V�}�ӳi���Z��c��$�Q�7,�@  @�IK�RZ���,�5�w/ߙ��u
�O6X�6^urt�w$6+,���9:�o��V�6���i5n <N�ك�:��s%���!��ll    XZ��}���݁�s]���|�  :KlTʓ�'J?	��ԩ�S�-hO�����~���oH���)�,��:��!y���3_����JC�N 4�P�S��Yg XY��\V]���p�:    ��6rf~}��PNoV9��u8��!���t  ����RhXgt sa,�u���8h#�}�s�*�vwԺUZ��m��5_���]�
��v ��Ŵ�P*Zg X!1j�ym�udz���     4��mt�P���{�{���J���8  �$�VR��Xgt��;
c����@��e�+��3�]��[�Y.������v �~Št� �Ժ���|����3��9�    h�^����^��H���������   X91*���K:Q�ug^0q���X���0���2�q�W��J�v�t�ak���X��1� x*�<��([g XV�,�3��.��9?a]    �b���_�.T�o��=�=@�r�}�r�� @���z�:�C�{2i��{n�u	��X�u��9;��d���W�t�ZN�c�n <�X�(T��3 ,�˒>�d����=�9     ,��3�G%N��8��uД|VIߐ  �"�u�R�:���/�򯵮@��I�r��O�j�燒�n�����Ç��x���R���w1� ؏�*�/�+ڀ��������̅��/��u     �e�YW�J#V�*��HJ�{�f���Y�  :GZ*Ji�:�c���y��-���@{`��2�iۇ�t�uG�;t�_#�s�h1� �@��!��6U�⩝?d�    �J9�cB���Aw��9��!���  @g�sk����]���.A�c�6��uI���n�v֕Mt��Cr|J� �jC��b� �_�6�X��� �T�k(q7�$w��M���u     V֜y��>����
1���J���x  �Q�ܸ��܊������s��;��-hm�: ��%�5b�}�:��p;�Tm��ln �_L��9� K#��_v]��,��od�    ��&wn�Aal�F��s�s�J�K ����   +��e{�#:ZT8e�M}ʺ���Y,�Ȧk79ſ��hw}=Ys�uZ�� &*�/J�n� E�o�Lr~����f�    @��p�
�^`�X��rI�:  `��T���uE��>I^3~�fM�h�〭=����#I�Y����T��80�z���R=�j ���ʌb�d�࠸�F��c�ۭK     hk�̿<F].���[ 3.QҷV\#  :AZ��ҪuFg�~:�t���o�����:|Oe�n_v��,��8`�F�}�n <�ب1��4��䕅���b�    ���ؙ��0��T��1��{ 1U��ZW   ���k� V7b��K�u
Z�8 �_u�I�{�uG'X���:-��ݿkJ��� ���Beں�"D����
�'�R�e�?X�     к\,�����G��ϓ�ǺXi�^RLk�   ��e�%�\���>w���-�hM�=��Ȧk��Y���U�]z����hi��oה�Նu
 ���b�b�`�4)��V�uŃw��     �Ď�pewQ�?��%NqȺX1.QҷVr��  ���s��9�H��t�p�拿a�������k_'�ʺ�{ؠz���hr!Dݿ{Z�u
 ��z���@Kq%�}6����S�5     ��5/��j�����-����\�W�g�u  ��
���q�
H��CQC���9c]���د����`��7I�ߺ�ݭ�����^�4����h��v ���ByJR�.�T�������|쒯T��N��    �*��Q-�{�='��.�aE�$'o�,�P�K�r>c]  �|�WL�RL�K�8��������6�c�F7m�ZҟZwt�c[��n^ ���(�d��) ����RZ�� �Qr;|�9��K    ���}�I��?,ų���hg.Q�7,9�s  ����-�C3pI�k'n����h<��I�����]��&6�/���n��+�?���,�< &����� �#�}ù�=����պ     <��[_]��S8ͺX..��ϭ��   XFQ�ܸ�u$E�I)wJq��[���qO":�)1ܾ"Fs�	hr��n ���9� O&�{��7Ƕ�&��     4�­[�Z˟�}�)�?d�,��(+6�  �3'�e6�Y8�5r�/J���xJ/�	�۸��t�uG'��e�n��:Ml|��=�%� @ˈ
�))��! ~Yt{��Nz}��?�w�     ��J��yW��n��\Q��vR�u��bZ���$ǌ  hS>Q�3{�,��=��f�r���M�47�P�8������K$��N��������:Mjj�����Xg  ZH��*��3 <�/+�*]�'����u     X�5/y�j��]��!{�{���2=�A�  �e���RZ����D���u=��/��u��x��s�����"�NНMt�ӆ�3Ф�+uݿkZ!F� @��iM�T�� �s�����
�\��u     X�g�J|�L1�Fܚ�6�{V�es�   �"��
�P5���\��i�p~ٺ͉w<ƺWm���臒�8��62�����x�Z�{�Tn ���OH1�. )�}�gܟMܜg�      mjhC�y�����_�n������  �e�ΎK
�!�E�����f���Ā;ct�5/�WXwt�l�u��r|
�Kꍠ{�T��/T ��ӊ6��F��ű���%     `e��������?w��b��U�7$FI  @;
�i�:ߩ7��|��;>��:��[�y�{��/f�}��2܎�IC�{�n ,HlTn�G��
�'��p;     �e��K�\�w'D��\ѺX�PW��YW   ,��Y'��\L˟[����Z���0^�}^�ό������S:A�N8bX��#���Qz`��f�5� @+�A���9���F篕��8����     �ֽ4?�H�a)�^Rb�,���e��3   �\:7.��:����Ή�ϲ�@sa���u�n{W���uG�X�:�Æ��3�d~2>��يu �Ť�I)�Zg )Fw���:��»�[     @sYsV��.��t.�ĺX0�(����.  XR�:�X�ƚf�3=o����Zw�y0������Y��!�Nq��k���Xg���,i��u ���ZI���h`����һ�c�ۭK     @s[{f��1ƏK�8�`!\�G>7h�  ��B�t~ܺO��ٴ����/x�:́�P=�\!��WL.�p;cz��p; `�bh(Tg�3�N3��+��x��     �@L���Rػ�Q��(W��TlT�e�  ���)鲮��a��k)EwC�;�ȫ�=݅�o��Nq�U���@�(U���)��S  -%*�/J�nt�U���e�˽w����u     hMg��v5�9����)k�<5/�7$�Y�  �G��*��x�g�9�㒫�;`�����k�.�7�K:E&�:�a9>y�To����`� h1�:�X��� :��)Qr�ޱK�.     �a���)i]����[���J���x	  h1*����Vs��Iw�{o|��v8�@:�Ȧk79ſ���$���:d��:M ���vM�Te�. `abZW(�3��眿Oޝ7q˖��[     @{Z�a��Q�����[��q]�����   K&��e�<��V�����s
��%��q��/u�\�+���[:��F�I�u��O�g5[�Yg  ZM�
�I)�,?#��<�?K_����k     @�*����˧��޺/K�y�����'���.9ψ	  h�3���b8�ow�|�����)���5�i����a�N���KO_��:M`�dI�'�3  -(Tf�%��]Ey��ȾsⶋvY�     ��2x��L\�c
�U�{|4#�(���  @;�J�&��Z���8_Vw�Y�x?K�:�h��+G���#�i����������nj�����Xg  ZPlT�mo�����˼c|��_�n     �m茭/s.~Z
ϰn~������3   ��Z��|��{�su�&N"t ��v��2�����I�r�w�R����  ��*��Z���K.�x�Ng�     4��[n+�}��(^����~QlTk� ���9�<��x�P�ދ�3`���s�9!����2�-�d���΀�FtϣS��9L X�P�RlT�3�v�:�>_w=��qW#     ���~��#W�<��&I�u�����K��!   -���B�:���%���6Ϻ+��3�iۘ�3�;:ͱ��Qo7g
:���5S�Yg  ZP��*��@ۈ������7�k�     p �6�礫��,�@��%}Ò��%   %T�ks�x*>���a�N��o�[�`���AF7]�21ܾ⺳	��nWq��v ��T�2k]��(��K��o��:��     �������\=G.��(W��S�ʌu  �As����8i����Yg`e���S�0��w9�d��i���`�u�L�W��^�  '-��CR�A��!�s�҅7}�#     ����p�H=�>.��YhS�{@���:  ࠤ�)���E�p=ϛ��=߱N��`��C�n��O��6�Nt�ӆԝM�3`�RKuJC�N ��P�W�2���_]&����     ���q��%w�s:պ�����%Y�  �E���2w_w��+': S�`�9�p��W$�o��i�z�lo�g��    IDAT�P!Dݿ{Z�F�N ����+��@ˊrS���8��-��_�˺     `�������׾���G��(���z��Йb�&��I���  �59�(�K�8 a$7�H�w�k�%X~\Y�|O�bɭ���Dkx�ԩ~:>�J�a� hIQ�2#�@��sA�9��g��$     о��0�s�vɝ,�,^*�BL��Y�  Z�O$ύ4-#T/\�{�8�:ˏ#�mn�ƫ�]r�8��✓N:r��ǬӌO��ha�: ТBe����"��]�ɱ�ߴn     �0r�egD�W���nA�q��]}�   �j��Y�(��V������,6����2��&�{�n�@�vn ,Nl�n���%N�U��    @'�yɭ}:Q.�Pr�hĊ��Y�F�:  `Q|�˖��Y��wYg`y1}��F6^s�s�;� ���G4<�|�$Q?~��z��a �E�A�|A��u	�B�-J�\���G�K      ����<2q��)��a݂�%}ÒcD  ��t� ��uXR�I���[�w�u	�Om��L��ͬ�uY'`��t|��v �����������(����ֳn     x���?Tؑ��}�):�����*-O[W   ,�˲̶���kۭ+�|~nS#�9C.�غ�S��d�����$��eM�W�3  -*�ˊ��u���kH����;�8���:     �ٍ��rCR������{�,���P���   X0��N�B�ڋ���o����p�X������t�uJ�:t�_#�s�X!�j]�>:��K  -)���:�� ���k��������K      Z����ω>nw��Y����ܐ\�[� @kI�R�[g`��SI��	�7��n�,-VL����F_�p��U�<�w�4D=�w��v ����i1��G���%�*�m~>��      �W�-���sݳ��y��{��BeJ
�u  ���Ž��cij�u����Qo�|O�T���#�[:U�;��[c�����M�W�3  -*�����@s�x��2�3�i{     �%����.�6�Y�-hc>��wXr��  ��CCa~�:��z^=����u	�Omft����#��l��>�[�k��0>]֣�9� @���`\��5 �/��O���O�m�ٺ     �����uc⧝�!�-hO.�#���   8`����X(����������u
�������O����n���:+�TmhW��v �bE��n~It�̕����3�     ���wl��gKϐ�ՒR���ب(T�^  ���N�b�t��\��:K��mdtӶ�Jz�uG'�&^'9l��eB�=�N�R� `qBuV�6o�4�m��G�c�}Ϻ     �m�?��p��N�nA��A��  @K�i]�T�����$��ޛ�w�u�m�Ѝۏh��ǒx"4�f�GG�Xg`�=R���t�: ТbZS(q#�s~&����s땒�Z      K�]Cs����>��w�XB^�oH�g�C   �R:?!���"����'�;�Ϊu����h��b���@��:�l�\c� �x1*���+����#�:����O3�     �n�׊c�-N�Ӣ�7�s�N�ByJ��:  �)q�L늡~�df��<6�����l;E��',�;��ae~�*Q?~��z��. ��	�i�:��(7᝿xb���-      x2ѭ=��?
!�s�ںm"�RһF��  �fӺB�`��E��ה�������к��$npi�B�,��vgnos��2� X�ب2�HrQ7t��D��     ���;�l������A�Hk
��
  ��rIVr�u����Ci�uGb[���k~�9����֭���5}�X&�ي~:>k� hU1(����Ut�������-[��:      7�!����	'[������.�_  �+Tf�%���������Zw`qX7��s�n�>�.�,�Z#��u �������dQ�!4r�1�     к
c���g��r��-h}�:�بZg   <)��N�AJk�O��x�u��-ld�ug:����tґk��D���vMi�\��  ��X/+T��3 Q���Ͼun�n     ��ސ���x�S<Ժ�������u  ��Jg�%�̮�ez��p�o���±��eE�b`{{���u1�ަƧ�� /�
�Y�
�B*��z�W��p;     @�)��oL����JrL�`��Bi�P @�rr�.��F�uk_�߶���1�ۢ֝{�c�c݁}����u�X���b�N ����4)�5�`�����a���b]     ��7�!�;�q�\<ƺ-*�RһF��  �fÍ�m�e\8|�d]�V6ݶ6����31ƭ�����LkG��2� X�P+1܎��j���>z*��      ��0��߹�էH�jI�uZPZS(38  ���t['`)��3����u��-hݦk�宷��>�9=�r|��Ja����g�3  -*�u�RQ��1~���X�-�-�      �93�[!�ϲ��Ჽ�=��3   #�/H���-�'e��2~���Z������������K�;�s�=���L���0g� hYQ�2#����kH��B�?��v      ����g�ܯ�ܱ@�^R��[g   <[��DHs1V�[g��1��bF7n;_N���ϭ_ӧukz�3���3����u �E�ʌb�d�,����8>v���[      �|�n���cL?�6w,�����Xg   H����XN.���������%xjlpo!#�����;�X}=Y�,��l��v ���F��v���mm/�g3�     �'31��kls�b�ʴb�f�   IrIVr�ڶ�(��O�{�G��K���Ե��I���9���u�H���ȕw �E�A�2m],3�#e�
c�w�<�0     `����ra,�N���(�{�{�*�BeJ14�C   $I.�m��%C���L����Sc��E���k%w�u+ו���:K���i��  ��P��"K�Ц~���Я�
��e�     ��2�3�u��cAbP(MJ��o �=�0��Vj�?~�ǎ�����z�E4��$�ʺ����G�]̕뚚�Zg  ZT��e�`Y���c�M�^�]�      ���o8�,�k7\������c����b��4��wh���   F�mpw��u
��S��Z�JI/�n��c�{X���H�m�x�\w�:K F��Y� @�
���@��r�����~m�6��     �4&�6-7��9��控�J�Sb�  �rNJ�l'�Q������+�;��poI��I9�<^����`�TI�:��  ��V�%qE*ڍ�۹䷊;��;�׭k      �^���rag��N�����A�K�
��
  ���mqG��J�O����X���1���־r�!Q�-�x��;�t%�8H�F�ީ�u �E�ڼ�֬3�%�s�3ewja����     @{����������Xэ����Bu�:  t0��Ph9W�{�u������n��)�ͺ�ן���C�3p��=���� ���i]�T߹�]D%?��wn�'�      t��g�ω!n��z�4/߳Z.���   *��bj����J�o��=7�����ܛء�!�?����ue�p���� )*Tf�p;�D��_��3n     ��������}婢'*3���  6\��:K-�=iy���x<ܛXçI�^�&���Z'� ��H�+�  �*�R�[g K���$���3���X~ƺ      �mz������I�Q���A3�
�)Ŕw�  `幄q�v���k_�[w�poR����#�F�<��n6�����%��: Ђb��X/Yg K�ݒI���[.��u	      ��
c��rI��Q���ByR14�C  @�a�{��R�z�1��Ca��I���,��T❺��u���*[g  ZQ
�i�
� ���
c[��s{~�u      �D
�\�Hq,�R�?�4o݃&�BiR
�u	  �$�K�Ÿ�(���OgJ����1�ބF��~t�{�u�\O�I��]�9��3  -(Tf���r�2���eN����%      ���عe���N����nA�������  �����]��z���Of݁}poF1�,�	�&����U��55W��  ��X/+6*��"�r�?�0��ES;/~Ⱥ      X��.���\� :�5�լ{�DBCiiRb�  X!.À{ۊi�+W>n��}�u k�U��p�poj��kdu�:�p�S��ԭ3  �&�J�����������7_�C�      �`�l��� �EI'X���$]Jrk$�  Xf1(��k]���|�����+��W�N��&�2!/�ۛ^O�[��\��v �"D��i1܎�J��!7���     �.��.�^��Y��Jr���>iMiyJ�� �2s^�Y�
,�\�6�99i�@Y���?��	G�+Ï����_Uo�� �0�:�X��� $:����Tܹ埬[      ��v�ֳc�����-h.��ϭ��   m�9�v��2}0q���ƺ��1��DR.?���x�p{�.3� X���y(E�q�})��L��     ��&ƶ��;5*�ͺ�!6�
��  ��\�e��ec���l��ۺ��%��g�Uۏ�>n[��^�+��U=�X�4D=�wF���  �ByR��B˘�1�Ӊ[�V��b      ���=wΕ��}���nI�#)k�c�.Ir�  ��p�+�J�XN1��eU-����[�t*�P7�$I/?����Ź�V�w��40� X�P��B�:8 Q��i���ߺ��-      ����[�;�N�ܷ�[`/��j��  �]9'%��lw�Q����k�[wt*����ۏ��j���,���.[g  ZLlT������jQ���s�[S����      ,M���]ػ�ף����&.Vgy�  ��K�-���F_�L_n�ѩ�u �u��}.Jo����9r�*�u[g� =R�c� �0!UZ*H1X� ���=J���m�oY�       �f���o�Q���n�-����Xg  �6ӺB�`����4����x�X�t6�[��G��8p]6���Z#�0�p; `!���4��hv1�_��[u*��      �ߙ�z��i�%7X��V(O+�5�  �f\�#� �I�W?e�щ�t�.s���u\w��V�{r^1ZW  ZI��K��F�r�蒍ű�[��|N�      �1uc~jb�Mr����u�D�ҔbZ�  m�II�:+ ���}��ϱ��4�z�5O���;p��xg��P�����Xg  ZHLk��9��IE�o�_��=Jһ�����Tu�=�If&٨���o��!@4�8	!r[n��LWѳ�+��@�U�(A&�=D����芈@��LwU������}���	�LwW��.��99�9��;��Lwէ����ק��ػ      &���/������-�Z�Tx�  �J��	�&���W��1�M���Q9eo���pCd���Ccv���v ������xV�����=c�p�.�      `���bm�ާY��.)z���%�f��;  �Pb�<.�螹����zw�NQ;9������I[�[p�v�آǞv�wE�H��Wk� ',�dO���1�;�M\U?r��x�       �b��מ�,�����n��PR�}�BV�.  �Β�ʬw6K61'v~�a�;ep��I9�7�q�Й,�%3�� X�[��1��-y��D��      @o��L͔&'Д��wXTj�K�C�  `�B&e\q)�SN�k�3����NS̿$i�w��Swj��m�xEL����J,� '�R�ԨKJ�)�7j�~�:3�[�!      ���{���6�;d�7��M(���)+y�  �!��K��靁���c�����ڻ�SF�=��ĸ}(q�}��-�� N�)�Ÿ��,|Z�ē�      ��:=uS&=M>�݂MfQ�Y�;  ؐP��X�bk�i^�1X�n��ܰO
?�݁��`�>�b2ՖZ� �!���Rʽ3��B�tc}WxR�����      ���t�����'*�~߻�̢bk^2��  �ub�>~��U�_�k��1����&���A��݁�)�x4� �-��� �Ί���0J�ߪG�;�      ��c���!�ŧ^xݭ��
i�w6I*��*m�#�� ��	Yy�{>07>,��n�m�.�Ne|g���^�ۻ2�g�;�~%�d��T�z; �DXRj/zW �$��7��      ��v������K��[��R���;  X�P��N�&��{������Q�Zwe[�?m���O��)�
<��fGy�� �G[��@�A-do��Ω�T���      �u��~�6{��,do�/(�F�  `�J��tI�Yy�w�(c��I�<��-K��_�t�w�g�DI���N������Zi�� ���Yg�;c/�'�~�vt��%       ��*�Mf����-�$�I����  ����+5k��tA��ݗ�~�u�]2���I�v�_&��Cm�̗ˠju�� �Ge1�uV�30�����1��v      `8T�+�$O�e�݂M���y�̻  �P*�{��ȔR�m:�R�.E,v7Á�$��;S.��2���-� �����Z�ċ�p-do��~�ح�Y�       'n�h��ڮ�=�B�v)$�lF�  `M���qGVt�ܻ{�˽;F��x�-��;�1{woӷ���;��_�)�� ��ւ�h{g`L��=Y��d���'�[       l̾�?/Y�{��y�`�����d1�  �&�e9�Z�Q(M�7��=�_��n%���;&�w�
l\9��e՗ی� �(u���Ɣݚ��1n      F�����!m�!)��l��Ql�X  ��B6� '���l��;F1�Ӯx�s��w6�Swj��m�x��}��N�3  �bW�9/^x�f3���tp~��ۼ[       ����Nm|�Wd���J�9�Pުl�n1�  �b�Ԭyg�K�X,N>�;?�y�Q�I�>3�7y7�7��T�r�˸ ��,)�Ÿ���.����      ����X����Y�BY���AY��;  xD!+�Í1�w�W����>�w�;�!�l��F�����.��  ,�%�P�lᖴ%���t�/�K       �_���ǂM>���w�,v� ������+�)v�+o��1*��QP������ɣ�[]� ��J�)v�30^�)��6S�h�Õ�       ����_��>Sy�)�N
ɻ}��  <�Pb�>�R��Ӛ��;cT0p��W��$��wz���`�]h�x�  �,ve����p_�Jϩ�T���w(      �X
V��Le�|�)T�k�G��؜oX �o�wt����������Ĕ�,�E��_.�"/�V�� x��Z��'f�����G�>�      �������\~��ɻ}��-F�  ��Bi�;ެت��A�Q�b�N;p�w�e��-.���RK�
  ��[�E����kg��=��_9�      `p,>����gIٍ�xcsT1r  2�_���o<ƻc�1p���K�Y#&c�>b2ՖZ� ��:+R�zg`�4����L�jU*ɻ      � ��o浙��!�^(�%��	#w  ��B�2��cϊ-Y�5�1���طx�)�^�݁�c�>f���  dEG�mxg`,d�`����#��z�       |�#�?4��J�w��I�*6�q  H��;$)�x��7|�w�0c��c]uV���^Lܽ�ERu��� �IQ���]��g!���v���+wy�       ���g��<�	
���[�')Wl�3r  RV�.�@���a�b�����mm6[_�t�wz)�    IDATs�w�ػ����w �72�F]J�wF���J?];r�7�       l���}����
��݂>�&TھG
ܛ `\Y��HV�rԶ=�_����w�0�;�j��/�����v�"��̸ �@��̸}�}&d[���      @/T��n�D��p�w��K�   +{`PXQ
ݕ�3��^�T2�^�<��ݽ��yW  ��-Y����(�?.�gU����       ��v��?X���0�݂>`� �XY�;�b������zw#�=���N{�L�ٻ��w_�v��F�; 0@,�J�%��(S�Z(��6=��n}Cû      ������3��J��J��=�1F�  ���I���,f����:0p�����	,�ݘIwWW�3  �ĒRkA��@?��2�~�>=��       �.Xmf�R��BS�zנ�R�ج3r `���:�݋N;p�xw��z`߁��t)<ջEե����; 00����٠B�wab��3���;      ���=�KK�d
�ϻ=�
F�  ����]�Ab1��!�a���B\oqf\��PĤم�w `�����r��Y�jM�S��/��      `�,��yR+<U!{�wz,����8� ����;��\�����w�0�h��x����ߐ�[�_����0v�:��f��� �U�ېu�=��+j�So՝�qB      ���;o+Z����[���ǂ�GT�nB����(��(nQ 0�,�R�x��e�����O��wɰ���Bx��uyp�|���� ����+�,{g`Ԙ�H��Z���}�       ���t�=�P�QS����ĢR�.c� ���mx�w�8������1,�*ڀ�ܰO�yw`s���}�1�k�� ���T(��30bL٭Eiۓ积�W�       x�ٙC=�����nAYRj�3r `���X.:�k�+��Ha�5��zw`s0o�<���c��  KJ�yI����������y�G�<�       �ح�����=�B�v)�B��8�އ]�  �/��;���O�r����1��ә�߰E���������Xht4����  Sl-H�C0"L�j�.��T���7w       �͗��t�!�^$<{d��^t�C  @?0p����̊�/yw�봸�t��ӽ;�y����n�t�ܲw `@����^�����*�U����       kU�>��Hg���-�Sj-�r� 0z����Y��l�7�'�A�W�:�^�݀�UD���Of�]�K�\� HJ�Y�������4k�ٙ�_�.      ������R�����-�Sj/�  ���x$VlQ��F�AǗ�:�v��ϲ`��������N��;�xg��{��.4�3  ��R{�;�!����g*S�!       �;N9��J�]#�GDزK���  ��JͺwY6ќؾ����|��wʠ��uH�~޻�//���/K�.�v �$Ɋ�v�),�L�g�      `���T��R�
I��5��,+uV�3   �R�=�6^�1���Ѿ���t�w6_���	#�ݍ�kv�; 0 ,�J���������G�;�       �2w���rv�)��wzú+J>�  ���E�=n��1���Q(�׊_����2p�"&}�آb2� �3K�Rk^&`�,�H��Y�3��       �V=\����ؤ?�nAoX����H  Í�N@�w�;�?�1�����|�;N����UI;�[��&J���zg�3�K�-h��{�  �Y*����a2lH4eo��T��C       `�Y8�k�G����d$��6e�N�8 >Vt��Y�&�;�}����/k{�.����ĖW�q���cR^$��
�v ��"�vl���J�0n      0��է+oTVz����k�qV��Z��,  È?�qb,�{��՗xw"�'��JYA?�_+mٽp�|C�%^S��gI�Yg܎���,������a�       �V;2��a�W�[�qV����H  Ã?��)uߠJ�=���r���?�RI���V�;a��-�tl�� �Ƹ=`!;&[O�N���-       0(����D̞h��ڻ=;��y�x�<  C��;����w���΋�;��~޻���oHm��{j+�  o���R*�K0�L!{[}z�yՏ�m�;       ͱ[+���{�)���nA���{+�� 
Ɵ�XSjw~ѻb��a���w��̲Oyw`0�y��ڱu�;c�,4:�kv������q{�]�����e��9�~�       �\p�Jz{��aJʶ�Q���%  ����,ozg`�d�v��]�W�%���' ��j���r�;a�ԗی� ����>��ٌ�      ��է���&�3��w6ȢR�.��� �@�;�,�:�7{W��+o�+�
���FG1��>Qs�-}un�q; �;��ذ�S*M<�~���z�       ������d�IR��l�%�漬�z�  ��a)z'`Y�w�e��>�A���Q�_%i�wGL��b�;c(�o�ڊw ��%�f�q;�/dأSή�r�׼S       `X-��i���Q�lTRj��r�@ �@2�X�!/��;cPv�����z���z�`�����}̩*e|	=3������0 c/E�ּ�
��h��Z��Ly�       ��p���V��A�za�.e�;�3  ���W�yW`HYV�f��|G���o\p�C�b1n�C��tl��1��"��.0n ��ۛu��X+Yi���      �ׂ�g*S*e/U�x|���βR�'� 0(��6 �bR���;�G`���n���[li��{g�F;��_�W�ͯ �����<v��E�)s���w       ���-�߳�=[
�y�`c����^��   G �a���{�o�������a�~�=�ҹ�lw�-)&��ե��x��S  �,�۱�_�){r}��Y�       u����6������{�`c,o*�$�a  ��%�ؠ���R�����?���I
�ly�t�E�1�1�+ǖ���l|  �Y*���۱>!{Om�㞽��J�;       �E�c�r�]���t�w6Ɗ�bs^�y �#.����ϪR�7�p���8yrr�ݒvx�`8��}R�=m�}E-4:�ZuEW� �,�J�y��sk-��T?R���!       0�N���7��/K6�c���M��}��� �f�+sD�w��؇^��/|'��LN�L�۱Kͮ�2�46��W/�/�+ǖ� $1n�X����<��       �6=�����X!ky�`R�بɸ  ��J�q;z�;��yWxb��M,��OyW`�,6:���u���*%��bK�����F�; 0 ,v���۱v&ݕ�윹���       ���-S�R�#��^�l�E��,��%  ���E/Y̟���;��ᅁ������%}�w�S�[����k~e���fR}����]�=��1�T xtV��q;�*�c)dO��>���%       ��>�V�Y2��0���{׻ ��`��;zȒR����^�?H�����Lw�.�{����}�k���ܲ��" ��h+��%��'�Q�>P�Ξ����       xh�+w�������-؈�:r/��!  �<+�Pz�ȯ��K�y�w���w� 9��M�I�n��@^$՗��I�&���U�j�m�5���R[Ed� x ��J�E1n����֧+?����c        ������n���}�_n���{�~��Cyҹ �eI�Y����I��l~���]�نgq�	�,�J���c��m���y�qς�W:��6;��[ֿ�U�=�usvg �o�:n_�v�M�
�tU}��F�       �Z�OWި��3fʽk�~�]Qj/��x  �=���oR��z�M���1��έ�w���$��N�hʋ��FGե�Z�B�L�R�R\���Bե��V]��BK�n��� ����Yg�;��¬�tAmfj�;       �>��?���|��X���ݻ�r)E��)��  %�7�Txg`Yܹ��}��[?흲��N��}W��@0}л�gۖ��o���ɒ�o)k�DYY�F�fR�[����h�Zi�*b���/ ��I�Yw�;C'�lQ.=w���/{�        6n�y����E���n��&U�v�2�  FB\���-�#�&��z�5����L܏���W�g{w ��e���rI�r��R�r)�dy�?C
A�BP���L1��UĤ"&�ER;/�ɣ:ݨd�g �]j/��w�N�eK9\q��
��       �����މ��4Ȟ�݂%e��(de�  ��ŮR�����s��fo����.�,�%��ߝY�9��  � ��Z�-��k3׾V
|�       Fс���O�^蝂��m'+�&�K  Z�f���~�����Iʔ�Z��  �L����k-�__���j��       0�n�tkӕ�Jo�B���:YRj���w	  C�
�E��ؽ�K޽߻c������/}�V�^��  0P,)����.�P	Me�ק��w	       `sԦ�~U^",���)�d].� �VVt%�~�`�DJK����,c?po���K:ջ  ``XRl�K��]��rL)<�v���x�        6W�h��!��3��݂�K�%���w  C��w�H��W�R���X�M>�^�   00RTlԤ�{�`�X�\����*�       �Q�9�Y��4I_�n��Y�Tj-H2�  �%Y�Cl��b񘽟�q�w�f���+���
z�w  � ��+6�E���Tl;k�h�N�       ����[�0��O����n��Y�^}گ%�  Z�[�Ca�\&���zWl���+駼   �]��<�v�M(�~�����M��)       ��p��[�v��L)�c�l@�FJ�w �ñ����|��~�;���o%� /���A�w%m�n  �dyK��(>U�5�Jv�v������8�       x��;o+Zw|��m��W'�S�{�N�dE[�4����� ��dEW�7�30�,KY�m}���.駱���e��N��   ���X����JW�>v��x�        Y������k̔{�`�,)5�eEǻ �������'��ez�M��4�w3�ܻ  �Sj/�:��.s��t?�       ���ԻK��|)[�n�z%�ּRg�; ��`��"��K�}{g�»���r�~���~Igyw   �0�ւ,oz�`����r����k��;       0\�f�f2�sM����uW��K��� �qg��c 䝟�N觱�'��   .,)6�eEۻC%�S�<qα#o��w	       `8��\�ϊgI�3�-X?˛��yɒw
  >Rds��`��}�%�����2v�3ϿaK0�I�  �M��b�.Ůw	�JvxW+�=��_:�]       n�[��j��1���݂�]�f]�
�  6]꬈��` XR�#{�}��˻J�J:ջ  `3Y*V��Ј5!���]|�m>~       艅W��>K�����
�f]�a% ��TȊ�w�u)^q��7l��臲w�f3�^���g  ������Z�ģ"q��B����Ե��N       ��O�f^����'�����%�漲�')Ll� �דּ� <P��Y�,.���^����;��   �źM�ּ��D�B7��ק���n       ��`���7&e?')z�`�L����Y� ��,沂��c ��+��a��)�^�1�{  �+���:K�&�-J�ys�S��N       �����;C�]*��݂��nC�9/�y�  ������R���/~�c�;zm|���V�Az�w  @ߙ)�dyӻC��.M���ʭ�-       ��R=R�hI�7��݂��f]J� ��[Rʽ3��f1˭3rW��f�~ھ�H:û  ��,)6�<k�}>Y8g���O{�        ���̡���֧��[�)_}�*2 �KJ�e�
����U���&|��fI
z�w  @?Y�5>5�51e�謅��;�[        �:��/Lj�YR�G�l�E%2 FD�H��3�G��o���;���Kc1p�������   �bE[�Y��G>�ąP���N=k�Õ�        $龙��e��LS�g�-�Sj-(u�!  ��Ů,ozg '�;�W{W��X�C*�DRٻ  ���Tj-H2���{�Ӈ��͕�w        �h��J}���W���݂���2�c ���R{ɻ8a��sϸ���2�,؋�   zϔڋJ~���t�:}�+����       ��t��6]y�I�{�`c�h+6�%K�)  ���]�R���`�D�U�wG����}���<�,��  ����ب��w	����L�+�3S�        
����Pz�XG��Ul�d1�. �QY�e݆w�fV��{7������ �H��+6jR�@�I#˲K�f*��       �Z�OO�]��2S�z�`,*5벼�] ��3Sj-xW ���=��_�wF/�����/}�VI/��   ��[Jͺd�;C����G�ӕ[�[        X��-��+g�IZ�n�F�R{A��$ɼc  �&���&C,)���]�#=po��K:ٻ  `�L����^/�a-L�n)�H}��w�-        l��_�X(g�J:朂���؜�,y�  �,oɊ�w�!����	遻��Ļ  `�,)6�e�����Vg�g*��.       ���+���&�1˾�݂�]�FM�
�  d�Pj����=uou�|ف���x���xw   l��\�Q�b�;C�,�۸Eg�����       @/��r������쟽[�A�uY��. �33�֢$�,��`yg�����=��%��;   ���Rs^�蝂!c!ݾ�g/|����       @?��2kҹRv�w6*)��:<� �#���{g ����i�w�F���]�^�   �>��YVj/�Oc���ԟ.���׵�K        ��Lei�N9O�>�݂���RkA2�N ���Y�I"=Vl-uxgl�H�O{�;�����   X3K��yY��]��cR魵�k_�J�OF        ��3WwjO�e!��z�`�h+6k�Tx�  ƀmY�'�`D��E�	1�w��%�   ke��بI�띂�-�^_����;       �MW������4e�y��R�ԨsM �Ws�֒w�7�����m��5r��;��I�.��   X��m(5�E�3�e��OO�û        O��ʔ�����N�^Rj-(u�� ��Z���#�RV�+�#7p�ͪϗt�w  �	��؜�u��K0��V�J�V~׻       �AP�>�k�e���»gݕ���w
 `T�)�8@���R����5r�`�  `�X�5)v�S0��%������G�K        $sG�~;d�)4�[�qV��u)1D l�)�楔{� �#���w����X������"�<�  �GcݦR��'��^s!�Ϫ��s�        Qu��o�e����K�b�&+��% ��eJ�E)�g	�IRj�^�]�#5p���&�;   �����:K�x�"���V6�#�#�ʻ       �AV;:��L�\Y��nAXRjՕ:+�% �!�ZK���l�B����V#5p�t�w   �ñx�e��w
�U�nOa��#��;       �a07s�?�,�c�W�[��]Ql�K��S  C"���j`|������i�k52��t�;�]���   %uJͺ�
�)ٿ�=}a�^�       `�ӕ/H��e�s�-��Ql�d1�.	��:    IDAT ��^��M���)��Cw@|d]%i�N� �gI�9/�,K2�)��7���#�n��U        ֡>S��;Α�Oy��G,*5�J݆w	 `@1nV���R���P�>���n   �FV�U)v�S0�,��'�ó�?��E�        ����J5L4�)e�y��WL�YVj-H��c  �q;�u��{�e�9�k1�}/x�K�~�   I��R{�Ұq��~����;o���S        Տ�my�N9�BvĻ�cE[�Y���; 0 R{�q;�`E�B��{H�*�   I�T��x�Jؠ�߮�z�*>%       @�1su���q�
�݂J�R�&�[�%  7��Z��ࡤt�|��q���^�dRx�w  �u�J���r�����t�R0�        F�͗��L兦�7�S�K��^Tj/J��, 0V����q;�P,��N-��#�'j��}v��$}�w  c���J�%I�P�1Yv�6S��;       ���>Sy�I�{���,o)6�R��) ��`i�����.Z(�z7����[Wy7  ��eyK�Q�$�BT�~�v����!        ����u�L�u�豔+6k���� `��x�CM�w	0�,���Jٻ�D����/}�V�]��  Ɛ%�����&�;E��U����)        ���Le*��7����KJ�y�6Ob�Qd1?>n/�S��`�)�O��,�1��f�}����;  �x��j�m��S'+�������w
        �l~���C(�FR�nAoY�Tl�s�
 F�m�f]2���"����'b����  `�p�=��B(������K        �T�>��,�_(Sǻ=�ǏX� ��u�J��t`킊���K��fh�g<���t�w  \mG�eK!Vg�{�        ����>�A�KW�o�KJ�y���E�02���Rg�;Z���}񮳽;����m鹒vzw  ���v�I5%=�zd��-        ���n��S˲�daŻ�gyS�Q���; p�,)6�ey˻z)�^���h�v�̮�n   ����
W��ss���h�c���        �>=�g�ҏ�4�݂>H�R��P ���\�Q�b�;���;�����{�o�ʶv�I���  F��b����`�3髥�mϚ����n        'f���Rv4��z��?By���'Iaho��Ȳ����y� #$�<���}�u��]�p��l[�"1n  �f��YQ�S�����ɲg0n       `�T�\�)��3�p�w�Ê�b�&�=B  ��^Rj/�q;�k��ڗ{W<������  `�X�QlTe�����6�s�V��        k7��lb�9&}ջ}bQ�Y�J0  K�b�.˛�)��
E~�w�#	�ku�U7�T���$m�n  # E�β�h{�`de�͂�=7]�        C��;�������-�lB�m'KYɻ Ǝ���6J�)���,������_{�w�C��n�R1n  fJ��ի���7�g�Q�d�       �h8v��_��tI�{���R�ب�r�G�Mc��^Rj/�q;�R(5��+��܃���  `�Y쮾 �]�D���OOh�Y�n��z�        �ީ�T�Vi�R�y��SRj/(�%�=E �'K�b�.˛�)�XIJ��nx8�;`-v��]{��OҤw  B)*u��؎����S����?��E�        ���W�;��'B��nA�eee[w+�&�K `�nC��@!�"��߲��_Q�Ny����>Y�Kĸ  ��%�βb�ʸ}g!����g3n       `�-�T��l��i��Y*��u�nC0�G,�^m�,��['K�����e����'�  �01�ncu�΋M��}r���~|�ʊw
        ��Õ�B8�L�݂~3YgY�9/K�w 5�[�����)��K1]���P�w���s��!Ί�  �X�Vj/K�S0&���Oj���y[��        0f�^��])�>���n�f
[v*��� �ŒR{IV�:00By��L{u[e�>�74�'��\1n  ��b�ج+��ce����       OՏ�m���y��/�[��~�]��$�DX�VlT��Ɗ�{�l�i��]�.�N �U&YZ�+EY*d1�_�X�!֒d��K�RkA�Y�V�T!�n��|�%��¿x        ����*+�w�t��}»�$v�5Y��.��eiu��ZX�R8)�^���`�;�D�񼛶��$���,�R\��������7�MV�$)d
Yi��L!d�����ߏ��81)*u�_4�%�\A�U���R�p         I:����U�HP�q�l�Pުl�IǷ  I����Yf��0�������FC�����/��C� F���c��ו��a��%)+����A|I!+Ka(~��ϒRg�a;��?�>%\Ÿ        <ؙ�߰�jf�y�`�Lٖ]
ۼK ���B��$E���l�)�����w{�ܯ�pB�]�n����bWVt�>f��T,J1������4~�P(��8��v��}��d��q;        x(w�\�с��OY	J�{�`�XRj/Jy[��'�>� Ɖ�RwE�m�M0LR(�KIz�w�����߰eiW�����- ���b.+��ؕb����)��ʫ�ޏ��!��81)*u�1 �?�=E/f�        չ���t��.�N�f˔m�;��aEg�j��=��M����������0�Ż��3[��^�eEW��U�F�Ri��;���B�m�����v        �F�VʧnMT�%�)pP�Ti�n��]���K���]`#B�q���=��n���"I�w��)�Ի��2Y�Vj-(��*�������LJ�,o)u���5��Y�Fm�˼%��:s�ւR���v�P~?�v        �f�U�Z;�\��;bw�=�nC��	`�X���Re���;��w��q���h๕�;K�v� �Ê���8�ɿ��
��ciu�^tVG�ݦ,v���ٻ�8I�����s���꽧g�F�4ha&`�5��1X2��%�^/�A�B�˵lc_0\r�k�Z�I,1�#;�/c�q�H,�@ �4�]�{-O=�������MU������j��=�|�ݵ�|�_�%39�$7��@a���ٹ}�kܾ1@�Ǫs~\w���u        '�;Bc���:66�,9�(v��Iy*�R��(�4w C���B�Xl&�l�����C�	����>I;b� 0 �6���Wh,n<9b�n�l��n��K���7��K
�5Y�JƓQ�����P����X��x�`��Oչ�[%�!        x���vu����?����B���\���ar��B�*�v�4 ��앱#5�w�{m� Ⲑ)4W:e�֊dy�H[�岬)K�5�kG:o��\���R�g�S���xs���8&���܁��        ������%op�[bGA<��_UY֌ N��BkM����݈�@��������cH^p7sW��  ˚��5��Y�.���B�����벼-�r'fcZ;�q8s�Gjs�wPn        ]u�u�����7ǎ��,��{{cI� 0 k��>/K�D7������CHR;���}��>S��R� ���M��R��ʴ�!`���y*k7di]��S�M�yɹ�!1 ,d�t]��ܙD�m����U�;        ؤ���o~�'��I���qQȎMCvI�c00,K��)�[�s���>���cbx\.��� �e-�֚ڱ���X�잧?�uI�ExR�KJrIA/ȷ��w�!�i�4�	1���U���9        �&W�����_&�7ǎ��L��)o7�G&䊣���,d��Zgx!�-�BxY���cx<&�&v �gYK�zU��H�}��\�5e�U�zU�����Bkuc�w���f�y7�ƒ�y��2�v����*        lΪ��Er;	��
�e���,d�� �j,(4W֫�ہ���=�����c�Ȃ��7�?�%}O� zǲ�Sr�ؾmLyO�7
�G:%�Ʋ,���x[�!d&ˎ/�/m���g�!�
��¡��c�         [�-��Չ��A�;
D�*�W�+��{f
�5�k�v]t= �к"z�����h@�8E!Wh,)4jLt��,�e����S�7^�[������#'�7����!���zYx��x�        ����jCo�����d���t]Nt��B��|}^�����c�}y�.v�ǲ����kb� �M���e�u�dO����\R����y_�j˱�ɲ�,kq�
6��Y�L?�J�(        ��*��e��\���Q0`\"?2!W����3Y��<cy�0 R�Vm�6�Q�6�v�
�g\���ԕ$����;,KZ+S��u�X��%E�o����=�/�B{�ʲ�6�t�K�x�2{�v        00���f��g����` ���Ȥ\�;	��c�vS��F�����K����{��n�mۍ\.����r�֪,k�N�M+Hy�)_�������^���h)���Lʳ��4O90���ua��7�r�v        08n���k+?0��os
��&�5))u��I1v" C���� NJ���(�e�]-����
麬�.�� "Y���鸇���w�<|�4�oh�dy&m)ow
��m[��OT'/�N�\ǫw        0xn����?x͢j����q0��T�^����	�� �e�p�$Y�_s�k���u݇7v OQȕ7��<��8q.�(�'��DrGO}�t�΂,�Ǌ��g�.��-�\r�V���
��       �@�`�Gj�p�9Qr�r��\i��; I�e��b{;v C+inӶ�{�~�c��*��x�����s xj��Ph�����\�t���+�'�sr�wJ�.�C��)�Ǖ�s��Evn����'�G|���Q^�       ��pƵ�����^;�@2"_�+�b'�w&k7�:�v ]�#�X��=���w!Ʀ���;����BsE�5c'z�6ަ);6����\��Qxw�?�N���D�x����l����ce�����c'�H���q�z�Qn        ��۷�\���T�73�i����y0��B�%��|iL�Xր�@�mf
�,��X� �!/�D�]fW�|
.�5�+L��+�o\z�����ym\?�[*i�,         '��*��/�\F��Kᅱ�`��BsYj�ɕ�䋣��l 6
i]֮���&{I���N>��m�4/)���	0Sh��ڍ�I  xB&�7cӯ��-?ǃ        j;���������];���+����
��a ��SYڐeM1j@o�z��i�Q���s�7|<嶽Z�ہ�`!S^�Qn �?|�q%�v        �,���ms�e���Y0lL�55�k�
��ء �(3YZW�^U��dYC���^��Vz~����n�폝������^�B;v  ���Rh�^�p믯�N        �-+����v��2�;���֪���΀ô.Y��
�c����\���Z����\��"ƾRp7'�ձS x"��ZSh,I�E `����r�U����I         �m�3�Zu��J�{bg���S�֊�#�닲v��;[��u��
���]}- �{I�m]�Mm�>|���s x�7���;	  '���륇?]9;	        @/�\������bg�&�r���GR����,Ȳ�B�IG�@1�j�i�*��i3�}���3 xl����Wy� 
f�J
���        ���C��f^(���;6�Ж�k
�jg�tkU���,v2`� k7K���� 0x���������}��n�+bg �ݬ�P��$�cG �I��7���U?�����        �/˷]����4;6����u�FM����E�t]��ɀ�cA�֕����-k��G 2����3z�}�����c� �H���9*�'O �!`�&I���*ߊ�        �ߪ��r��+D�=gRޒ�V�:�Ʋ�ݠ�<�B��|��|�BkecR;�, C�����ܓ4y��b� �2�ƒ,]� �br*�_5���         �Ń��\�_irK��`�\�5��ޛޱ�Y���
���mb}A�Z�B;v2 xJ�����3z�]�];���7�� ��gr�W�n{ם��         Ķpk��\-i5vlQ����ޏ(4��uY����؜L��
�����7�d�dy�p p�,���cW?��^pw��3 �N^�Iy;
  '�䖼W,��cg        G�n��T|���� � ˚�֪B��|�����Bs�)��1d�d�F�}��:�k�t�)� 6+�������w�����tv� $��
���[C ��ox_z�����;	        ����]��·kej��<�I�-k���:��^Sh�vJ�y[��1P,Ȳ�Bk��	퍍B;�L `�0����~�~n�h.	���? ��M��x� �IR��#����Q         ���������()��x|A�SY�>���r��9M
_z�L��e�-�����N �.��vQ'�K��;��u��(� ����
?z��{>;
        ����;��N�OJ.�����ɲ�,]Sh,mL{?�|�ڙ���˲T2~��Y�e�B���XV���|�pg:{kU�5)��g�su��};h��k��R��]w�:,iG���uYk5v  N�����:���I         ���7�����������%�ߓ�ˑg�">3Y�:M��c�98 N�/�;�_��^�޳eǗw<G�ہ((� �����Sn        8y�C7|`��JY
�;��<=6l��I��|���Q��}D��3)Y�%�7���F��)� ����6w�ݛ�<���VZ��t=v  N��Wjs�ߎ�        `XU�*��}e�~&v���Sp�sY���cS������w� ?hl��r�m�n�r=�� �.��"I�ۏ���%��x{[Sh�����1  89��z�P���1         �]u�������_���L�V�8��7�䑅��;��ƬSX�Й����)�@lf�y����k��=�ڛK�n�&i<���V�˲v#v  N�s�?X8t��b�         �<��^��?t�;	��8/�mߝ�F^�s�{���5��If���q9<|���q�C�b ����ON��/��z�(ܫI�{(��a
�eY֌ ��✿y���o�n�        `qV�W���Q?!���Nl*�Q����y�O<���{��9u��������ٶ����;����݉��w���Wظ��p�=<|�	� ��%��z�����FQ
�y�WFl9�� ��T8T��M��o@         ��J�m��]�ڜ\xy�8 $)t�����S�Q �/����(�m�L���/�Մ�
�v ��1�gj�u�uy�,         ��=s?��M]#�/��  ���-<�/��c�����������/�Մ�,kĎ �I�W.�ktK%��        `����������;cg  ��3ӳ��O�'���_$���}�-$4Wdm�� �!c�+iA�y�J=v        ��b�����&���Y   0�̞vƵ��6}/���K��'���֪�M/ 0\L���ܫVo�,��        ����<�
�����   `�9+���K{�M��A/����VZk�t=v  N��#Iq���\�۱�         lU˷]��D�j3-��  �f�z�E_�O���s���{[EH�e�Z�  �$��br����'v        ��n~�/%*]-9�:   ��ɞ��=�B߇    IDATZp�w��K���V�uYk5v  N�o8�k������I         �1�{�Fο�L��Y   0�Bxv���k��ɾ���[���� ��\�Ľya�         �T=t�ϼӏK�cg  ��qn���9��}-����~�lv��
͕�1  8I.x��U?y��N        �Ƕ0w��K~1v   +Ϯ�ua/w�_����Q��69��
�%I;
  '�����^���c         ����-��_�s   `�x����{���v$�K%M�k?`S�F�=�N ��qɯV���1         pb�s�w��ߏ�   ��,<����������~�lj�7%�c' �$��W���)         pr������q�   ��^�޷����q/`s2S�X�B;	  '��iu��O�N        �������?;	   ��^.߿������I�沔��c  pRL�s�4�f�Y�,         x�n��#]#�/Ď  �Ȝ�{Ƌ��h���K������ْN��^�f�+��;  '�����+���V�,         85�V�r]-s���  ������3{�x_
�!qLoNAH�e�z�  ����
�+ks���Y         ��?]9����&�@�,   ��y=�Wk���nο�� ��eMYk5v  N�|�/�~�߉         ݵt��L�6�r�,   �äg�j��eF�x
,o+4z 2��������Q         ��s7}�%��Ԋ�   �gf�j��������.��>�fcA��$)�N �	3S�9���*;         z�z����>�QIy�,   �3��z�t��{å�F{�����ƒd�� \��ma��m��         �?��Ŝ~>v   ��3;K�VJ�X����酽��lBcE���1  8I�����o�         �ڡǜ���9   �GN�m��i�X��w�����LB�.��c  pRL���s�_��         q�U��s�?��  ��)h��^����w�DY��Z��c  p������\�         �ka��w�ܡ�9   �y�E�X���=�~p�L��r`���)4�b�  �$��T�<�F�Y�$         ����r�]+�;
   z��.�ź=-��\����MÂB}QR�� �f�����?ڎ�         ���*����$���Y   �k�^��ӂ��{^/�6S�X�,� �fr��x�­��;         ��m���_m�cg  @��׋e{Zp�܁'ZkR�Ǝ �	3iQ�p�§��_H        �1-z�7gWI~%v   �s;'_����^��ܝ�����agYS��ǎ ��s��8���m7�;
         ���M_rNo6S;v   �F�.���=+�Ͼ��S2]Ы��ag!Shp�2 `��N���*;         ��¡�'��C���  ���ޝ��5��౅�¥�\����)4�%��A  8aA�_Z8t���        ��2���%���s   ����s��f�
�ץ�Zv��"�} 0L��,����S         `8U�*���b�   @w9�s��f�
�f܁�bi]�nĎ ��3�gչ�&v         �����n��;   ������=+�Kzn����m��j�  �03�w�M�Ar;         ��-���D���?Ď  ������fO
�����˒.����в��X�D? 0,���vz�}wT���         `sx�J=)��4��bg  ���rgH��v��\쨵f�^*�bm �ęF
N��TNLEo*%R)��T𦂗
^*�Οi�/)�Zr�F�G��$�'/���{��̤,HfR;�\�N����u�L;Hypj�R����)R�w�� �t�C��ի���j�$         �\����ó���j��wҶ�y  ��9�R�4Rt*x�b���
NŤ�Q.8�TH���JI�[W.:I��:�.(礒7���V�����?Ƕ�IfA���̔�S��������_���ܔf�V�Ҷ�Ly0�B/�]@|N���:�6�owkɞ�]�?C��������i�`-H�E�hb�N��hQשSfOL�S��n4�'���~����;p%��~�3�G��c�O�Y���ʜZ���;��V����S#uj�N��R< l�·���t_�          ؜j��t玫��z��!9+�� ��ђ�h�i�$��x�}���q~��6:|N�%��	�}jN������:�a�y���mS�mZO�9���iP��c�k�M�4���,P��p�!�����%����$��Ƌ���i�d/�L%�XQ��(��M�O�a���jtt�?�m8Z�7�G���~����=���_������:����z*�gN��z۩�9��N9� 0t����޸p�/��        ��m������Ɵ0���d'� D֙�>1�59�4Y���*{M���JN�#N�E�dOos��/���0^���=}ty�#�TϜV����i���2��Ak-i���
��)�#��t���vk���M�lλ���fF��FL�#��d�4U
�*��KOm��fs�S�����<�ef��\c!(<�� [��z[Zo{���ն�J�S~�  �ɹ�g8;         ���C7���+*���M��  ��xM�M�z͌z͔�fƼ����G�Fz6iR�����i�(i����N�-�bӴ�0�4�VZ��f�r�s9�smփ0 �����zRp7�^���c�h�)�fF�fFL�#A����H�x�;�~:Z�O�D�b�	��h�=���d�<�T��B�_�ȜVS��TZj:-�N�-���w ����v����        ���z{��ۯ��/~,v �j
I�m�^�ƼfǼvN$�);m��KO4i��נ��4]���N�q��{8�Z۩V�Ճ�"�b#�J�TO�d�����x���\����?������^�O�K��m����r��i�l*x����^�{
�}�rt�������G��K��>kG���r�i��Tky���
 ��o����T�         [Pu�n_��,�^; lF��D��mw�1�h�������E�Ĵ�Y��O���Ms�jݴ�4��X�U����@a'&�;���u����'/�
�}���rA�1�}̖M�GM�%���j�s*
�[�Ϗ+��e������z����5�9mz-6��m�S�0���ra        �8n�.����|���R�$v V�5;�hǄ׮�D�'�vOx��b'à*%��&��&�:��;�>��Ҕ�릅u��Z���\���v��)�8�s�����^p��_"=��R`�J����c�Sd�9f�14U�N'&I%I�]�?�}<˴m<�YY�<oK��I+-�j�k�鵰�9ߦ� O���+���;*��Y         ��-�Ż�g�|�������;v t#�D;'��L�g����f�hp�;���4]v�`֩S~/�LZiI��M�ׂ�W�փ��߷0��s��ߏ��C�fҿ���,傴k,�=�]c���M�GF���)˲cy���n��d&��NM�j�k��5�p���8&�$���*w��         ���+�ɇ��4; ��B�ݓ^���6�h���(�=�ܤj]z`%�C���+�փ�,�޷ SV�?8�/~�ݍ�~����朮�����������=�g,h����؈���#���v[!t��-���^Ն��F��;���L����?t��          �������͒����`�s�kf�Sh?s���f�vN8&�c(���+A�=����Z�z+�������ڧ��n�U��"�s^��;7�J��g<h�x��ƃN��*��pI�DI�hdd��uGK�c�Of��3���B��H��p��uϔw [�%J~�r;         U�`��WU��B���Y ��F��N�Jt�L��3�t*rx6�ɒt��wx�-/7��WL�Y���r����,���)3gI�J����\���#+��uq��P�N�V�Lf�3֙�~���;
������n��e�L�R���z����z����a ��z����1         �'3{��~�Y���9 ���J��Nt�t���%:m����ڂI�u�wV�\���J��Z&3���go\������X��ܗ&
�x�����N��;t�dgB{����B��B��r�,I23��m���vO����r��u�ֽ\K��@1 C�9�¡�$UbG         �T�2{��߻����� �S5>�謙�Ξ-����1����vN8�H���:��V.ݿd��R�o/�:��)���I�D���Z��w���GK��i�x��A{'r��O�9�R��R�$�Sx��\��vM����Vm��������z��z�����'����          C�R	��T^����H���q �D�ݓ���^�y��N�trtځ�2�Hlw�`{ARA�FT�K�Z
�9��K��mI�`��խ��Zp���{����\gN�:s2hz�p*�sǦ����J��,�d��S�.NS�����zp��;k�Zw�T�����;*��A         ����m�����5r���� ��y�u�T�sg:oG�Sh�
�d��v�K;ǽ���K*��(�Šo-�1�Z3��x\��Z��w����蟉�錉���r�3�Sh��
�Si�3fR=�������}k�龕D�m����L�r����*��          OEm���WV��_K��� &G�=��ق��HT.��mvT��z����RC�����L��r�2Ὧ��-�;�Îzg�h:{�3����\3ent@lG�ccc23�i����ΚI�¬�Z��۫N��$:\�<T�;3���ks         8�*�8{��~�Y�ǒ��y l-�{�Nt�lA�v�s��$0hfF��Q�g�)�3�}T_���f-��˹-&���3�޵����$��Cw9��n�����w"�9ӝ)�ǂ����!(MS�Z-�ig���뉾�����Di;!���\�C~'v         �[���=��;��o��uֶ��ߑ��]��;R@�-6�{�����V��<P��&᫵O���n��ź��]�}x]�h���zfʦ�3]�-�ɠ�q�����,S��R��R;�u��u���}ˉVR�^����s����         ���+�Q
o����39���ق�����{%�z�M)��+N�.����L��B�X���|����V��w�x�����^�@��$��s�3��1�}�H�،�s*�*����P��j�tֶT��S-4��[�o%�R�g� N�������b'         ��:��Ϯ��cg0�v�w
��L�k�ǎ�
^:w�t�LARAk�ӽ�\�Vs�W��J۱#!�Mz^A��)�֢�q퇾�;�ѭ�6��A��:g:���\�.+������Z���4U�!ݿ��+^G�<a�T��LzQm��;	         �+�W�k[!�>/i_�, �϶��.�U�3v�s�����I_��to5��j���'�Y{`������ӵ	����2���Hb:g:輙\�M�gJ;��x�U.�U.�ef�JS�6�ҳ[--6�o,'��r�E&�81�骥�)�        `s[>�k���+����uNӱ� |�&�z�΂�������i *��&��&z�y��e�S�{!ӷ3��Lw<��������-�ӝ��}�Lٴo[��3�J�8�9���hdd�X�}�LK�KS��ҽˉ�]J���N
` �k&.����7�;
         ����]��������rֵ.��c�X��v���=�����q �ɒ��Ӝ.=��<���1}m>�����$��G%���tq�{�k[|���Ѡ�fs�?�k�X���� ����Sm�����Z��M�,%�{��F;)�a��w9t��b         �����|jە7��7�^�, �x)Ѿ�]����g(���K�m3��-�O���������S=���,Ď�?Ӎu�8�ݝ�-�8���ɠ}��.��5Y� ��S�TR�T��Ą&'S�6����i�;�^__J�e���!`�rɯ�:���1         ���o��r�,�3v q��};Kz��E���o�:#�Hv�K;ǽ^|vY�M�+�A_[���R[!����y7Xw9�޵�X��Ο	�p6׹ӹFڤ �����驖����z��olLu��St`K1������N         DS�L?5�y��)�*v ��t涂�uZI��*&tf �3]�^p���,����kA_��t�B�|˔��t7V�^�]���^J��3]8��������`08�T.�U.�5�f�[�dWC����(���c��[�F'�Dr<A        ��V�������tq�8 zgz4��w��E͔)�<��Y{�����4/�����m}��V�e����ug�{w��+��]MIŮ�7 F����ؤ���� N\��j6�j4��β�k�����(��
l*&����js�o��         �]�o:?S��N�;��)&^�v���%�=C��pʂ��U�]G2}c��v��&ؚ�j����NW&����ޝR{���#�i߶�g3�3�+��`H%I���q���kj2չ;�Z��t�b��T-�x�=�2��r;         �HG殿w�����B~й�3�تv���%=�D�� í�M�.�YP
��6�;��z��v{Lv�0Սe�Rp���k8���3�3�)�_8��8�� �J��J��&&��O����=���Z�{eLu��y��9?W���A         �AT;t�Ϸ���H��bgp�Ӆ��z��%�=C���T�҅;L�(*����h���>�*����"78w����(�s�r]�=׾m�J	�N ���^�����T�3gzA��{jNwULu�������+��         dչ�q���[cgpbvNt�ޒ��'���l!�3훕���|ZQ_Y�ݿ��VCTv6ݍe�Rp�޶����I�;�)�_�=�h�R;���P(hrrR�>�ҳ�4���\_�t߲����2�o��@���c'         ����9���������y�oGQ�sfIg1� T.H�����=%��Gt��\w���r*�;����2])���m��o�>��.ޞi�De ��S�\V�\��d��v6T]m��U���
jd�x$�U�~X�ʀ?S         �?�n���b��d�Ď�a�D�>���Q��Ȁ ���3�.;���fI��P�;ʴ��J8��9W��:])���3��M+J϶��������qt�����v�4��Ӛ��f���h��ѱ@l&-&ő��o}�J�,         �0Y�������q�}N�d�<�V�w����-��yz� p¦��K�I��s=�V��| ӗ�j���ю1��ܝ¬)�#M�s�r=}G�}�r%<��S���ؘ���45���=����'��R""0�%���[�}O�(         �0Z<t�?︪�#�'$%�� [�s�;F�³�:c�A� p�N�0���D߿oT�\��|�������Y�\f68wsn[��������_�#�hap���fP*�T*�41���ن��-}y���jAi;�u���v������         ����[g�Wnt
�*J��%{Jz�9EM��Z ��t�t�LQͧ�Յ���;�R��=G�~����:]9q쒫��szZ7�:A:�ǝ�o����8}Ҿ��A] �3�{�J%MO���i��[Kr���Z9/>��r��U�;         �4�����|�dϊ��̦ˉ^t��^�̲.�U�H�~	 �Z�K{&�^xV�ѿ9<��Ω�L�da�_�,m����^:���]����n��$ڒ:����Ço��L����>� ��S�\V�\��TK�����2�ӑ�(b7    IDAT�M^� �f���6�࿎�         �L&z�꨻X����l6{&�z�9%]�+M ��9����?U��sz�G�ݮ#k��Y�m
�岬+�џ`��t�]y�u݇�Y�3��֣9g_��>�B�?�/o;|��~�7�"I_�ž ��e�����]h럎��:/O�n0�[��?��+Gbg         6����3���퉝�Ι-��t��& '"H�����_��u9M����o�<=���?&���܍�6ʺ2�]Ҷ.�sԚ��l�;������}����9�� S�P��Ԕ�5�k߮��Gݷ�cG���{^wx�r;         ���ʷw��r�>#���y�a�Ӿ�E}�9#:m� of��t��W.|�J�Q��v\��/Us��Ph�ukc'�t�9��/~��Ic]���������.���O��s��ζ �S�$�&&&t������Ѓ�}�׽��B�p�p19����          �ّ�>����,�p�,�0���{��޳��6� D D�糶p��J�_m��#�I{��-K߮�}�����-\\��橬ѕ��I�S��-'�*飇o~�_���T*%I/;�} =����ؘ����-Yj�2}�Z��� 3�[���9v         `+X8t���^Uy��m�� ��{�Kv���J�.3� �	_��˒~[�oo�o?_y���?���>Ս�Q�<�?{T��z*�����b;�=|�;�;�r�$MMM�H��S� ��9��e��{F��hLo~F�g�̔��x��w�і���w���]-=XT�# }�"��51AA��c<)-�x�j��Z�C��kNr���p\8��hc�����{Q��F���f����D��ݬ�޹���>V��>����6�?���K�yC�      ��L�����\}�t��fU�	ƫ�6/8fH�`~X�q�ƣfr���x��'>�_^���jp�?Gc蛳��w�ι�ޅ�9E�g`�ޕ">q�ͯ�XDʳ��n��Mɍ��)�?ix8�Y�3N�{��Os|cK3ڳ��s��ݻw����.�      �/����j�pw#��"V��u1Ш�����kc�R;��SUչ�^�o[�������w_yjx:�w�c�7���[�Sn�+��_�<�����>�r{DDJ��r= �744�"~󨱸�v�w�Fw���i[s0^��co�(      �{?Һ/��#���@iͪ���?z�X<��!�v�y*�t�\�xd�{sh�Ս�%����]3\5缀}�w�}^����������v���} >њ��G��mo�kpp��BA�rv��[����N|��ftJ�2rj^��k��t      X��yΛ_�I�,�JH)ű�obc;��uɒ%{]~�廻vb�U������w����ψ���Fg�OW?�鿸k.c�ܐ���]��iG��%�������W�z��<;������8p���{ٮ8~����{r|{�sz��;�u��      P�߱��z^��ȝ?*���J)�� �>t(�)�,$K|��3#�S];���������^����ij�k�ԮK��{����f5����;c�`��"����6����7�jr��>�n���>c�~����q���?	Ew����<#�16�N      <b������zr��9��@o�8b��8簁�k̾Y����:��+�������FīW^t�Սm;.�w�6ڻ����9���|�T4n�����}�Vg��M�o�i }444�����Ll��q?��(�T}'�zI���׿�      ��h�:��j]��_H�Jǁ^8t��8����w��v��,��[���3&�v��#���j�g�-{~~x���z漻;]��GG�7K� ��v��߿������nWtg�i[c0=����Z:
      �g{�N�Լ;>�)��e�%�8爡8dE�t ��]UվW\q�d� 31ۂ� @��OZ�0����K'�nH�\U�)�     @�m�p�Q�WGD.��j�h3~���x���� �K���<�t��Rp��RJ1::��<.>�O?���S��j���/      xb�o���ݥs�l�6⷏�?8s4��G�`��w��yUp�{�;�,���K)Œ�8��eq�U��;��]"rT�8=_[:      0}g�k#�(�f�Q�8u�p\���8��fT�t" 
���fj^ݶ�����"�S�s P^�ݎ{x(��G��֤'���釻w�:u���>Q:      03�?�m�슝_J��T:<�#��s��eå� P�F�u��}�t��o�o�U:  ��h4��������c��\:<��᪙�Sn     ��駛�xJ�EN;Jg��r�����x���� <Z�ݞW��Vp?�t  �e`` �<pY\x�p<��v,Pt�~RJ����R�      ��MlZ�O��ה��j�p�۱�q�)#q���V	�O�{��jGę�s POCCCq��q٩����10o�p,t95޻eӆ���      ��䦷�YD���s@DD�������g��S�o��@�=;�J���yS�FDxq
 �)��#q�Q���8|y�t$��+�זN      tϒ��U9������v�>C�O�s�fc��(g�o���!�k��SJ�� ��PUU��x��	K�G�X>�KGbQ���4����y���I      ����'Z;���H������=ֈO�?ˇ���v�����k��s��*�����l�q��ť���������1��4�S��[[w��      t߃�����^^-N_5S<��x�c�z� 3WUռ�bϋG�6nܸ��hLFD�t 槜s������N�][���y�ͫؼ���9      ��Z��7�%E�M�s���P<눡ў`n<����:���k��޼x����g�r; s�R�V�������|(��ĂU}@�      ����7�T�^:�^c����x�����ew�u�ɥCL�|)�ϛ�� �[�шc��4.;u8�vP'�ŝ�y#���KJ�       �%��qa��;���p6R<��x�cq�r� ��٥LǼ����誑�8��eq�	�8x�m�tC��48���?��V:	      �?��[?�"Ώ�.���������*�N�B�R:�t���-�mo{�^�����<)�0�LMM���=>��"�]:�T����ۆ��t      ��}���WvR�/K�`~Z:\�o5���(�,��}```�ڵkw���xj_xṽ� �_�f3N\�4^q�P��o��OQCջ��     `q���Q�u��?�0�:cL����9�NMM�Y:����g� ��0>:�9vi�wl#��N����41W�N      �71��T:����f\t�x����jZ�@t:��w�k_pO)�S: �GUUq��c���G��6wW����L���v��      ��-�]�j��9��Q���R��j8^y�H���> ���ͮuo��ۿ�������s�M|kW��p�o��:)�nټ���I      �zY��7��r�戬�̣�5ֈ�3-�� �쬪j�W\�p� ���w�F���3 �x����F����'�z�4�՟*�      {2�i��s��J�>U���W�1��@iC�v���!O�NG����qΑ�q�Ƀ��X.�Z�>6�y���)      ���<#�̩�T�����f\v�x<�����@������Z�SJ���`�H)�+���S��7V����^ʑ�i���i      ౵Z��=𒈸�t�hT)�:t$.;}4��l�>rε�h���y�M7�k׮{��X��}pG�ݿ�os�ZLr�]Q�3y���-�      ��~�[��c꣑r�t�g���x��C�lD� �Zڱm۶�VkG� {R����w�>;������ǅ���9�T��/&��F�      ��-w��9�?)���jV�ܣG����������SK�x,����}�= 4��8������8`�tz����7�N      �?�w�K�js���A˚�3��ăJG�'�R�mW������_ ��}��E���%�Y��更헔N      �W)�޵��qW�$t_U�8�������X>�9 ��P�e䵼��p�+;���Q�> ���'w�m��#�Y�[,��cg������JG      淽^��b�ԧ"�P�,tǊ�F��ؑ8h�� �KJi�֭[W�Z�]����Z�U���3��� ��<i�P����8q�#5�)�      �0q���w��s��0�<}L��y)�<�dɒ�K�ؓZ�YSJ�]y Odh��9f<~���(��9�Շ&6oxO�      �����6�H�J�`�F�������@�t ��N�S��v-�qv�  0)�8j��x��q�J��磜�t��/-�      Xxv��uI��Q����{��9G���������v��w��˚��DD�  B�9�|�����MŮv�4LK��1�|�ĭ�?_:
      �0�|��<-:��L�Kg�6�8���8m�W���lݶm��V�5U:�/���F�qV(������U�q���q�x�-cOR\��      �����~6��U:Ol�%�x��c�� ,DK���O*�Wծ�^U�3Jg �^�{�`����8kU��+T�%Շ'6���K�       ��Mޞ��\:{V�g���N�����`�:�t�_U��{���3 @�4�xƑK�%�Ÿ���N���qq�      ��{�΋s��K��і7⢓G����m`�cw�V��n�i("N-� z�}����ơ+�\9v�Ըprs�祣       ��֏�}��r�ݥ�������>OZ�( z.�d���ٱcǩ1\: ���P3^|�x���j���T]3�i�?��      ,>�m^����ͥs,v)�8��xɉ#1:��| �����#J��e�*���	  襪J���F�'����˩n���zW�      ��5���o�)�Q:�b56XŅ'��3���{ ��u��Vpz� P�ꕃ���b��Zݚ����t      `�Kyw#]�#�]:�bs�ʁxՙcq�
���8UUU�wm��9�O-� J�ₓ���C�s�^�r�j�t��>��Y�(       [ommiF��i�t�� �g����4�ֶ�x�k���Q:�#�,YrLD\U: ��R��Wē�������.�h�K՛�ln�M�       �x�w�h��sS�KgY���F����� �׹����~���Q��Q��? ��f��x��c�zy�n�L��ؼ��c       ����cC����9�5+�Ug�������"��C<�6w�sm�R �Ƈ��ऱ8{M�>7�"G����)��      �kZ�Nj\Q�_:�B�R�3W�'��蠽� ��RJ��rצ/W�� ���J���F��c�Y:�B�:UU]6q۵?.�      �L�v�#w.����`l��4�>�� �Gg���Zܫ�������I� Pg?����O�uJG��rT���ZW:      �t����{"w�S��فK�q���1>T�}� PG��m۶��jm/�w쪪j����Z:҈��:'�(e��9�29W��      0]c��՗K瘯�;`0.:eD� ����%K�("�&����Kg ���٨�9ǌ�o9�Z��e>�~�h�8ni�*�      `�ni�F.�����2�TU�s��3��� 0M�XZ^��{��i�3 �|r��x��#16���"��ۛ�S:      �Lm����JU���9�с*.<i4N}R�t �WrεXZ^�w�7�t:��E�`�, 0�<�������w[�t�zK��Llj]\:      �\����-�鼨t�:�I3�;~$����|��m۶��j��Ҋop�t:��r; �ʲ�*.9u,��o�t��J�w�����1       �*w�9��K稫��KNUn��[�lٲ�J�(^p�9?�t �Ϛ��{�H<���f��;�Q]t�'Z�JG      ���ͭ�Gn�,��]:K����G����F�F �o�N�x����<�tf� ���z(�?q$��j�ȍ�ډ[��t      �n��c��"5�Z:G]�T�ғ��7KG���ˋ�#�� `�8t��x��c��xn������7���1       �mr��?�\�Y:Gi{�5�姍���#�.*�������_��  ��*.9e4�ާQ:J19b"�͋#R.�      ��R�f��iK�$���@\v�h,�s �c��w,+�h�=�T�� �@��>e4�Z3��G���z��m���t      �^����W�Z[:G���♇��yǏ�@c~# �W5��Ӌ(9<��Ԓ�`!K)�3�7�����>W�_Nln}�t      �^۲i��"US:G�4�x�q#����� �BW��]����� ���`\x�h�.��{��3\��J�       �j{�:"�W:G��T�ғG��}��� �bpf��Śn7�t�Ю]����R `1ypG'n��ñ�v�(=�#�J��Y���|�,       ���3#w>�R,���+G�Gb�H�}� �h�l۶m{�Z�N������w�>%���o�Wqɩ��f����R�Rn      ��ͭ�T��t�^8xE3.=mT� �k���������真Zj6 ,VC�/9q$N8p�t���Q}rb��w��      P�����gJ����N��f* ��]��Yp6 ,ZU�xޓ�㙇���9�h7_�r�,       ŴZ�Nj^�#��t��Jq�!��c��Q)�@	)�b]ow X���f0~���h��5R�?M~����      P��6]����xM�sѬ����F��.�7��<T��]��o��v�}O�� ����`;��W��C����\�?w�^^:      @�����ˑ/(�c�F����Gcղy�� ������׼�5��=�ȿ���%� ���e��䔱X12��AN߭v���      P7�H��H?,�c&V�6��S���F=��I%����i�� {�|���N��+���LW������Vߟ      ���ͭ�Gn\9M��2�V4����b�|[� \UU��[bhD�� �mx����8��7P:�4T�ۼ�3�S       ����?��]�s<�����8��f ,*E������sNqJ�� O�Q����F�����8җ&ƏY_:      @�M���7樾\:�c9u�P����hT�t `ϊ,5o�{�ҥK�����= ���+�1�H��ɺ���z87;�{�|o�$       ���/v��|�gS��"r�^�}�������| ���{�{>�я>�ϡ}����� �̜�z0~���EN�i��7N���o��      0_<�i��:�j���c��<�~�!���  ӐR:��3K�O+0 ���n�Yj�FD_��۳�&7o���)       �6�靑�;K爨N�:�)4>Z:	 0=)��/7�{�=�� �C��n���o������
�#�/�H�T      ��+��@\�s<X*A��`���'6�>XU��J�  f�D��������qb?g ��񫯾�����6������o�~R"HjT���ܺ��l      ����[[wU��k��龪�����wFDLMM} ".� ����������>%"F�9 ���ң����C�|-7�̈�[��Q�<q[����L      ��h�m�6��@_���ݩ��[n������zk�yS_s  ��R���o\�ϙ}-�7���� feWJ郿���ںk�9~VD��=]�}�Ow�Q��s�    IDATf      ,|�;��~�ʩ����Y������UU��=] �O���k����Pp�y ����+������s��T��̈�=NѩR��[?�Ɖ��      X<~�w�ɪ��srT�ɻ�~��������n�z{D<�� @w�n�=�|z?� ���O��KkۊX���Շz� ����Mo��g�      ,R[n��)���݄��������,��Z��ko ����[��hD<�_� �Y{�����D���;'Όߏ����G��32����?      ����FzmD|��禔�r�xQ���5��?��5 �RJ��Z�����6hll섈h�k 0;)�]u�UM�íVgbs�9һ���su�ݷ\�p�      ���skk{�/��v���Uu��Mo��h�:����m�>�vk> �3�###G�kX�
�qJg �7�'�'7�y]��-��Su���?׍�       xl��q�sTޝӪ��������Vk*"�ߝ� @/5���5�o��R��P ��=�u�֏����ͭ9��8��+��7��       �ie��&r�׹���Ӊͭkfy񌗰 E�m�y?7�+�@ͥ��{���5��'7oxk��ED��9��4P]���kw�v>       3���kw�@㒜c�,.ϑo�ؼ���ο��+??��� @�,��Vk8"���, `N��d��ۯ}WU�6"ufr]J��|�����      `f&n]����fxY����6�}.�SJ9"n�� @_��sN�ԗ�����S"b�� �Y�oժU���A����?���ў���'��[�1      �����7圾:͏��j��6mxg7fWUuK7� zjٍ7�xX?�����i 0K)�����,�?��7����j��%�iWjƥqKkW�f      0C_�����tq����l��x������n�^�n�SJwu�< �7������ӗ�{J�/ `�r������~�_WU�9���ӟn����n�      `f��p�9U�9MEռl���͹)��s�P7� �/�ԗ��6� [�m�vg/����D�.��S��K����i/�      0s�gě#W��W=�؝�ꒉ���M/榔��� 躅����j朏�� `Nno�Z;zu����3R�pnv.�[�o�j.       3�juR5xqD���/�H���E[6mx_�ƮZ����W� ]qJ�9�zH���E�P��  ��s�����6|(�ꅏ�O�NTo�������\       ff˦7~;R�'�����λ����r���ߎ��z9 ���_��^�y�=�tJ�g  s�shh�~��c��E�~'ru��w���L       fn���1��X��y[6��R<O)�|9 07UU����^H)�� ��߯]����6qǆ�E��)�k&       3�ju&"�ѿ�v�n��������_3�;%"���=��'�a 0K9���r;      @�����V��#���~� f������ӂ��7��H)=��3 �9��o-       ""RJ(� xl)�{=�����눜�h/g  ��R��������       SSS�EĮ�9 �Ǵ������z9����s�� ���=�      @m\s�5��>Q: �ئ��z��i�=�tB/� ��h|�t       �e��@���#�ӂ{�8< 0'_^�n��K�       �_�l6?��9 �=��tw X�<�      @��u��7"��t `�r�'�����o��}"��^� �MUU
�       �R��w� P_G�Z��^޳��Ν;mo����W\��!       `O���; �Wc||��^޳�{JI� jʓ�       ��W\�݈�F� �c�YW�g���: ����6��        �'缹t `�z��w X|�t�       ����z��'�V�5G��l `�>�v�ڝ�C       ��y衇>[K�  ����s���=)�/Y��؈��� ��y�      ��k�Z�RJ/� أ��|�;���=)�眏�Ź ��5�;Jg       ���9o*� س��N�ɹ�8T� j�_֭[���!       `:��; ��q�8�'���z ��ͥ       �t]}��wG�7J�  �h��s�O�Ź �ܤ��      �Wrξ��z�Ig���n�aeD��s�9{h``�ӥC       �)�@=q�7�t��^lp�� ��ck׮�Y:       ��ҥK?�� ������Q�>���v��� ��v       ��/�|wD�Y: �몪�zw�܏��� �5����        �d� �S׻�]/�WU�� 5�s��u�_:       �F����t ��r��.��S���n�	 t�'�      ������#��s  ��RzJ���j�}�ƍ�"by7� �B�      ���w� P?�n��Ʈ�ǻZp���y `��T�       0)%w ��v���yW�9gw ����]�vg�       0��㟎���s  ��RzJ7��v���� ���9�}�       0W�_~���d� ��圏��y]-���lp��i4w��        ݐR�x� ������o��Gu�< �+�[�n��K�       �.�� ꧞����C"b�[� ]qgJ)�       ݰu�֯DĖ�9 �G���|��:�k���1�: 莔�'�      X0Z�V'">Y: �h�F���:�k�N�ӵP @�(�      ���} 5��e�]+�����^���+�]:       tSJ��3  ��s�����Z� 芏�        �v�W~3"~Z: �(����sNqt7� ��+�       X�RJ9"|' �R���ƍWEĒn� tG����<       ��o P;���o_э��Rpo6�O��9 @�|oݺu?,       z!���� �G�J��+���Jy �+<�      ����7��{���9 ���s�J��+���� P#^�      �"��� ���s�� سN���       ��RJ��@��g�{���n� �]���W_}�=�s       @/MMM�}� �����w��]�E�^]� tAJ��3       @����o�� �B�y�ƍ����9�;���� P#^�      �"b	 �Gj4G���n܏�� @���?�       }��� �G����9�s�
� P�z��_��t       臩��ϔ�  <J��)%w ��ϖ        �r�5��?*� �ws�Ϲ�ލ @w��      Xl|W �Q���j�#b�\C  ݑR��5       ߕ@}�sNs9`N�e˖͹� t�ĕW^���!       ��:���; ���u�]w�\�S���n�y�< �5�M)��!       ��֬Y��Z: ��fsN�9�s�
� P�-        �����oG��,� ���v��TpO))�@}(�      �(�}g 51׎�\�G��z �kvo۶��C       @	)�ϔ�  �B��s t͗Z����!       ������ED�t  ""��o�ᆕ��\� ݑs�$:       ��ڵk�(� ����o�ᆑ�^<�{�ݶ� j���ϖ�        %Y �QE��s�xVRJG��Z �����>W:       �d9 �G�y�]�Y�c�z ��~p��W�S:       ���tlp���t:���
� P^�       W]u�"�ǥs  UU6�k�0w�C���5       �w�+  ��9�� �U����9       ��%q PG���Y������+f; 莔���۷�t       ��ϗ  DD�A7�p��l.�U�}``��v ��n�ZS�C       @l۶�K�{t (/����fs�
�)%w ����Jg       ��h�Z�#⛥s  ��Ϫ��j� ݕRRp      �G�]: �@_�9gw ��      ��RJ_,� ��t:�+�϶M t��m۶}�t       ��N�cY �@_7�G��; ���V��)       �䡇�JD�.� �]�|���n�iiD�;�a @��=q       ���j툈��� ĪV�5<Ӌf\p߱c��� P_,        �(�di �W-[��_4���Й^ t_�Y�       ��[��:��a3�f����[� @�=x�UW}�t       �)K� �:�Κ�^3�{Ji�L� ���)�\:       �ђ%K�;J�  b����#b�,� �˫�       �1\~��#�k�s �b�RZ3�k�`~�*5       x|�/  ���^3������ �F�a�;       <����q PX�7��t�M�DĒ� �j˺u�~X:       �Y�ӱ< ��{�ƍ3�Ϩ�k׮53� t]���       �V�^���x�t X쪪Z=����� t_J�K�3       @ݝ����Z� ��UU�fF��ɇs·�( �u9篔�        �����N��f&��Q�=�d�; �R�j�       0TUe�; �7���
��f�� �kǶm۾[:       ��v�9 (,��f&�Wp����Vk�t       �:��W#"�� �Y�y�L>?ӂ��3�< �]^�       �t�5�<w�� �Y�6�_��{GĒ� �(���       3��� `��{�ƍ��O��^U՚Y� ���^�       LS��w� PXUU�����~��鬙U ����       3PU���@a3Y�>�{Jiڇ =q�UW]u_�       0�TUe� 6�e��.�GĴ�� =�n       ���:���p� ��M��>�{�yͬ�  ݢ�       3t���#�_J� ��,��f�����i
 ���J  ���Ǯ�>���6g�CR%[�\�
I�6E��.�m��A����.�`A�ݹ�@S&��WзiP�v
[�*�rdQ_4CΜ�za����e�:�����9$�;ba=��     ��r� ������< <z�8:l      ��Lw� ��#_p��7�O<` ��m��g^�       `�� &O�>P�@�R��* ��y6�m�       �hmm���  S������|�@�q� �ƫ�       ��:u꣈��w ���|���|�@��<�? ��Tp      ������; L�A;�*�GĿ~�$ �C����        ���; �Uk��A�w���A�1 �p�����       `�e�O{g ��;���Aܟ�  ���:y���{�       �%g\ :��u�Zp��Cd ��^z饭�!       `��Z�����}�gϞ]��g: ��      �!���+��� ��w�yg��K�ܷ����h�  H�       ���  6���_��K��K)�� Gf:\      ��ad :�a�n���Z�w ���       #s ����3ӂ; tt��u�k       x2�� tt�n�w Xl�����       �	w �� �t� ���      ��|���#�Z� 0a��~� 84
�       ���f���Y� 0a����< p8j�?�       3�� ��Z���k�
� ��0�       �h���N2s�n���7�x㙈8�� �e>�[p      �G(3��@?O�;w��^_سྲ���< ph6�^��^�       �8����� `�677�\q߳�>þ� �����l6�       ���|�����s ���9¾g�}>�[p�~~�;        <n^}�����9 `�����_y�Y ���z       �ǔ;y �d�/��Z��h�  ��?�       S?�  �����=��/3sϿ �Z��4       �s ��C-�g� 8<��\�       ��9 �g�����Z��; �������!       �q�����+��f�#��#� ����l6{�       ��Q)E� ���l6۵Ǿ�/�x≯��{ ��d�W�      �!y��/D���9 `���<yr�!��
�{N� �ǫ�       �p��~�_��kW]� �8����        ��Z��9 �$3��^k���� �!       ��y ��
�{�% �p��5h       p�j��������w-�����É �^�t���!       �1g� :y�ww ����l�Y�       �8�Lw ��wv�Ů��x��  �s�      �C�����{� ��z����	 8<�֟��        ��_|q��� �����ZkF�- ��R��;       4Pk��u �����z뭧"b���  ���       md��; �q|6���;��qܵ .�g       h#3��@'O=�Ԏ�������Í �f{{��3       ����n� 0U�u�w,�g�w �����Ƈ�C       ���{g ����|����� }|0����!       `
�����3 ����^k�q� 8\�VO�      @#?��>����9 `�2s�����ݾ ���d8       4��5">� �h�Q���w�{ �w       h�]= ��cg}ǂ{DXp�>�      �-o[�>��n� :��*�      @C������q�]� �0�
      ������-��Z3"�p�q �{d�C3       4���� �����x�g"�ȡ� �v�������!       `b��@ko����w�������Mx ��y"       [__w_ �lnn>{���)����{� �Z�'�      ���~��W"��9 `�2�q�{
�a� :�LO�      @F� �w X`�       ЇQ: � 3���g��w� Є�;       tPkug }��^kUp�2���       Ї�; tp��ء ��tX      ���@7�/�G� ����       `�J)��  STk=Ђ��d �t��_��       �h{{�W�3 �D��S 8t�        SUkuo }�]p��ff>�. p��2       t�ꫯ^��+�s �}���Qp?}���14� DDD�ի�       �/�t ���ٳg�?��;
�kkkO�� DDd���       ���= ����uG����˓m�  ��)p       �֪� ����^p���; t��       ݹ���qܽ�^kUp��      �/w� �Gf�����/�6�qtH      ��J)�����G�-����~�;       L�w �cς{DXp��6^{�O{�       �)Sp�>J){�-�@{�       ���֖�{ �㎑v� �Yf:       @g��������; LM�u���	 >�8      ��2�f�{� �	ڽ���
� О�;       , #u �����{��d  �}�;        F� �� �H<�       ��> t�{�="�j ��̴�       ���� ����[��gϮG�z�8 0q�8��w        ���Q� 0A'f�����
�yr�� �i����        Dd��; t��3�<u�Ϸ
�����>q `�677�      `d�;| �`kk�V��V�}Gw h��l6��w        bG� ����H5R:    IDAT
�y�O �4O~      ��X]]Up��a���^J�� ��Z�      `A|��_�c� 05;.���h� �Lw       X/���<">� �&3ou�-�@_��        ���: h��j� A�ա       ���@{;�3ӂ; �g�       ��| h,3o�����\� �s(      ��m� �ގ��D�, 0i^k       �E� ���7������� .�       �X��@c
� � �󹧾      `�x; �WkUp�E����P       �ł; ��� `~�ҥ��C        ���h� �Sp���l6{�        n�A� ڻ��~�����X� �Ɂ       ��˗��@{�f�Y��Qp��ώ�� ��q�        ��f��fD\� &&��׏G�(����D�< 0Iz        vt�w  �����7
}� �$9      �b��w  ��������|�� �9      ��Lw� �����Tp��,�      ���*�@c�����8*�@{�       ����@cw�-�@{^g       �ɝ> �ws����|�c ����        ���*�@c7G�KDD�Ղ; 46���      `1�����Xp��v �)�8      ��Lw� ���q�c ���|~�w       �^�8*�@{�#,�@7+++�       ���� ڻc��֪� m]{��7z�        �� ��촗���-a       XP[[[���=� ����       ��=zT� ڻ]p�Lw h�A       ԩS��E�F� 01��7?  m�Z�      `�y;; �u<B� �(�8      �b3^ �Z-�@/�      `�e��} h(3�(�� &'3/��        ����� �����A `rj�
�       ��.�  S��ke6���8�9 L��;       ,��Tp��j��-�G���Y `��      `����n �f�ّ�����;	 L�C0       ,6w� �������0
� �X��R�       ��J)������������ �e���      `����n �a���󣽃 �9      ��� ��Zp���C0       ,6�u ��Z�Lw h�!       �|>w� �mmm���Pp��������!       ������ ��0GK��h�  01Wf���;       ��R�w h,3-�@�       ����w hlǣ%3��-`       Xp���� ���\+�֣�� ��8       ��;u�Ե���; L�Z�� Ж�;       ,w� �P��h�Lw h�R�        ������,�@��      ���� �̵Rk=�; L��/       ,��t� �Z��R�j�  01Wz        �Wku� mYp��2��       ���;  L�Z����) `J�qTp      �%Pku� m-��� e���      `	xK; 4�Vj�G{� �)q�      ��a� �Z+a� �Q�       �@��? �uT� +�8�      ��v hn�d��; 4d�       ���� `b�J��H� 01�       �j�F� ���J�u� �d�_       X�� ��%3�����m�_       X����D��; 4�����       K��z�w ���J�U� �v횂;       ,�R�;~ h��:��Tp���~�i�_       X�8�����
� ����^zi�w       `�֫�3 ��d�P"�� ��n       XG�q� �Z�Rk�� �8�      ���L� ��P2S� �Qp      �%q��%�� �V)�� �x�       ��l6ی�y� 0�9��(�� ��l�        �w� �H��H��#�� ��l�        ܗk� ���C� 0!�       �\��@#��A� �L�^       X.�� ���JD��A `*j�
�       �\��@;���Z���      `�x[; 4�� -9�      �r1f M)�@c�       �\��@;
� ИC/       ,� Д�; 4��       K$3��@;
� И�;       ,w hG� Z�T7       ,cv �NQp���qTp      �%Rku� �%"J� 0!��      �%�m� Д�; �TJQp      ��� ���w
 ��q=�       ��]? �S���R�C/       ,� �Hf�c�  0�V�^       X.����Z�h� ��       �%3��@;��%�       �\�qTp�v�w hK�       �Hf^� &d�� ���;       pp�Vw� Ўw hI�       �K)�]? �c� ZZ]]u�      �%2���� `B,�@Kׯ_w�      �%2�1; h��Z-�@Ckkk�       �Dj������K�Ղ; 42��C/       ,��|�m� �N-��� �lmm)�      ���]? �SKD��S �T���{�       ��w hj,a� �pႧ�      `�9r�]? �c� g���w      `���� �T� Ў/       ,�a���  2�̴$ m8�      ���� M�Rk�� m8�      ���� M���w       X2����D�w hÁ       ���֖�~ hǂ; 4�e       �d�����@;Ղ; ��n       X2.\p� ���^       X2��l��y� 0��Z��w       XN�{ ��Kfz� ���        x �d����d��      �rr� ml+�@#ޚ       K�[������
� �@�U�       ��; hf��Z��Os      ���v hf�D��; �1�        <�v ��v	��@+Gz        �j�  0�V� ��z�        �q� �R�J�U� �p�      ��t�w  ��q�Kf*�@
�       �d�y�!"Vz� �)�̭
� І�;       ,���{�z; 4Rk�.q�w �^       X2�i� )�l���� � 3���        �w h�ֺ�� ��Z��f3+�       �D���zg �	�(��; LœO>��       Kdw� Ўw h�S�       �\�qt� ��Z���R�C/       ,w� �Nfn���� �����       K�]? �������t�      �%� ��Pp����;        pp���q-�@K�8>�;       p_��;  LEfn�q7{�����;       p_���R�f����� ��(�      ����f(�@3�8^)�0\� &���       �������X� �b�+e>�+�@;O�;w�D�       ��2ӛ���#G�\)�y�w �����.      ��� moo_)W�\�� ���|�       ��<�;  L���ǯ��l�[�� �T��B�       ���q��� `BƏ>��r��ծQ `Bj���;       ����F� 0!Wg��x��~�k ��_       X�;  Lȕ��Qk��7 L��;       ,��lv$"^� &�v�=3-�@;�{�����!       ��;v셈X� &�v��� ���+W�x�       �0��; L�Ո��K� �}�w        `w��?� &�b���ŎA `r�      `����>��]p��c ��?�        �]f�I� 0%��I�w �"3�]�       ��j�YkUp��j�#n�o~  ڨ������Wz�        ���[o�O�� S���F�(�ߜs �Y�z��7z�        ���� ��8�������|�0       ���o{g ��)�\�Pp�n2S�       �;} h�f��DDd�'}� �$9      ���Zp��J)�F�(���h� �s      �s�ܹ�B� 05[[[��� ��WΞ=�\�       �m׮]���ѭ �Y[[�q�?�W^y�jD\� &hǿ�       �m>���� `�������;�2��S �2w       X �w� �ާ/���Vĝ��t
 �Uku(      �Rk��� `�n��+�@G����lv�w        ����_���z� �	��eWp���?~��z�        "�a�� }�[p��*�@�;        ���� �(J)�       � j�����Z��7�|������u �0�Z��;       L����W2�s �}��n� ���3g��N�       0e�.]�fD� &�V�]� ��Rʷ{�       ����� `��`��Z��w       ���tw �(���qH      �N�y�!"�c� 0U�0|t�Ϸ
�FD� �����_�       ������ӈx�w �����o��V��ԩS�"��.� �\YY�O�C       �e�7�@?�^{�7?��~�a  ]8,      @7�;  Lؿdf��A� ��;       �7��J��۽s �T�Z���
� � j����o?�;       Lɉ'�,"�� �*3���]p�u  ��k׮���!       `J2�ozg �)�����w ��̿�       ��֪� ����� ����       �T�>}����V� 0e{.�g��; ��ܛo��G�C       ��R�KD��� SVkUp�E��g       �Ff�������Qp/�(�@g�       Ќ;z �lς���~���j� �Cf���o���;       <�Μ9�BD�^� 0u�8����(��f�1"��@G��c׮]�v�       �8+���� ����+�\���_��Q `����       g�����  ��]ߩ���~ 4Tk��3       ���ܹs'"�?�� ��]����������9s���       ����������s  (���% ������       �1��� ��Z����� t�0       ��l6+�w�s  �����8~�& ��?�я~���!       �qr�رoEėz�  ""b����ʊw X%3��w       x����� � ���=���܇a�eD�&� �=�R�      ���zg  ~��ѣ�/��:u�Z��7m" ���gϮ�       ���g��^f�a� @DD\����wOo���{DDf��y ���Z����w�s       ��`�� ���̬w�pǂ{��� 8(�k       x2���  ���N?ܱ�ۗ�.�s�����!       `��9s�Z�� ���Tp�%ubǿ�       �܋��C  ���^J�šF ��?�        ���;��������ꢛtUEIL�"(��yf�g��a�e�	K�^�0��#������cB@6�� �YT`�e�Q��FԤ;KwW���c��z��s�����oչ�O���|�I�RzZ� �[x� &���V:       &Q�۽OD<�t �ORJ���8q�#� �j~~~�q�#       `�|�=��  �ɚ�]v�Mq�H� �5�9?�t       L����J7  �b�s���pʁ�I_M �N����m�#       `�,..^�RzH� �[|e�Ν'N����SJ_Y ��n߾��#       `����<#"R� �[�p�/����~ (#����       0a�Y:  �V9�/��k��眿0� `#�����]JG       �$�t:??Z� ��?�N;pO)��C @1ۖ���R:       &AJ��� �Bgڪ�v�^U��; ����       gW�u�RzF� �;�/��k���t�M�� ��z��KG       @������8�t pJk�����#�+#� 6��9���       �f9g! Z(�t�}��z���v��s>�2 (�9�       ����O.� |����SJ�t_?��=�d� ��n����       �F۷obD|W� ��θQ?���l �zv�        h��ҳJ7  ��s��~Ɓ��> ��Rz��C�fKw       @�t:�{F�ϔ�  N-������a ��{�|��O(       mRU�s#q �^���8q⯇� SJ���       �-r�)"�W� 8��`pƍ��_~�?D�ׇZ ��8p��JG       @�z�GF�E�; ��:~뭷�p�o8�����wH1 ��m���٥#       �r��: ��_�u�|�oX���sC� F ����b       6����s��zj� ������Y�9gw h��v�?]:       J:q�Ŀ�9�S� 8���Y��g��� �����W�       J�9?�t pV�}ff�� ��鋋�w)       %t�����(� �Y�y���n����<�" `T�<�^:       JH)�B� ��2p���xD�0�" `dr�/(�        �v�����xN� ��q߾}_;�7�u��s���{ �{`��yD�       ��o����]�; ��Z�&}U����; L���..�        c�� ��[��� 0]�������#       `:��#r�.� ��gW�M�����|fc- ��l=~���KG       �8�K� 0QV�I_��}yy�� &DJ��Çϔ�       �Qj��n�� ��䜇7p��+�_�P 09���~�t       ����m�# �U���/��j�qU��>�� `�RJ�       S���*"~�t �j�ݱc��j�q���Ҫ�� Z�g���}JG       �(���?!"�{q �k٢�z��s��; L��+�       L��`��� ���^U��Z_ P��<xp�t       Ӂ~(���� ��������`�����o���#       `�fffvGD*� �^UU�ޢ�z�w�ޯG���U �s�ź�W���       �f�~��#♥; �59v�ȑ/����:x[��� @+\4??���       0���?E��� ��|�����~��)�O�� ()�|I�       بC��F�ť; �5��Z�yM��� Z�ѽ^�A�#       `#�9�8�t �6kݠ����\[ �9��       �A/.  ��Z7�k��OF�`ME @<���ܳt       �G�4����(� �]UU���۷���� �6�:33��t       �Ӯ� �����ݻ����i��s^ӂ h����u]o+�       k������t �.kޞ�y��R2p��t����疎       ���"b�t �.���y��X� �����-�#       `5���{D�sJw  �s��Z?����̌�; L����J�       X����]��t �>)�5o��<p��K�&"n^�� �v�9_�sN�;       �L�����9�,� �� ����~h���RN)���x �5���W:       ��رcGo&��    IDAT�]Jw  ���}��ݲ��y�1��T< �*�K       ��,--mM)�b� `C>���k��X�� �v��n�a�#       �TN�8�܈�W� `�r��ڜ�k��RZך h�����       ��><�s�S� ؘ�n��5p?z��'#��z> �Ɠ�����       pG7�p�S"�� ��������Għ��Y �5����       �F�9UUui� `þ�w�ޯ����G���x �U���v�S:       ""�����\� ذ�������:�� Ze6"��;       ��s�/� ��X��|���`�w �)��5MsA�       6�^������� �ƥ�ֽ5_����[n���X^���֘��}�#       ���(  �����i#7M�x�F�  Z������.�����t       �O�4���w��  ��{���z?���OZ�� h��[�l�;       ��R�  `h6�1����c�< �9�_X\\�W�       6��i/� �G7���SJ� h�m+++^q      `�RJ��t 0<ݘoh�~�ȑ�Gĉ�� ���^q      `\z�ޣsΏ,� ���L��{]׷Għ6r �*�VVVv��       `s�9�R� `xRJ7^r�%_���GD�?��3 �VyQ�߿w�       �[��y\D<�t 0<�ؖox�zB h�;�KKG       0ݪ���� ������ 8���n�>�#       �N�n��D�CKw  �Պ�/���OG�э� �ʝRJ��t       ӧ��*��˥; ��lݺ��=d��;v���>��s ��������/      �t���{fD<�t 0t�]XX�y��lx�1����֙YYY�KG       0=:4^o��4�M�P�)��� �u����~�t       ��ȑ#Ϗ����  �/���㜡ܫ���a� �N�9�j�       &_]��"�%�; ����a2����]��_�Y @��\�4�*      �d���QD�W� �[�9��a4���I^q�)�Rzi�       &����r��Jw  #󑺮��q�0�CyR h���#;���Jw       0�n��}q�� �h���lXgm��R��� ڧ��n]����8       6����{EĞ� �H�����fgg?ǆu �:���{v�       &�������; ��ɳ��>�Æ6p_XX8��y @+�Z]�甎       `2,..�?"�[� ��ZXX��a6��{DD�yhO� �tﹹ���       L����&"���  F���<l����P� �V����޽t       ���v���Jw  �5��P�+++^p��7_U�KJG       �^9�RjJw  �7�;p���K��R�q�g �s����\T�      �v��z�."R� ��/���O����#"r�2�3�֙����JG       �>u]o��N 6����رce�g}��R�а� Z�i�^��#       h��������t 0zUU���������� 6��s�sN�;       h����e����  �#�����޽{?��� @+=���?�t       �u��:"�R� ��7�|�G�}���)�2�s����u}N�       �j��Gr�;Kw  �R�h]׷�ܡ�#"RJŹ @�䜿~~~W�       ��G�l� `<r�#ٌ�d�>�`s���/����       ���i��/� �O���Gq�H��{��#�Q� �O���-[���t       �W���"�S� ����̇Gq�H�;w�<>����zV�4?]:      �񚛛���  ��S�w���Q<��{DD��C�: h�W�u=��/       h�����qy� `�F�� ���l ��2??���       ������#��� �x��&o�~�-��YD�� @;�;KKK��      �)��t�)� �]����������[SJ�� @k����㗖�       `trΩ��_�n� ����%�\��Q>�.���Gy> �Z��t       �����]D�t� �����Q���G|> �Nۖ����       `����΍�N� ���>�>ҁ�֭[?��� ��RJ?����X�      ��:~��K#��Jw  E����`�����c�g�� h���v��KG       0�~��E�ť; �b�r�޽_�#���1� �P���#���       l\]��`08[J�  e��F���}0��&�R��4���       `c�o����xX� �����z���� ����Q:      �����ߝRzY� ����Ǐhԗ�|�^������ Z�1�nwG�       �'�܉����  �I)���_���g���F�= �n)����Kw       �6�~�'s���t PV����g,����� �ڽgff~�t       �w����`p(���* �^�3p?��>?�� �V��^����       ��7������ @q�WU���h,�;v��?0�� �Vےs�o9�T:      �3����N)�J� ��d��ݷ�㢱�٘���7�� �V��i�c�       �l0���8�t �
��Ec����3�� �vK)u����Kw       pj�^�)�� @;TU5}�ݻw�uD�͸� Z���U�#       �NKKK���t ��p�y�}b\��m��R�r h��6M��      Z����݈�W��oz�;V�u�X���� ���\\\�K�       ���i?_� h�����y�X�'N�x_D�y' �j�ZYYyi�       "�����+"R� �=��z�X��eW\q�7RJ�s�w �wq��yD�      ���رc/I)ݿt �*_صk��y�X�9�?�� @�UUU���N�C       6��i~8���t �:׍�����}' �z�����t      �fT�u�RzUDl-� �K�y���{�D�M� h���K��;      �1���{a���; �ֹ��[n���/��}�Ν'RJ��� @�m����'       �U�4Dį��  Z�u]�:�KKȮ/t/ �b9�Gn߾�E�;       6��sJ)�""�K�  �s��Ľ��E�a������N�sQ�      �i����S��q�; �v�9_W��"�={�|)">S�n ��r��TUuu]ץ~      `�-..^�s>P� h���߿��%..6�9���� @�=|���/*      0�r�i0����- @;圯-uwɁ���� گ��+;��E�;       �M�׻8���� @�]W��b�m۶�QD-u? �n9�s������b?�       L����#��; �V�e�֭*uy�����±���R� ��۷oQ�      �i�sN+++�����- @����ֻ��/�^[�~ �媪����\T�      `����D�cKw  �w]�ˋ�SJ\� h���9UU]]�u�_�      �X���术,� �����K�_t(�gϞ/E�'K6  ��۷oQ�      �I�sN+++�����- @���e�]vcɀ6����� @�UUue�����       ��i�G�cKw  �R��tC�{J�J7  �s>'���C�͖n      �����O)��t 0r�זn(>p?r�ȟE��Jw  �!7�|�KJG       L�C�ͮ���6"�\� �7����tD�{]׃��Kw  �!���^��S�;       ���ѣ�?Q� ��޹s����UU��t 01��_�����!       m��t�s�[� �(ו�h��}vv���8^� �����[:      ��<8WU��1S� ��-[���tDDK�7GćJw  �#��������       ms뭷�����  &��.�䒯���h��=""���� �dI)�rii�{Kw       �E�4OJ)=�t 0q~�t�7�f�e˖k""��  &�=�?���       mp����� X���~�t�7�f�k׮/F��,� L�'v��痎       ()眪�zeD|O� `����ݻ?]:�Z3p��H)�f� L��үw:��Jw       ��4�SJO(� L��������^� �H۫�zm]�[J�       �[��@UUJw  ����V=Rު��ɧ�?W� �H������       �T����`�Ɯ�9�[ ����]�v}�t��j��R��t 0�.�v��)      0.���K��� ��z{J)�������A��� &J�Rz}�ӹg�      �Qk��9�/� L��R�ۭ��ݻ�#�� �ĺGJ�59�T:      `Tz���q�t 0Ѿq�ȑ���v����rJ��; �ɕR��^�wI�      �Q��zK����ݥ[ �������KG|���#"�A랺 &΁n����       �6??�҈xx� `���Z��n����.����z� `�ͦ�ް��tn�      �a��z�<缷t 0�9r佥#N���;v�D�;Kw  �ǏE�      �a�v�w�9�!"fJ�  �꺾�tĩ�r��sn�� ��yz��{N�      ���9���oGĽJ�  �/��ڭvk�[�n�È8R� �|9��l��Kw       �W�����t 0����^W:�tZ;p_XX8�� �(�#�u]o+      �V�^�"�WKw  S�=7��8���#"rέ}� �8?>??�T:      `-����s�o��;�n �CJ���V��9�wE��; ��s��^����       �Q�uUU��DĽK�  Scevv���#Τ�����G#�}�; ��s��N��Jw       ��������Jw  S�CW:�LZ=p���9��	| `�l������ҹ�C       N���=:�tE� `�L�6�����;"b�t 0U.:~��+KG       �J��;?��战)� L����rM鈳i��}�޽_��?.� L�MӼ�t      ��u}���["�n�[ ����.����g����Io)  L�^��yD�      �o���k"⡥; ������1)��q�t 0uf��zS�4^>       ��v�;"�_� FaPU�[KG��D���������Jw  S���x��ÇgJ�       �W�ӹ(���� �����ݻ�\:b5&b�QU�D<� L���x㍗��       6�n������GĹ�[ ��s~s�՚������5q[� `j�M�<�t      ����^?Z� �Z'N�8����51�����#�Jw  Sk&"~���ܷt      �yt��}�� �T{�W\���51���T:  �jw�����nw{�      `��z�G��^V� �z������ѣG����Jw  S�)���S�      `z5MsA�����t 0�RJ����w~g鎵���{]׷G�5�; ����i���       �S�߿sJ��q��- �t�9��_�£�;�b��'M�� �dJ)��i��-�      L��s��9?�t 0�RJ������ѣG�_-� L�*"���t�[:      ��^o_D<�t �)�������#�j��u]/G�[Kw  ��]��z{���^:      �|�n�1�� ��Rz���±�k5q����`0qO� �)���S�      `r-..^�RzSD̔n 6���\O��}߾}_,� lOn�fo�      `2���;��E��J�  ��ߞ��,�9pO)�8\� �<RJ/o��gKw       �%���kr�.� l*oٱc�J���ȁ{D�`0��'���UE������J�       ����$"�^� �\RJo,ݰ^�t�F4M����� ���'N<���/���!      @�5M��xKL�C� �D�aϞ=�I)��!�1�?8�n�  `������߭�zK�      ��z�ޏG��b�7Z ��I)�qR�����`0xCDL�� ��z���\�t      �N�N�9�wD���- ��RzS醍������?�s�X� `Szq�4/(      �K]�۪��&"�/� l>9���{��O��؈��GDTU5ѿa  L�_�v��)      �C�9���]-� lN)�חnب����̼!"�Kw  �Җ������J�       �5M����� ��5H)�N鈍����%�\�՜���  6�s���7Ms��!      @9�^�))�_*� lj�ٳgϗJGl���#"RJ�)�  lj?o���N�C      ���t:���ED*� l^9�K7�T܏=����� ��������,      ����⽪�zG����- ��v����;JG�T��>�Rzs� `s�9?�i���       ƣ��n�J�  �ޛv��}[�a���{D����kJ7  DD����\�      `�><�Rz}����[  ����-����������� ��������n���C      �ѹ��#�I�;  "�3�w��H�a����I�-  �s>'�t���Ⅵ[      ��k�fD��t @DD�����4U���"�D� �������W^y�]K�       �����W��  8iy˖-�/1LS5p߷o��RJז�  ��H)�vv�������[      ���t:��9�.�lw L�w�ڵ������Akڞ� &ޣ�?�ڜs*      �_�߿_J�m��t �7���.�0lS7p?z��"�oKw  ���{��KKG       ��4����u)��-� pߘ��}W�a���{]����  �抦i^P:      X�~��xgDܯt ���ް��p�tǰM��=""����  ������X:      X�Ç��7F�O�n 8��K��T���������Kw  |���xS�����!      ���x㍋��  ���={�|�t�(L��="b0��t ���9�3�i���-      ��u��}���  ��s~u�Q�ځ����#�X� �S�WD����޽t      �z�޳RJJw  �Ɖ�[���tĨL��}����,� p���u�����!      �?�v�?�s~MD��-  ��Rz����ߕ����GD䜯.�  p?q�m�]�����t      ��v�R�݈�R� ��.0JS=p��[������  8�G?~�꺮���2      h�~����ҵ��t �|mnn���4�C����#���;  �����#      `�Z\\�p0\�]� �,^�s���#Fi������Kw  �I�y�i��\�      6��i�r]Dܻt �Y��`����6�����>"�_� `~�i���      �����������-  g�Rz������tǨM�����*  �JW�z����      �iW���fff�)� �9�C��aS܏=zMD|�t �*T9��7M���!      0�꺮���~'"_� `������;KG�æ��u��.� �Jw���v:��     �i477׏��;  ���;w�<Q:b6��="byy���R� `�έ���~���!      0M��������  k�����ۥ#�e��/��#��  kp��`�����K�      �4�v��D�/��  X�?8���6��=""�t�t ���������{�     �I�4�RJ��  k��6Лj�~�ȑ�k�)    IDATk#⋥;  ��~+++�ꪫ�Q:      &Q��{ND�FD��-  k�R����Ͽ�t�8m��{]׃�ҫJw  ��-//_�W޵t      L��i��s���d[) `:��رc�t�8m��VVV~;"N��  X����^{�����!      0	��y|D�1"��n X�+++W���M7p߿��F�5�;  ��n��w�u��t      �Y��{t������-  ��{�^z�WJG�ۦ�GD���n  ؀1??����%�G      �B��}X�����p 0�rΛr�J��sN�^��[  �+��{G��Q��r�      h�N��cUU�?"�Z� `�zϞ=?�RʥC�m������ L��󿙛�{u]כ�g:      �v�~��UU��0n &\J�o�q{�&�GDTU��ҭ�;  6��sss��9oʿ�      ���t.�G���n ؠc����S:��M;pߵk�?����  ��5MӔ�      �R������zDܫt �^XX����lځ{DDUU�J7  CJiw�4��      0n�����D�y�[  �!��[�JJ�Jk�����;  �dq�޽�KG      �8,..^���򁈸�t ����޽{T:��M���I���ٻ�/�����O�ܐLO�FQ�$�"
."����*G����u�kV/Qp����$HB2=���Cý�������g/P���\�u�W�EDP =q����\?]�I�$�������<�ӧN�W�?�  g�A��     ��;��666~;���v9��m��w��uCD�fw  �EG��(;      6�����:��oF�C�[  ΢�;���ڶ�8p�ֈxsv ��TJ��     @5Ms�����.� -Sk}ݝ��mm��#":��JDL�;  β���h�      gK�4Fć¸ h��;v\�1�#���}""ޗ� p��RzF�      ��q; �f���<x�ϳ;�����j��d7  l#w      f�q; �v�[�;��i�4��"�;�;  6C�ui~~���      ��q; ���`0�a���_���  ���;      �fyy����a� �X)e)�a����N���� ��RJ�5M���      �j����icc�7#��� �M�׫����1M���^�w��z<� `�]�4͡�      �+M�|�d2�@D|sv �f���z8ޞ�1Mܿ�d2�>"ֲ;  6�Ѧi~>;      �����y��߈�Gg�  l��Z�k�#�����XXX��R�;�;  6Y��W�F���     ����t����{J)�"� `��СC�1mܿ�Z�Rv ��R�2�$;      �?�s2�����n �
�N�U�����+�����  �;k��h��_g�      �}�Z����k#�G�[  ��o�z�?Ȏ�F�w��rMv �9'"��cǎ}Wv      �����RD<'� `�*�������Έ�%� `��WJ�OM�|[v      ��x<���zqv ���.xOvĴ2p���p="���  �*�����6Msav      �C�4/����  �b��۷o#;bZ�ߍӧO��۲;  ��C#�W_}��g�      �nM�<;"��;  ���n����if�~7�9�Z��  [�[���?p�UW= ;     �v�F�>"�%� `+�R�|����gwL3��b2�,GD��  �b߱s��_�F{�C      h��h�C���GD7� `��Z�u������XXX�xD| �  �J)7?~|gv      �p�ر��t:��-  	�7�4;b����k�  ����'O����iH      ����Gu:���Z��n Hb�|��@��4M�ǥ�Ge�  d(�\���/��      `6-..>����ND\�� ��c�~�q���2�\p?w~�F�  Yj�GF�с�      f����y�n��ø ��J)W���3t�y��PJ�9�  K)ey<?3�     ��q���kkk��n H�竫��̎��gh����k�+�  �:����yRv      ӯ�Zn����G�S�[  �����zvĬ0p�j�������  Ht��x����C      �n��x���3�  ������bv�,1p����o�s� ��=pcc�����     `:���D�|v �����ʎ�%���JD�� ��C��������     �t�����zmv ��mmm�xvĬ1p����������� �)𘍍�w�����     `:4M�k�7FD7� `
��K.���Yc�~�"b=; `
<ymm������J     �m�i�GGĻ#�~�-  S�����Jv�,2D�����""ޑ� 0%~b�޽WfG      �gqq�!�x@v �������7gG�"�{��r4"jv �4��.4M��      �����y�n��#��� �)Q;��8;bV��K�~�c��fw  L���i��     ��������ߙ� 0-J)���z��1����d���  0E:q�x<���      �ƞ={V"���  S�Xv�,3p�����sD�^v �9����G�� ;     ���4��R��� �)�[�~�w�#f���}TJi�  ��7�ر�7�=�5�!      l��i����  �6����Yg�~����j��O�;  �̣���/���!      �]ǎ���xK� |�?��z��1�|ɼ����$"��;  �M)��sss^�     h���Ňt:��DĞ� �iSJ9VJ������,ؽ{�["�/�;  ��K���E�      �w�]w�\��}_D<4� `
�277wcvD����ֺ�� 0�j�׌����      �����o����xlv �4��6���?����g��ݻ_���  �B�Z�ۖ���     ���w��q���ew  L��=��sߘ��gɁn-���  �R{'��{F�у�C      �g��y~���� �)v�E]t2;�-�ϢZk>�  _�7�R~m8��     ��9v��S#��� �)��n����&�g�`0�l����  S�����\k-�!      ܽ���Gu:�#bGv ��*�,<x���mb�~��ZG�����  �b�g�4/ˎ      �]y����xoD�?� `�ݺ���z�Yf�~�:t�"�w ��QJ���h�ew      ��VVVv�ڵ��� �iVk��ȑ#���h�M������;  �X)��aii�{�C      �b�O��6"��� 0�n�v�WgG����&����;  ���&�ɻ�     ��k��ŵ��ew  L�Z뵽^�o�;���}�t�ݫ�w ���������     �yRD4�  3���ݻ�Ɏh+�Mr���OEě�;  f����^�     ��5Msa��]�+� `ڕR�=p��g�;���}�R�F��  3�9��xv     �v���tND����u�-  3ඝ;w.gG����&�����+�  g��z�����gw      l'��2�L���n ���W�޾��7����U��� 0vN&������!      ��x<^�����  ��M&��숶3p�d������  3��k����f�      �ݱcǞWdw  ̊Z�����:���ܷ��ӧ�W� ������^�     �f�����N�ƈ�f�  ̈�w���z�0p�w^q��� ��S��     �F���{k��g�  ̊Z���Tv�v`�Ej������  ���z�i���      h��p��v�o��o�n �!�O&�qv�va�E��M��� �ҍ��.--=";     �-���^�Gv �,)��faa�/�;��-��t^��  3����W���     �Y�4�3"��� �s����(;b;1p�B�^��ַew  ̘~�ԩ7dG      ̲�x�ȈxSD�� ��:�۷����v��W� �}MӼ$;     `�F�=��wE�y�-  3掍��c�ۍ����z����;  fШi�'eG      ̚R����� �YSJy��������n��R.W� ���h���     �Y1�/�����  �A�J)G�#�#��~��"���  3补�_>q�D7;     `�---}O�u�� 0�J)W�z�OfwlG�I:��0"New  ̠'�t�M/ώ      �fKKK�L&7F��� ��RJ��]�'��z�,���  �E��K�����     �i4;o���e�  ̨c�^�o�#�+�D��WF�jv �*�����g�      L������R��� 0�j����ظ6�c;3pO4>[k�:� `F=`cc�]KKK�d�      L��h�Cqiv ��*��baa��D��&�ɨ���� ���Z�5�      ���ѣ�R��� �uӮ]�^����'���� �YUk}�h4���     �L+++�w������ �YUk}�������ܧ�m��vmD��� �YUJ��رcߕ�     �emm����� ��g��v�/eG`�>������� �v�N�s������C      �Z�4?���  �q�����ܧ�޽{��3� `�=bcc��      [iyy�Q�� ���~���������ؿ��xYv ��{�x<�(;     `+���mll�-"�d�  ̸KK)5;��g�>EN�<����Xv �,�������;      6����rD|gv ����`0xv������Z�+�  ���Z덋��{�C      6�x<~fD<?� `�u:�˲�b�Sf~~�=��  3�[���Jv     �f����Z_�� �����>��3p�N��  Z�9M��tv     ��4w�Z9"�� 0�j)��|9�)4~+"~3� ��o��۲#      Ζ�{�^O��  h����fG��ܧT��95� `��Eĉ�px��     ��j<?��:�� �����2�)��������� �x������     ��b4=������ ��J)o���W��[__?��  -p�i�ˎ      �7��a���ֈ��� �8�Ȏ��O�����G��  -P"�������     �{jnn�pD�Pv @K,���[�#�k�S���\�ew  ���"���pGv     ��ZZZ���fw  �A��3���ǲ;�{�S���}�ֺ�� ����gϞ_��      8�����L&7F��� �6(�>�����L&���tv @�R.��O��      �j&��#�a�  -��{��.;����},,,��R^�� ��Z�/---=0;     �4M��Z���  h�Rʡ�������3p����#�gw  ��7M&��     ������#b)� �-j����������ψ}��m�Zgw  ��3���#      ���p�cccㆈ؛� �����#8s�3d~~��#��  mQk}����ò;      ��޽{/��'dw  ���^��#8s�3��2�� �������_:q�D7;     �i���Z/��  h��#���3�3���,"~)� �E�t�M7y�
     H5��D��"bgv @[�R���M��3�3���\ZJ��� ��(���i����      ��N�����  h�Z�gN�>����=g�>�z��''��rv @�쬵�����9�!     ���4��Z��� �&�N���Bv�����:��s�F�_ew  �E)�Q��įv    �-����u�(�-  -�񹹹�fGp��Ϩ�.��dD�<� �e^4�$;     �j�emm����-  mRJ9������;�3�.x]D�qv @��Z�F�у�C     ��[ZZz~D�hv @��Z?���ߛ���g�>���۷QJ9�� �2.�ώ      �mii���c�  -S��� ;����}����_�����  h��F?�     ��p8�1�Ln���� �6�������Av���{L&����dw  �I)����ew      �gϞ�"�_fw  ���˲#���[�СC�o���� ��ٻ����Zk�     ��رc�YJ�$� ���7eGp���D�۽���w�  -�䥥�fG      �0wu:�_����-  mRk������������z���.ew  �M������ó;     ��777�҈��� ��)�\r���/dwpv��H�ӹ2"<�  pv�M&���Cߝ    �{m<?."�;  Z�/���7eGp��H��;G�;  ڦ��}sssew      �i8�bD��n h�:�L^�o߾�����o��~8� �mJ)G�;�-�     �왛�{YD<&� ��n8t��ogGpv��Ӌ"b=; �Mj��v:�7�8q���     ̎�x������  h����#8��[h~~���Z_�� �BO���_�     ̆���ݵַD��� �z����_fGp���T�۽,">�� �6��+���#�;     �鷶�6���� �B�s׮]��l����z[Jfw  �M���Z�O�8��n     �ױcǾ+"��  mTJ����wdw�9�[����MD|,� ���p�-��$;     �N+++�;��["bgv @}����Zv�������۷/���� �6��+��ytv     0}���.��o��  h�����gG���[n0|$"~%� ��vG�N�8��     ��h4�����  h�k>���2p�����K)�� �B�{��7Ȏ      ��p8�UJyCD8� p�}z}}��l>�m����7�Z�;  ڨ�r����ó;     �|{��=ߞ� �F��Ç�Bv���}��t:����� ��������~]v     �kqq�[k���;  Z꣫��oɎ`k�o�^�T)e>� ��J)O�����      r��N��}}D�/� ��j����p8�ak�o#�~����� �6��^=���     l��{�� "��� �Ro����/�l����#  Z�A1Ύ      �����Cj�Wdw  ��j�۽4;��e�����gw  �Q)�Y���G�;     ���cǎ�#���  -��~*;��e�u��a��3�  mTk}�u�]7��     l��h�����;  Z��v�zUv[��}:x���K)�ew  �ԅ�N��<;     �\W]u�J)�dw  �؋8pGv[��}�:y���#�fw  �ԁ�i�;;     �<;w�l"��;  Z��`0xv9ܷ��p8��D�Fv @u#�Ǐߙ     �}���"�g�;  Zj�����#�cྍ���R���  h���z뭃�     ��ZZZ:���(�-  -��^������os���E�?  �������Gew      gO��e�� ���o'O�t�y�3p��Vk��q  �����_]ku�     Z`<?�����  h�I��y�p8\�!��;1??����� �6*�|�4���      ��pة�^;�[  Z�5�^���#�g�NDDt�ݗD���  mTJ5M��     ��777����  -��ӧO_��t0p'""z��'"�� ��zP����     �޹��+���  h���#G>��t0p��<y�hD�iv @�R�7����     �s�v�G��Z 6A����~�m�Lw��p8\�t:Ϗ��� �B�R���p�#;     8sM�<)"~&� ���J)�/�خ���"�^�å��gw  {+�    IDAT��c������     ���y��UQ�[  Z��`0������;_����"���  mTJy����C�;     ��nϞ=#��  -���'O^���1p��\|�ş.�\�� �R�u��&;     �{����R�/dw  �U)�%��������;_����#���;  Z�'���fG      w��zuD�ew  �ԍ�~�}�L'w���p8���� �6���zeeewv     �嚦yZD<#� ��n�t:�����;wi~~���R���  h�o9}�� ;     �bw�Y��  h��z��'�#�^�ܭ����"� �MPk�tyy���     ��v�w\���  h��^p��/s�ܹ[���@  l�s��ׯˎ      �����#J)��  -5)��h߾}�!L7w��~�c��}�  mTJyz�4?��     DL&��#�~�  -��~��{�L?w�H��}ID���  h�奥�s�#     `;k���� ����������w�H���DD\�� �R�L&�;    �$���~�dw  �؋>���f��;g��ɓMD|4� ��7Msav     lGsss�"⛳;  Z���`���f��;gl8��R~."Ng�  ��9��     �����C#�Pv @K�͎;^��l1p������qv @K���h��     ��t��&"�dw  ����/�����w�]�vk��� �F��W���     �;v��"b_v @K��~�Cv����{���wD��E�$� ���}�޽�ˎ     ����N�sMD�� �����>��R�C�=��+������  h�Z�W^y僲;     ����ݻ?"�� �RG<����&w�]�v-D�-�  -��ݻw�#     ������Z/��  h��r�\���2p�^;p������gw  �Q�����;�;     ��v��uyD|mv @�u:��۷o�Fv��������/"ޞ� �B�R���     �6M�<�ֺ?� ��J)W�z�?��`��s6���Ύ  h�'���gfG     @��R�#bgv @�����bv�����l0|�����  h�Z��p8<7�     ڠi���>5� ��&����õ�f��;gE�߿!"ޛ� �B�����#     `�---��� �6��^���'��v0p�Y__qD�fw  �M)eaii雲;     `��Z{�� ����=�ܗeG��5����zIv @��ZϝL&���     �Y5�\k=�� �Bu2��袋Nf���U��v���� ���i�     3��8/; ���t�СdG�.�U��p����܈�=� �e:�dG     ��i���J)?�� �Bu���Av�c��Y�����R��  -����G�#     `��Z��#� �mJ)/:r���;hw6����bD�av @��Z��Ǐ���     �Y0����#�  -��~��������M1�#�yq:� �e�uuu�y�     0��a�ֺ�� �B�ݱc��#h/w6�`0�hD\�� �6���ѣG�&�     �ٞ={����  h�R�/���Ogw�^�l��'O�����  mRJ��;v��     �i���tN)���  -��~��+����;�j8��R��g�  ���M�\�     �h2��G���  -󩵵�gG�~�l��`�?j��gw  ���J)WfG     ���F��Av @��Z/��K�&���3pgK�v�m��� �6����h4zBv     L�R�+#bov @˼i~~�W�#�����p����܈8�� �"��2����     �M�<:"��� �2�<}�t?;�����-�����4� �e��4͏eG     ��X���  -R;��s�9���w��ɓ'������  h�R�����wfw     @��h�C�� ��9����Svۋ�;[j8Nj�ω��� �����՟ˎ     �,��RJ9�� �2���q(;������~��O{��>�&� �E���<�5��Og�     �V;���CD��  h�I��y�����e�����N�^���Z�'+  Ξo��    `�;j��� �6)���z�gw�=����R���s#�s�-  mQJ9t�W>(�     �����s#�۲;  Z�㥔K�#ؾ�I���>Yk�gw  ���w��u(;     �����9qiv @�L"⹽^�Tvۗ�;�����TJ��� �90��ώ     �����qqD<4� �E���dG�������\�� �����fG     �f[^^�)e�� ���?9y��˳;���t�TD�8� �-j��qyy�Q�     ��666�D��;  Zb�����px{v�3���#�W�;  Z����qyv     l���Ň�R^�� ���+����w��#���  -���x���     �����j��fw  �����]������1>���  h�Rk�";     ζ�x�Ȉ���  -q{��y����Og��?0pg��w�Rސ� �?�4�S�#     �l���2"vdw  �A)e����(��)w��d2yID|<� �%�����     8����ED<3� �%�����ώ�/e��ԙ�������LDx� �{���ҏgG     ��0�L���]  �Z�gv����RJ�n�/e��T��z��gw  �A����p�V     fZ�4O����  h�N��܋/������3�N�<yeD|(� ��w�ޟȎ     ����zEv @K����7;;Sk8NJ)?��n �u�֗��    ��j��)�����  h�O�s�9��pwܙj�~��Rʁ� �xĞ={~:;     �R�K�  Z�t�����.��dv�w�^�߿���� �YWJy�p8ܕ�     �D�4?\k�W�  �����^�������3N�>��)� `�]877���     ����  �����^xa��g����p���/Dĳ"b#� `�]����;;     ��x<���=�  3��֟޷o�&3����1>RJ9�� 0�ο�;��     _M���Z/��  h����#�Lu���x����]�v=-"�� 0�J)�{����}�C��[     ஜw�yό���  ���z������pO���L��N�Yq2� `�}������     �+��Sk}iv ���e}}�@v�S�̜^���R� � `��Z�\w�us�     ��ٳg_D<6� `�Mj�?s�ȑ�e��=e��L����#��  ����u�N�zav     |�'Nt#��;  fܕ���ʎ�{���Y����Tv �;����7;     ��[n��'K)���  �aݻw���po�3���g'��s"�f�  ̨�ر�@v     ��'Ntk��ew  ̰�666~j�����C��2pg�:t���k�;  fU�����r^v     DD�|��ϊ�o��  �U�փ������������� 0�������     8q�D7"�dw  ̪Z�;���_�����;3o8�^J��X�n �Q�뮻n.;    ����o��� �+�������gw��`�N+���?+�\�� 0�t�ԩ��     l_���� �[�'��O�z������� g�>��?|�S���"��-  3�O�ӯ{��߿�    ��s�y�=3"^�� 0����OdG���;�r�9�0"�4� `}�d2ynv     �S���v ���������:U]Y*pw� �>�F�#���b �Y��Ą- �@C�:�{���+KHwWUk�3y0����G7��AŇ���"�MY�>tU׹��s#f饪>gy>��ׯ�s��u���^o5;���;e߾}�N��'">�� 0������ʎ     `�����@D|Gv ��hD<��R�C`+�3q���j�K�  c��ʎ     `��� �k��h���C`��3�����J)���  C��m;�    �t8t�Г"�q�  㦔�����dw�v0pgbu:�gG��;  �I��a���7dw     0fff^��  0nj�o���n���b���Z\\�l�ӹ."ֳ[  �I)�Gڶ���     `�>|������  '��O�����ٳ���������v�Qk��� �1��w�S�#     �l���n  3���<{������T�`��Z�����#�� �qQk}�cǾ�m�av     �gee�j�o��  3�5Ms ;��ܙx��:77�����% ��TJy��ݻ���     `2�×d7  ��w�޽�ǲ#`'�3>��t����� �qQk}I۶�     �R����.�\�� 0F>{��ݻ�;�X����v����  #�:??iv     �e8�n  '���4Msgv�w��`0����  㢔�#�     L��~sD\�� 0.J)k�~�u���ܙ*m�gggo���g�  ���\^^���     L����~ث  ��w=ztv�4L��n���qcD�� �1�c    �3v�С���ސ� 0&���{ڶ�Bv�4w�R�4o���dw  ��K:���     ��N�Ӎ���;  �A�u����ߟ�ܙZ��-��  c��Rz�     ���n��A�� �qPk���~��; ��;Sk�޽�����Z?�� 0�J)�9r��     ��]�v�0"�� 0�lff�%tL5w�����?�E�fv �������fG     0~ڶ=����� �1�Z�U�n���!���������RJ��� �QWJy����Wew     0^�;�gG��fw  ��aD����?���!"����K)���  e��s�?���     ��w�1��  c��MӼ!;F��;DD)������� p?J)�<�;�    ���}hOD|cv ��{�����fG��0p�{8p�3����|v �������fG     0J)Mv �������u{�����Qa�_dii��J)�F ���n۶s�     ����Ջj��:� `�m���>�����D�׻="�Kv �������#     m��pv �(��v���~?�F��;܋�`�/"ޙ� 0��m���     �^-//?&"�� 0�~���*;F�A
܋�m?��t�����[  FQ)����fw     0���  ��������0���>t�ݿ*�<#"jv �(*�t�     =�������;  F� "�ZXX�;;F��;܏^����֕� �������fG     0ZJ)7E�lv ��zA�4������c��Zߚ� 0����Bv     �cmm��Z��  �����4��ew��3p�ж�]�v=5">�� 0���v�mˎ     `4?~|oD<(� `��ѣG��0��$�t�M/�\�-  #f�����#     �׶�l���1 �?�陙��ڶ]��q`�'����A��G�;  F�޵���#     �5??�����O �j�/..�Mv�w8M�,�Z�[v ��9}}���     r�R~8� `��i��ʎ�qb����R����� �sS۶��     �X]]�w��� �QRk���`pkv�w8E���?��t�Dı� ��ݻw?%;    ����n  1���xF۶��7�p���j�O���� 0*j���     v����7E�%�  #dPk���[n�Tv�#w8M�~�u��۲;  F�cVVV�    ���ݰA �G����~����W>.�=z����  ��C     ����ꗗR��� 0B^���^�����@۶ù���k���n ��+:��     ��p����  ����=��0���-,,�]J�&"�f�  ��������     �����Y�� ���'N<uϞ=��!0��a4M��֧G�0�  [����n��A�     l�����"�k�;  F��N�s��7�|WvLw�"�~����� ��{vv�Y�     l�}�  #��Rn�v����Ia�[��뵵���� 0^ض��    �	u�С�dw  �������28�-TJ����ƈ�O, `�}������     l�N��� �l�����gw��1p�-�������"��-  �J)7     &���Wew  ${����3۶f���1p�m����WD\��-  ��t�ȑGfG     ��:��"bWv @��gff�r��7ߕ����I�4�mv @�������     �����Y����  H4��^�������Tz��+"�� �,��g���~yv     [�����G��dw  $��~���0��a�R�9��xwv @�Z빵�gew     �e^�  ����^�����t�����7����,"�>�  C��Ew�q�Lv     g�СC�SJytv @�Z�{w����RJ�n�Ig�;`qq�o"����LN ����×fG     pf:�΋�  �|fff�򅅅��C`��i��M����  �Pku�    0�VWW�."���  H0�����_e���0p��4͡���� �O\]]���     N�p8|AD���  �i���MӼ!����;�RJ�t:ώ�?�n �ae8�0;    �S���vVD�Pv @����z��0m�a�u���onn^�n �aO�+_�e�     ���Ǐ__�� ��J)o���id�	�����R�eq,� `��ڵ�Y�     ��d  찿�״m�������z�?��gD�0� `���Z�#     89����-�<:� `�t:����Od���2p�DM��J)���  �A߸�����     N�p8|~v ��R��v����if�ɺ���#��;  vJ)�a    �x�+_�e��=�  ;���z�������R�`0���x{v ������͎     ���ڵ�ٵ�s�;  v�O7Ms$;0p��ж�fgg�RJ�Pv �����ynv     ���Z"�y�  ;����`��;�P������ʣj���e�  l��ݽ{����ݻ�    �?�����xcv ������w.,,|2;�np��������Ԉ��n �f�b0\�    ��+�<?� `�]k�ܸF��;��^������ ��Vku8    0�VVV.��^�� ��6k�����wg� ���;���in����� �͞������     �S���E�lv �6[������s�0�v����Z�[�;  ��=�$     ���o�}WD<;� `��T�4�!;�w�0���ݻ���quD| � `��Z�y�����     ��`0�*"�� ��~w0<?;�o�0�n��OE��qWv �6yPD\�    �?��^ �$�눸�m�����Èk��/:��u��� �J)��     �8r��#K)ߛ� �M��t:�7M���!��3p�1��v�XJY��  �&�:|��Ɏ     �v���Ϗ��� �ND�5�n�=�!�3p�1���Vk��gw  l�R�s�     �����9��� ��PJYh��M���1p�1r�ر����  [�����n��A�     �j8gw  l�Z�r�������3p�1Ҷ�����U��� ��Tk=wvv���    �i�M `B��c��gG ��������ݝN璈�Hv �ۛ     0������Z��;  ���g�m;�N��;��n����pxED�[  �пZ]]}lv�e`    IDAT    ��)�썈�� ��>Xk���m?��:wSKKK�3"�Dĉ� ��2=�    �����Ϊ�>-� `}jss��~��������k����dw  l������ώ     �����D�Wfw  l��Rʵ���vp��a������Z��;  ��y?�    0-j�^� &E-�<����vvpf�a4M�TJ��� ��Pk}~v    �4XYY��R��fw  l�Z�^������3p�	PJ�G�}N)���[  ���:���#     &�p8|nD�� �-������`k�Äh��Ǐ�""�Wv ���t:��    �Fm�ΕR��� p�j�o^
�	b��[n�������� �3����Ύ     �T���WF�Wgw  ��wonn^׶��`��ÄY\\��N�sY)�s�-  g�N��';    `R�R��	 ����R.��������;L�n���Z�3#b�� p��     l�Ç�ˈ��� �3p��rI���pv���aB5M�˵֛�;  ��w���<*;    `�t:��� 0�6"��^����!������.��*� �<;;     `��q�3�֧gw  ����iޔlw�p\p�M���gw  ��Z��������     �w�y�E��� ��Qk}Y�4�)��^�0���ٳy����#��-  ��ˏ?~Ev    ��1;  �4�R�4/Ɏ ���;L��m?733seDܙ� p�     l�����*�\�� p~g0<��R�C��g�Sbqq�o;�Υ��� �SQJ�pee��    �q���������  8E���ظ�m���`g���v�冀^ǲ[  N�LD<#;    `<3;  �}��rɁ>��w�2�~��J)�Eĉ� ��Uk}N��dw     ������Dģ�;  N��"��^����`g����z�ώ��� p���#G�7;    `\�Zo�n  8Y��ϕR.o��}�-��3p�)�4�ϕR~4� �d�C�/     ��m۳�y� `l���{��d� 9�a��z�WD�Ofw  ��k����ώ     7���WEėew  ��ZJy^��}v�����`0�F�k�;  N�������    �qSJ�B& 0j�z��Oew ��aʵm;O��7e�  ��0     �`yy���}�  '������#�|�@�m�>77wMD�iv �xܑ#G�    0.j�7�} 0���`0xQv0|� ���p���ܓ#�/�[  ����泲     �A���R��� � ~{nn�m��C��`��o��G�ǳ[  ��3o���]�     �nyy�����  ��]333W-,,�F��;�O,--} ".��Av �}�������    �1���  �����p������f� ����g����Z��_q �H�.    ��;|��|)��� �������/--�]v0z܁{����7F�0� �^\q뭷~Ev    ���t:�F�y�  _���Z�����v0�܁��4��SJY��  �ssss�fG     ��Z�3�  ��F)��~����`t����뽺ֺ�� p/��     0�n��EĿ��  �5"���vߘ�6w�5M��%� �K<����ߜ    0jv�����	 FO�i��Ɏ F����R��ݻ�o�n �b�N��    �QSk�& 0jV��YɎ ƃ�;pR��ݻ1�)��-� ��R�Ѷ��    �{���|WDx� %?�������0NZ۶���ظ���?�[  �������͎     no F�?TJ��!��0pN��7�|׮]�.���e�  DD�R�     DD۶s�'� �o�����m��!�x1pN����'777/��;�[  "bϫ_���#     ��޽������ ����s�9�)ǳC��c������d8^�� L��>���_�    0�x	 ��wnll\�o߾Av0�܁Ӷ������'G�g�[ ����    �j��z�W�Z/��  ��_��'8p��8m������,�\�m d�����͎     �277w}D�ew  S�#333.--�]v0�܁3���������8�� L�������     Yj���n  �W���q�����d� �����~�ͥ��G�fv 0��     S�ȑ#�,�<:� �Z���>�i��e� ����2�^ﵥ�gGD�n �ҷ���<*;    `��8q�� `:�R>7/_ZZ���`r�[����lD�pv 0�j�q    ��Rk-����  ��F�������e� ����rM����xiv 0�n��;f�#     v���꿉����  ��f)��MӼ!;�<���h��%��� L���y�ߓ    �S�l	 $�����z���L&w`��z�~)����  �K)�a    0ڶ���k�; ��RJY������ &��;�mJ)��.���n �ʞ���s�#     ������#⫳; ����^���L6w`[�ٳgs0<-"ސ� L������     �͋� �{u�4/Ɏ &��;��ڶ]הRޖ� L�:    �D;|��|D\�� L�Z�����`:�;�m�ϭ��_�� L�K�9���    ����t��ew  S�W�;vc۶��`:�;��������0"ޓ� L��O�8quv    �v�^� v�o���]߶��`z�;jaaᓵ�﫵�7� �l��;    �DZ[[��R��gw  �̓��ʅ����!�t1pv\������̅�� `����>4;    `����_�� ��*��~��ʶm���Lw E���h)�	��� `bufgg�ˎ     �^� ���O�8qq��?�L'w M���pD<!"��n &S��!    0Q:���� `b����ƥ���?�L/w U�4w��#�c�- �D��Ç[v    �V�t:7DD��  &ҟmll<��������;�nii�/#��Z�'�[ ��t]v     �zjv  0��?;;{�q;0
܁��4�_D��Għ�[ ��RJ��Z�ی    ��w�Сo��o��  &�_���<ᦛn�xv@��;0B���;����Għ�[ ����+++�Ύ     8S�N��� �V�3".\\\����d������?��^G�[ ����    ��f  �õ�'4Msgv�3pFN����R�E1�n &��m��    [+++�ߐ� L����'���f� |)`$�z�?���#�Xv 0r��~wv    ��R% �U>OZZZ�@v��1pFV�4�O��/d�  ���8�    �R۶�Z�� �D��Z��������b����i���t�ǳ[ ��Vk�Ӷ�lv    ������ވ��� `�}6".������?����v�o���`Dld�  㫔�U�{��ew     ��R�*�3uw��yr�4��@܁����_�Gĉ� `|u:�@    �X��eʫ�; ��UJ�\D\��vߑ�p2܁��4�/�R��� `l]���vVv    �ɺ�eʯ��  �ֱ�pxi�4��p�܁����~6"�G�[ �������'gG     ��N�s]v 0��_k}\������Sa����i~9"�n ��S�     N�=/R>%� ?��7�Z����3��T�c�i������n �K���Ç�gw     <��Ǐ_��  �ί;v�)�~�Xv��0p���������>1"ޟ� �����4;    ��t:�=� �����શm��p�܁�v�M7}|ff梈��� `|�R���     pVWWϩ�^�� ��R��:���m۞�n8���[\\��N����lv 06.Y[[;?;    �lnn^�ew  c�=�N��n�����3e�L�n�����."6�[ ��p������     ����\��  ��Ow:�+]
Lw`b4M�[�fw  㡔rmv    ��Y[[;���� �X،��u�ݿ��*��D��z���;�; ��Wk�xmm���    �/u���'E��/�TJYj��� [���(��z�9�<'"�2� yg���_�    p/��  �¯w��#� [���8���D���� ��Rʵ�     _���o�UJ�,� m��u:�g�Rjv�V3p&R�4\JyEv 0�j����y�    ������ `�m����C ���;0��=��Z�[�; ��v����/Ɏ     �G�֫� ��Vk��~������b�L��m��N���� `t�R��n     ��h�v6".��  FW)�m��W�; ���;0�z�އK){�; ��v������     �{��E�Wfw  #�Z����ٳ���܁����^[k��� `d�}���K�#     :���� �H{Q�4wfG l7w`*�u�Y�"�� �h*�\��     L�;�c&"���  FS)�uM��\v�N0p�����ݵ����� ��K����ώ     �ׇ?���G�Wgw  #��Rʋ�# v��;05���["��; ��t����/Ɏ     ��p8�:� Y�n������b�L����ň�Dv 0zJ)�f7     өm�N)��� `$�n��{Mv�N2p��-����fw  #��Ç�gG     ���������� ��9>33��K)5;`'�S�i�_��_��  F�9�N��    `��ë� ��SJy����{�; v��;0�N�8�dw  ���zUv    0]j�%"���  Fλ�;�C� f� 2���o��IOz�"���- �Hy����#��;�s";    �����]JY��  Fʰ�z����! ��L��`���� `��7??av    0=:���� ����~�o�L-w`j�m;�t:{#b#� ����    ��Pk-�7I �+�|�s�����L��T�v��*��fw  #���o�}Wv    0������  Fʋ���7Ȏ �d�L���>����� `d|�ѣG�    L�R��� �Hys������l���۷oߠ�rsv 0:j��    ��pUv  026"�E� ��� "���/�Rޖ� ��Rʕw�q�Lv    0�����#"�!� �֟l��}� ��� "J)5"~8"6�[ ���5�Ї�;;    �\�/I ��㛛�/ώ � ���zZJ��� `dx    �6�V�A QJ���o�+�`T�|��Ǐ��Oew  #��ZkɎ     &���ʣ"⛳; ���'G�����Qb��En��OE�˲; ����#G�<&;    �<����� `$k��ڶf� �w�/1^���  �y"    �&�d  �J)?����(�`��|��mO�Zo��  ��Z��n     &����R�� ��kff�G�# F��;�����o��_��  �}������    L�R�S� ����7�t�ǳ# F��;�}��6��  �p8�"�    ���˳ �t�۽{���# F��;�}���,��dv ���j�    l��>$"�� �*��߻w�Fv��2p��N綈�Tv ����+++dw     �ovv���(� @�?�v���0�������gK)�fw  �JDx2    8c^� ��aSJ�� ����=z�U��  �C'    �L����O��  R������gG �:w�ж�zD�$� H��#G�<8;    _Ǐ�$"�; �4�333/Ύ � '����bD�Iv �f������    ��*�x) ��kߛ0�NB)��R�� @*�O    �i����wE�E� @�c333/͎ � '����v)����  �\���vVv    0~��'Dă�; �4+����0.�N�p8�G�0� H�{}}���    ���t:^��)Uk�����Jv�81p8�~����_��  r�ZB    ���Z"��  G���񅅅��; Ɖ�;�)*��8"��� �R��F    ��#G�|GD\�� ���G��&;`�����iWgw  )������    `|�C/C��*��ܶ�zv��1p8���Ogw  ;���0
    8�g  )���v9;`���|�ֺ�� �Rʕ�    �x8r��#"�_ew  )^\J�� ������E�'�# ���+++ߔ    ���pxUv ��J)��4͛�; ƕ�;�i������ ө�zYv    0�j�Wd7  )~4; `�������WE�ǲ; ��UJq(    ܯ[o��+"�q� ����^���� ����t����Zgw  ;����?�?�5�    ��:묳.���� `gu:�g7 �;w�3t�ر���  vTgss���    `t�Z�	 ��M�n��� �����m��R�m� ��r8    ܗ���s"��� `g�×e7 Lw�-p����D��; �u��Ç�#    ��Sk�0"�~ S����KKKo�� �� [�m���p�; L�sJ)n`    �/@���������Ia��Ev������� ��rH    �m�v"�� `G�j��}Gv��0p�"{��ݨ��<� �Q��m;�    ����;�q�� ���a3�������🍈�gw  ;�+�9�    ���Z��`���i�?Ύ �$� [hϞ=�����)�
    �b��˳ �SK)/͎ �4� [��ѣ����  vF)��    `4,//KD|Sv �c���z�0i��X۶�Z�[�`z<����ߖ    �����F������;�6h����� `g�R��n����{{����;�]{�$���<I �@[�c�ql��#!m���_Нk�����ԧ��f�S\�pHB�8$�@��!�$���<q�� %�Ȓlyf�Ջ��H������{�^��r�>{-    Z�?e  #��C�});`�A)�F�]� �h�Z�cv    ��رc?o��  F����;�# &��;��\v�eG�; ��+�\s���gw     yz��[� ������Ɏ �T����{��"��� `$J��sv    ��-� �h���۳ &��;�mݺ���; ��px    Sjiii[D�lv 0���?�0���h���gJ)G�; �����i��    �������+� �N���v�!3p�~�o���dw  C�c�Ν7eG     �Wk��# L��8p�� ���`����Nu:�_��  F�!    L�Z뛳 ���ϥ��0��F`yyy)"���  ��?d     �u���+#�� ��}��ɓʎ �� #����݈x{v 0t�9r��    `tz�ޯd7  #q{�4���i`�0"��c���� ��9�   �)��tޒ�  ��O�<��� ���`D������ ��,    ���~���Z���  ���rg�4�ew Lw�ZYYY���d����n{Av    0|333o���� `��YJ����ib�0B�~���[� �Pu�n���    ��u:/:�������}&�`���X�׻="V�; ��r�    �����Z�/fw  C��^�����ic�0b���_��dw  C��i<K    ����>"^�� կ.,,|7;`��$���5� ��o߾���    `xJ)���  �3[�n}[v�42pH077�W��?��  ����%�    �Z�d7  C���������id�����ݝ�  O���    &ԑ#G.��+�; Ŀ+�    IDAT����nw);`Z�$�������|v 04�^\\���    `(�Cv  0<���8p��� ��� ��  ��-�    0�|��	�����n �f� �v���ވx"� �\    0awD�M� �p�Z�r~~����if��h߾}�qOv 0����瞝�    ���R~>"��� G��9�� 0���-//�'�; ���v���͎     �ˍ 0���駟�`v��3pHv뭷~���� �pt:�]    0!j�%"ޜ� ͯ6M��0��Z�����������    �1w�رk"��� �P�XYYqI%@���������  ����Ύ     6����F �P��������� ��d1;  �N��+�    �����Z��z����g������x(� 
�^    0�_�dw  Cq|aa��� �?w�v�;;  �7�u�]?�    lʿ; �T�� ����EN�<������ `�:��7gG     ��t�� ��C��Ev ?`��"M��#�ײ; ��p�    c�i���֟��  ��zwv g3ph��'O�+"��� V)�����ew     �}��=�+� ���:u��# 8��;@�4Ms:"ޞ� ��3g�ܘ    �_����� `(�6M�ώ �l� -����; ��*�8   ���� L��<y�# 8��;@������� `�j����     �����OFĿ��  �MӜΎ �\� -���ߖ�  V)姎;���    `]ޒ  \����� Vg��Rsss�� V�����    `]ޜ  ������>;����X)�׳ ��s    c�i��u:�=� �`���{� 8?w�۲e��Fķ�; ���٥��m�    ���ܹ�Z��� `�=}��'�# 8?w�ۿ��R���  j�����    ��x� &�ۚ��gG p~� -������X��  ���P    ƃoy 0YN����+;�3ph�����#�#� �@9   ��[\\�Ɉ��� ���Zkaa�� \��;�(��-� �+�9ryv    p~�N痳 ���v��5���3p�/"�:� �R�/e7     �Wk�# L��fgg�o ƀ�;�����  `��   @K---m����; ��)�ܓ� ������'O�'"��� F���wH    �̳�>{SD���  �ɝ;w~$;��1pMӜ.��;� �gΜ�>;    8W���# L�Rʯ�۷o9���1p#�^�m���  �!    �P�շ; ��u���Ȏ `��������"�� �`�R�   @�,..�dD�2� ���r�-�̎ `���L)�m� ��\y�ȑ˳#    �p1 L�Z�=� ���;������È��� ``~1;     8��; L�R�#sss��� `}��L)�F�۳; ��qX    -����-"n��  �ײ X?w�1��v�YJ9�� ��6M�5;    �x���]D���  ⩧�~�xv �g�0�8�T���� �@�ڵk���    @Dxq &F)�=MӸ@`���~���� `0j��    �|����� l��;�����8"��� �C3    Hv�ر�Eī�; �������������Z�od7  ��;���    �f�~�E 0!J)��n `������̻J)��; ���v����     Ӭ�j� ��镕��gG �q� c���O�Z?� ؼN���    �4M�5"n��  �w>�tv g�0�:��'� `�Z�{�h    ���ر��E��� `����-��3ps������~9� ش];v����    �R^X�������G�# �w�	��t~3� ؼR�C4    ��� L��g �y� �̙33� ��9D   ����_ZJ��� `�Nmݺ��� l��;�x�[��O�� ����;�,;    �I��-� �@�o���'�# �<w�	QJyGv �y333���     Ӥ��K� ���Z#���0p�����fw  �f�    #r���n���� `��znn�ϲ# w�	QJ�~�
 �ֺ��Z�;    `<��WGďdw  ����  ��`�lٲ�]��� lB)�_;v��    ���=� ��=��t~';��1p� ��r�7#��� ���z���    `��}�� `��Z?0;;��; w�	���=� �oOv     L��ifJ)7dw  �SJ���0� fnn�#�k� �ƕR�4M��5    �ݻw�>"vgw  ��>��`L L�RJ-��3� ؔ�ر���    0�z���� �����R�# ,w�	����ΈX��  6���p    ���rSv �)˵��ʎ `��&��Ç���~2� �8�k    0<M��D�� ��||nn�[� ��;��zwv  �q�֛���?    ��]����; �MyOv  �a,0�N�:��Tv �a�߾}�k�#    `����� �M��֭[?��p�L��i�-��?� ظRʞ�    �D�NgOv �)�ۿ��� ���`��z�wg7  WJq�    ؽ�޻��z}v �q���d7 0<� l~~���Jv �a7?~��    ���ɓo��� ��=z�С�dG 0<� ���;� ��]��c�]�    �ˉ 0��]J�� ��;���ޓL�� `c:���6    �Z�� `�j��e� ��`�:t�"�� `��d    ��h�fkD\�� lا����>;��2p���wg7  v���ǻ�    0	�o�~mD���  6����� ���`
����G��� `C.}�'�Ύ    �I��v�d7  �L���Pv �g�0���N�Z� � ؘ^�wsv    L�Z�� `�>������ ���`z�;;  ذ=�    0��E�u� ������d7 0� S�ԩS_��  ֯�r��޻%�    ����ʛ"�� `C�|��^��� F��`J4M�/��vv �!�N�8���    g��=� ����޽{{� ���;�tyWD�� `C�d    �83p����t\�0E������."�<� ؐ=�    0���y^D�)� ؐ�����uv �c�0eJ)��n  ֯�rý�޻%�    �Ѯ]�����ew  �Wk}Ov �e�0e�{�ߋ�3� ���<q���#    `�Z�d7  ��e˖�eG 0Z� S��[o�ND|4� ؐ=�    0�J)7g7  �?o��ofG 0Z� S��M 0��   ��=z��Z�Ogw  �WJ��� F��`
�޽���O� ���R�o�fkv    ��Z��DĶ� `�N�R>����L�}��-�R>�� �O�u����ߘ�    �ֺ'� ؐ���>����L��e  ���tn�n    �qRJ�M �P�ն`J�L������G�7�; �uۓ     ���ѣ��Z�� ��m۶�Qv 9���޽{{��dw  �SJ��i���    0z�޵�{ ���߿�Lv 9����� `��Z��޽�u�    0J)7d7  ����mZ ���;�;x����� ���Z�   ���� ��ۧO���� ��L�RJ���?� X7�r    pǏ�Fě�; ������i��� ��L�n��I' 3��k�%�    ���_��k#��� `}lY 0p�r���_��  ��w�u׿͎    �6��z	 ��?��%/y(;�\� DD��+ ��n�{cv    ���; ��R��������  ��; ��vߛ�  ���9    ����  ��%� �q���/G��dw  �b�    �q�ر�G�K�; ��+�<>;;��� ����� ��+��ΟȎ    �6���.� �1Sk��RJ��  ��; ���7� X�����    ���`���}�3� |�����"�s� ��8�   �U�� ������Ɏ ����Z�_����ޘ�     ms�ȑ�R^�� �]���� ���; ���t~/"jv �f���;.͎    ���!"Jv �v�nץ� |��; �w�����R�4� X����̛�#    �Mj��g7  ��7���_̎ �=�8K��/b`�ܐ     mRJ�1� X[ �b��Y����#��� ���;    |�ѣG/����; ������ ��������#"���  ��ڦi�fG    @�Z�����(�<2??��� ����s�R>��  ��%�v�z}v    ��`��ZmT 8��; ��v���^v �6�~���    h	w /� �}�8�-���͈��� `mJ)�    �zǏ��Z���  ��K���� ������Y 74M��;    ��c�=vUD\�� �M���� �� �*�| "jv �&�߹s竲#     ��`�t:���n ���X����^k�\v �f�    �j� 0V����|v �d���|(;  X3�w    L�� ����~��R�; h'w Ϋ���� `�n�    �,w�u�+"�'�; �5s�" �e��y���5"�&� X���}��/͎    ��n� 0>�q�ԩ�fG �^� \P���� ����}O0   0�j������`�4�� ������$ ��R��    �ķ1 ����n ������������ew  k�f    �Α#G^���  �䩝;w>�@��pQ��g7  k��cǎ�Hv    �R��ƈ(� ���Z?�o߾�� �����*���x�����Ɏ    �Q*�\��  ��G� h?w .��.{8"��� \\��a    �ƥ 0�۶m�ǳ# h?w .j�޽���� ���);     Feiii[D\�� ��}���?�@���&��g7  krm�43�    0
���WG��; �5�Hv  ����59u��'J)��; ��ڱk׮+�#    `���`<�R�G�# � �I�4�k����  �ġ    S���[ ��G<��� ƃ�; kVk�pv pq�V�z    L�� `<|$; ��a��z|4"z� �E9�   `�;v��#��� ��J).U`��X����oE�g�; ��z�ѣG��    ô��� ���ggg�*���a��z�E- �_���Ύ    �a�t:�f7  Wk�h)�fw 0>�X��e  ����^   �D��^��  ��G� /� �ˡC��_��  .��b�   ��j�f&"���  .��ɓ'?��x1p`�J)��  \ԵM���   ���}���FĎ� �>�4ͳ� �c ֭��?� ����K/����    0�n��� `MlL X7w �mff澈8�� \X��w�   �D��^��  \����ǳ ?� ������Dğdw  �   �	�r h�/,,,<���1p`�<! ��   ��s�m�� "^�� \X��c� �'w 6���},"jv pAW.--�Ύ    �Aڶm�uQ�; ��ry" b���>|�Ɉ�Bv pA����7fG    � �Z��n  .��^~����x2p`3<% ����     �� ����Ͻ{���; O� lX)�SR �r�Vw    &F�4���j! ��M	 f���=������  ί�zm��dw    � �޽�ʈ؝� \Poyy���# _� lX�4���	 �X)�_;v��    0�^ϋ� �~�ַ����# _� l�'� ���:�   `"�R|����%`S�ؔ~������ ���   0A|���+���)� l����7"�� �9�   `�;v�G"�U� �=���O�yv ����M��[ h��wdG    �f�z�k�� ��MӬdG 0���� �@�͔R�Ɏ    ��(�x� �φ�M3p`�v���PD���  .��    c��zmv pa+++�� ��3p`���۷�gw  ��   ��Uk-� �ݗώ `��0(���v�.;     6���~eD<?� � � �������av pA?~�ȑ˳#    `#J)o�n  .����0p` ����>"��� ��C@    �U���� ����t:dG 0��R�_�@��   0�������}&;��`����Z?��  �_����    `���y^D�:� ��Of 09��n�{D��; �ՕR^�4�Lv    �ǎ;���-� ����1p``8�TD|.� X]�u��;���    ��(��!� ���.��G�# �� �'� ��ޘ     �tMv  p~��������� `r�0P�VON@�9   `ܸ� ��V��2p`��m��pD<�� ��s�    ��{�ggD�2� 8����Of7 0Y����������; ��jiii[v    ��3�<����fw  ����Ç���d1p`�j�����ں����    X/@��qv  ������v�� �b�~ߡ     c���[ ��� g����8q⑈�vv p^�d    ��@��z��� �<� \�4�Z맳; ��zcv     \�w�qiD��� `u��/>|��� &��; C��t<A �u�ѣG/Ɏ    �ٲe�"�dw  �uv  �����p�; ��L��{]v    \H��Cv p~�N�6��0p`(<���fv ��R��A    Z�7, h����� �L� E)�F�� ��j�   h;߰ ���r���'�# �L� M)�ST �Rn�   �͎9�xYv ��Z��� L.w ���rv p^����;weG    �j:�� ��\z�0�04�RD|+� XU���^�    ����� �b�N�� &��; CSJ�� h�7f    �jJ)� �^������� &��; CUk�$ ��5�    ��Z��; ���� L6w ����  �   �:w�u׏Eċ�; �ՕR\v�P�0T��bD|+� Xտ>z���#    �_*��1� 8����� �l� U)��Z��  VUz���#    ��\�  ���/,,<��d3p`��  ��a!    m�w h��� �|� ���� ��J)o�n    �����A h�R��; Cg���:t���� `Un�   �5���"�ǲ; �խ��ܟ� ��3p`�J)5"��  Vu���⋲#     "bffƋ� �^_=|��� L>w F�U �^��k�     "��b� �e��H�0�V�� @K94   �-j��U@K�~ 0*� �ġC��6"���  ���   �6����x}v ��Zk�?;��`��(}:;  X�Og    �����#�� ���<??��� ���; #�* h����;";   ����v�4 �e����02�n�?; �R333   HUk}}v p^�g 0=�����GK)�gw  ��:;    ��� �Sw F������~:� 8W��u�    L��� �U���C�����0p`�j��e7  �2p    �ѣG_/��  Ve��H�0R�^�S� ��.����4;   �����\�  -�2C F����ZXXx<"��  �Qfff<   @�R��� ���+++dG 0]����� �B   H�� h��u뭷~';��b�@w h�)�Z    IDAT'��    dq� �P�����3p`�z�ާ� �U�.;    �鳴��;"^�� �����0r� ���Ç���G�; �s\�4��#    �.�>��UQ�; �s�lٲ�� ���; )J)~� �e���WdG    0]:�����>���� Lw R�Z����ݮ�D    F�7) h'� R������5� 8�U�    L��� �s��}w R������_��  ��0   �����{�D�� �9�K)gG 0��HSk�K_ h�Z�U�֒�   �t8y���-� 8�g���NeG 0��H��t��}v/..�<;   ��qUv  ���� �^� ��v�DD��  ���v_��    �Ը:;  8W��0���e�@�[n���hv p�~���,    F��� h�^���lv ����l~� -SJqk    CWk-� h�R������2p U)��� �n�   `�9���� �l�V�����le  �xɑ#G^�   ��s� ���
�f�@���]D�cv p�Z��E    ���� ���ʊ�; ��HWk��� �l�N��"    �� �ϣ�~2;��f�@:O[@���   �as�; ��C� `�@�N��`v p��    �m����Z�e� �9\R@:w ҝ8q���tv p�W5M�=;   �ɴm�6, @�z=�����tMӬD�g�; ��tw��yev    ���j� �������ˎ  w Z���+ h���    �L� �>��K)5� �h�N��+ h���    �L�w h���  ������������ �,   ����m��� �l�w Z���V���;���  �rU�4�o   `�VVV^[�; �(��>q�� �`� @��%0 �ˎK.���dG    0Yz���� ��j��i��� �0p�]��efff^��    �d)�\��  ��f��0p�5j�ED��  ��   ��*��6� 8��; �a�@k���}+"��� �@����    L�Z�� �Yz�^�3� ���h��v1p   ``�=��x~v p��>|��� �g� �J��� ��eKKK��#    ��~߅
 �2��� �_2p�U��u�����    L�R�k� ���Z�n ����V����jD�cv ��V�j   0�5@�t�]w Z���֩��iv p��    �oM �._=p���hw ���  �,   ش�i:�����  ���v Z����)���	 ��5�    ���۷��ֺ=� ��Z�f7 �3p�uv�����x&� ��-..�(;   ����t\�  ����  �a� �ξ}��K)�dw  gyuv     c�7& h��/���/fG �3p��j���n  ���   ���	 ��/����ˎ �f�@+�R<� -��t>��c�~���{����'��!�"*�\�Z�o�1������z�C�F>�-���^�K�J1�����샤1Ɯ�}H�������
�O���]   �=���c�i1>�$)�0UQ 0!   ������Lv ��0U
� Lҋ/���R�f�  n��Zkd�    `5moo?[J��� ��l6Sp`���2) �����O��dv    V�7�  ���Ǐ� �D��)Sp�	���    |^�  ������ �w ��a
 &���   ���� L�0F�,w &�ҥK?,�̳s  7y�   ��r� 2�͌0Y
� LV���K)�g�  n�	   ��}���=ZJy2; p�Ս��ײC �N���Z�/�`:���~#;    �ecc����� ���^x�jv ؉�; ���� �遭��g�C    �Zj�� bl��Sp`���C L�|>�Fv    V��; L��A &M��I�ַ��f)�w�9 ��"���    X9
� 0!��:w &-"j)�g�  ���    �I�U� ��ӧO�2; ܍�; �~� �1   ��������x4; p���  �Qp`��`R�>s�̑�    ���0�  Ӣ���)�0y�/��!; PJ)���g�C    �2�`Z�%;  �F���;q�ąRʛ�9 ��"��    X]�)��t�k�?� �Qp`U�� &b��gg    `5�Z�`:^?y���! `7
� ���  \g�   �e�Z���?�s  ��Z���X	�08d�tX�   `W/���S����9 ��"¸  +A���p�ر�K)��s  ��R�8{��#�!    ���|��� �Qp`%(���{�E��G�9 ��a�ki    �*"��� ��/��Fv X��; +#"~�� ����     L��; LǏ"�f� �e(��J,��t(�   �wH 0FX%
� ��a� `:<N   ���f  n2*��Pp`e�<y�祔�9 �R��K   p��������pv �:�� �w VFD�Rʿe�  J)�;{���    L�0�  ���K/�t>; ,K��U�b ��n�X<�   �i���  LDD��ƨ  �w VJ��G� ���p   �wG 0� �w V��; LG�uV�    ؉�; L�� +E���r��ɷK)��� �Rk�jv    &�8 LD���� `/�X)QK)�7; PJ�H	   ���?x���Dv ��Rʇ/���;�! `/�XE�,�i�j��Ε    ���W�>[J�� ��v V�" ��G� �RJ)������   ����� 0����Qp`��f3�/ ��Z��    �wF 0FX9
� ��'N����6; `�   �;Rp��X,FX9
� ������ @)�֯fg    `Zj�F `>8u�Ի�! `��XU~� +   ������x:; PJ)�z; +I��U�� ��w�    �t�С�K)��9 �R�n +J���4��}e ��o��_�   �4�f3����w V��; +���ӿ,��&; P��Ɔw    ���" �� �*w V�/�`"£%    ��] L���N��uv �<�XY�V_�4x�   �}-;  PJ)��d ��K��Uf� &��;    ��jv  ���Щ `e)����ap�iPp   �|���}����� (e�fg ��K���u�ԩwK)�e�  �S}��   @�����eg  ������� �y)����  �졇z&;    ��� ��?O�8a0�����J��*���Z=^   �� �A������J��gg  J)/   �Wk�Zv ��R�k� �^(��҆ap(�iPp   � L�. +M���v��ɷK)�s  /   Z��+�<TJy<; PJ�u?��  �B������zv �<���3&   @��������� �O>��㷳C ��P> `�E�/� Y����>���    䨵�� L�k}��! �^(���j��eg  J)�x�   h�0�#; PJ)��e �{���:Pp�	��>��   ��n &����� p��Xy�.]z��2�� ������    @w ���Pp`�)������RJy3; �΂;   @Ӟ�  �ťK�~� ; k�� �ς;   @�^~���J)e�  �O���� ; k���Zv �<�ꫯ�   ����?��D�� kA���0�w �w��ŋOf�    `\�� �`�u���Z�w ����<f   4fwB 0�X
� ���'O����~v h]���   � `677-���X�V_"@2��   h�;! ����?�Av ��X�� �<f   4���tv ��L �6�X�V���|~G   А�_~��R�Vv h�Q@ ։�; kcccC� �=���Fv    �q��5��iЙ `m(��6�x�7#�rv h܁���'�C    0��l�~ 0��܂; kC�����s�-j���� Z�X,<j   4b� ����>��g�! �~Qp`��" �E�GM   �FD�� ��z��Cv �_�X7�e  ��;   @#� �$`�(��V�aPp�d�V�]    ���>�� 0�zQp`�9r�R��n@.�]    x��+�le� ��E�w ֊�; k����R���9 �qO�}��   ��u��5C �o8x��g� ��I����gg ��mnmm=�   ��5�͞��  �_����������� �l{{�z   ���� $�	 ֎�; k�뺟dg ��u]�q   `�E�;  HVkՑ `�(��v|� ��q   `�E�3� �u
� �#w �Α#G�,�\�� ��	   ��j�Ogg  �@ ֎�; k����.���� g�   `��9s�K���� и�<�Fv ���XW�P�\u�ܹYv    �G���  ߛ/����� p�)���~�  ���;�<�   ��1��� ��? ֒�; ��! �E�_gg    `��� ��`-)����ap��|V�    ֔q �� �%w ���˗�*�|�� �   `ME�q H6���������Z��~(��4; 4N�   `M�Z���  ����SO�<; �w �V�կ�  �/   �5��+�<ZJ��� ���s�=�� �A��u�W\ �멾�;   ��իW�*; P^�  �E� ���u�w ���C=���!    ����;�� Z�� �3w �����w H6�Ϗeg    ����>�� Zg��u����:u�ԯJ)�s @�f���N   ���� �u]g������ڊ�ZJ��� вZ��    �_q,; 4������� �E����X�D;   �O�Ղ; ���� ���Xk�֟dg ��Yp   X/}�w��'�s @�����Xk� �5/   �5r�С�K)d� ���`�)���f���; ��ʹs�f�!    �?f�ٱ� к�Pp`�)��֎?�A����9 �a�~��'�C    p��c $3���Sp`��r rmnnz�   X�z  �G'N�x/; �'w �^D�r �p,;    �ͱ�  вZ��� `�)���j�� Q�ժ   ��8�  ��� �~Sp`��Z�� Zǲ3    p�3 �\: �=w ֞�; 䪵��    ����~����9 �e: �@�����o}��R��s @�����   ��9�R�Fv h�0
� �=w Z�Fv  hU���W_}�@v    �! ���S�~� ���; ��3 �]�|�+�!    �g
� �("ވ��� ���; ��� ������    ܛ�8�� g��&(��
�< �e�   `����\� 4A��V8�@"�^    �� ��} �	
� 4��ѣo�R��s @�j�ǲ3    poj�� QD(��w �����o�R��� ����'   �
���`)���9 �a����� 0w Z�Kf Hb�   `�:t�/�� d�E��W�C �>h��; �y���    +h6���  ��y �
� 4#"���  ��G�>�   ����  �8w ���@K�  �b�8��   ��'"�eg ���< �w ��u�� $��fV�    VT��� ��y �
� 4�ĉJ)�g� ���ev     >7w ȥ�@3�h� $��   ���� @�߽��Kf� ��(��w �s,;     {w�̙#��?�� ���  0&w �Rk}#; 4��   �jr� �"B���(�Д��U3 ���ٳge�    `o��{2; 4���h��; M��f�j�<1���";    {���  вa���w �r���_F��� Ъ��
   �b�ap� �j��h��; M��~����� Z�u�w   ��t  ��cǎ�� cRp�E�l�<־    V�; ���s�=�� cRp�9��7�3 @�j�־    V�; ȣ� @s�h�w ��1   `�D�; Hb��)�М�l��� �0��   X!�����Xk=�� Z�u�� �Qp�9׮]�Yv h��/   ����a�  �Z�h��; �9}���Rʇ�9 �Q_����   ���w H4��; �Qp�U� ���ѣV�   V��; ��t����C ���h�ϲ @��aPp   X�. ��,"jv ��; M����3 @��~   ��a�� @��I
� 4i� ���   �JQp�$��@��h�l6s�$�Vw   �a�  R�6 �$w �t��U� ���   �
��F)�� ЪZ��; MRp�I����R�G�9 �QV�    V�?��?>ZJ9�� Z5�͌��$w Z�Kg �a�   `D�{ �������� �h�/� �#gΜ9�   �])�@��GD� �hV�Ղ; $���    �]��/�3 @�t h��; ͊���3 @ì   L\D���$�� 4K��f9@�_    ��p  ��> ���@��� RY�   �>w8 ���:�} 4K��f���K�R~�� Zd�   `�j�
� ��h �Rp�i�V���~o   0m}�w��ǳs @�"��'~�� �(�д��K/ �a�   `¶��+�lf� ��Zߊ��� �(�дZ�_z@�    �X,�� @c} 4M���E�[� �Q���?x0;    ;�> �c���)�д���3 $�t���    ؑ�; $�7z Z��@ӆap(�$~s   0Q�Vw7 ���:] ���@�N�<��R��� �(+`    �n  ��; MSp C Ha   `�"�� ���'��gv Ȥ� ��";  �H�   `�j��gg �F���~� ��h^��|v hQ�u_��    ���� @ Pp��u��� ТZ�gg    �O}����B)�Pv h����<w p8�a   `� @��8�� �)��<�����/�Z#;    l>�+�@��0�@��h^�u�(��� Р��|�;�d�    �O�� $Qp w (�w�Y)�7�9 �E�X
   01a� �\�rE���)��u� @����R   ��qg 9>�����e� �l
� p�/� A�u�   �ǝ �8�  �@� �;�  �   `z,�@�| P���RJD���  -��*�   LL�U� r(�@Qp�RJ)���! D��R   ��qg 9j��3 �(�@)e6����  -��   0-}�,�|!; 4�8 w (��r���wJ)Cv h��]   L��֖A ȣ� E� J)����WK)�e� ��D�S   �	���	  �b�x'; L��; ��3 @�>{���    \
� ��ӧO_� S�� 7��W_ � "��    �M�� 9t �w ���; ����)   �tXp�
� p��; �Pk=�� Z4�GS   ���w5 �@g �@� ���� ���:�    QkuW 	"Bg nPp�666�gg �y4   �� �F� nPp�>��R�"; 4H�   `"j�
� �`6����  S�� 7<���ۥ�w�s @�<�   L@��])��� Рz���w�C �T(��-j��3 @�,�   L��Ç�TJ��� ��������  WIDAT�! `*���� � �    0����  �:�  �D� nQk��/ �c7~   @�Z��� �Q�
 p �ED��� t��|$;   @�"�  �� �B� �د� @����x
   �� ��U �[(��sh��0|9;    � ��U �[(��-��C# $��k   �|�0����
 pw �ũS�>)�|�� ZSk�   �� ��A� n�� �� Ƨ�   ��K� �Aۗ/_�Mv �w �M�U� F�eg    ��������� �D� n�u��; ��ϲ    ��W^y��r4; 4HG n�� ������ ZSk}4;   @��� ȡ� �Qp���Z`|P   ��s �CG n�� �� ��    Q�u�g  AD��< �F� n3��; ����3g�d�    h�?�@ ���; ���>sx�V�    ��Z�� @ ���; ܦ��˥���s @kj�V�    ���Vw ���; �ٻ� �AQ   �D�w ߕ_|�w�! `j���|! #��#*   @�Z�� ߯"�f� ��Qp�;Sp��Yp   ��n Ƨ�  w�� w�fg �yD   H�`|
� p
� pg� 0>w   �$�Vw �n ܁�; ܙC$ ��J   @��ﻈx$; 4H7 �@� � ""`|�   lnn>\J�e� ��DĻ� `���>���wK)5; �dw   ������ 	����)���}���av hIDxH   �ax  (���)����s��q=r��9��   ��; ���'N\� S�� ;����� ���|8;   @���  ���  0U
� �3w �l6{4;   @�,���t `
� �� 0���m��    #�� 0>� ؁�; ��:�I YD(�   �lw2 0���I �(��,�����   �ϝ �O' v�� ;p����    F�� )t `
� ���b�0	 �Sp   �; ��= ؙ�; ��ʕ+�Rjv h��T   �����f3w ؁�; ���k����s @Kj�~�   0�3g����� ��z�꯳3 �T)��ݽ�  c-   `D `|WO�>}!; L��; ܝ_���"B�   `D�V�1 0��"�f� ��Rp��Sp�qY   �0�c `|� p
� pw� 0�#gϞ=�   �!�`d�~v �2w ��Z��; ��o�   �Sk�bv hM���� `���.��Sp��E��3    4�] �,"t �.��.,����ax8;   @+��s ��E ��Pp����� Ff�   `<�0�������Sp������� �Q   `$a� Ffl �N� ��ԩS��R.e� ��X   �����677��.�`wV�`DU   �Sk�� �_�p��! `��`��i Q�u+;   @C� ��>��~� S�� ���*���"�j   �x�� ��t `w
� �;�K QDX   ����z��r$; ��_�`w
� �_O��j�
�    #�z��{ YD��� �N� v�u�� �1V   F����pv hM�U v�� ���� �1
�    #�A� FVk�A �](��.f���% �K�   `� F: �w ��b�p��qm�}�
   ��j��`d�`w
 ��Ç;\�����   �Sp��u]��  �Pp�]|�߼TJ�,; ���
   �φa�Bv h�|>Wp�](��r>�  -�����
   ��"� ���>�? �](��"�� 0"��    �/"�E �u���k�! `��`	�Vw ��;   �������q� ��`	
� 0.w   �QXp�q� ��`	�	 #�A�   `�)���t `	
� �� 0:w   ��� Fd\ ��� Kp��qE��U   ��g� Fd\ ��� Kp���)�   �Zk�R��s @K���r�`	]�9d��,�   ���>ZJ�e� �����(����C& �hw   �}t�ڵ��3 @k���r�`	p��Yp   �_�0(��Ȇa�= �%(���?~����� ��   �� ����; ,A� ����av h�1   ���� Fv��� X��; ,ϗ� 0���Ν�e�    XW]�meg ��|����� �
�`y
� 0�x뭷�   ��j�
� 0.� X��; ,�a F����`v   �u�^ `\: �$w X��& ���:��    ����� FTk�9 �%)���"�a F�X,<�   �� 0�� ��Pp��}�  Z�   `�Xp�qu]�s  KRp�%���� Вa<�   �Z��� ВZ�� ,I� ��u݅� ��    ��� �N� ��� K�� ��l   ���� �� X��; ,�a ��   `��Z�fg �����)����a��� Z��   ��ܽ ��j�: �$w X���}M �:�    `�)������9 �%)���^xᅫ��ϲs @C�   ������f���; ,I� �Ɓ FRk��
   �Ν;7���� -�x� ,I� ��Bv  h��;   �>x��,�Dv hȕ��d� �U�� {����Xp   �����] `\� �
� ��V�N IDxh   �����] `\� �
� �7� 0�    �`6��w��[< 썂; �ͅ�  ��    ���z4; ����`o�`o:`<
�    ���:�. 0�Z�1= �w ��N ��V   �}0�{ QD��=Pp�=p��Q��޹   �>�w �� 쁢  ��0� 0�x��Gg�    XCG� @Kj�� �
� ��`\���G�3    �� 0.] �w ؃Z�� Вk׮yl   ���
 ���`o�`��s���f3w   ����z4; �d�X� �(��<xС F�X,�   �Z�; �w �w ؃��ۿ������ Z�u��V   ��,"ܹ ������� V��; �AD�R�'�9 �[   ����  В�����j�r�X� wT�=�����>�%�1,�"q	��
�IHȆ�{2����/R5�}'�]+3��� ���= ��e   �)ܹ @��߿�  A� I�wO (b�;   �� �����p�= �� �� P���   `<w. PGc  Iw ���� �("���    ^��� ��h  I� I��� P$"^͞   ���  Dc  Iw H�;|@�;   �x�\ ��� �$p�$�; ���&   0�� ��J< �	� Ͽ����V   ��>~��� �2�5� $9�@ޏ� ����   0�ϟ?ݷ @!� O� I˲8|@�   �\.w ��1 �$�; ��| �{p   �z��o�Z H�@R�ݿ��HD��   0���� j��=  �� �� P'"<�   ���� �e�; $	� iY�; i���   0PkM� �,��<�; $E�W@���   t>�� P�= ��@Rk�� �xp   �z�Z(  �,��$�; $]�W�; ��   `,��V�]c  Iw H���u��"�w�    ��ܷ @!_��<�; $����| Ա�   `�eY� PKc  Iw Hz���O���� ����
   0�/�@���� I� �8�@���{�   ���< (����/ �$�; l?f�  �߿��
   0��� �Hg�  {#p�z�̞ ��r��   ƹ�  �����:{ ��; l#p�"��Y�   0�� ��k�  �Gw ؠ��
 E�e��
   0H��w �cy l p��eq�"���]   �w- P��< �@� �� u"�w   �q� P��< �@� ��B���|��
   0�� P��< �F� D�C( �^�6�   �Zs� E�E� [��mlp�"6�   �c�; �i�� vI� �����b    ���HD�g�  {$p�m~�  �����   `����� `�� ��� P�w   �A, �R�8 `�; l6�@��p�   0�M� P�� `�; l�{�� ���γg    xAܵ @��� �	�`�; �qv   g�=  ȫ>��= �H  �i� ���[�    �q� ��9{  ��; l��3 �Q�   �r� ��u�@�� 6轿�= Ekͣ+   �8�� �Hz�w H��!p�"6�   � 
	� O� ۼ�=  ��   `(w- P("�1{ ��; l�Z�@�֚GW   �q�� ���� Iw � "�:{ 8�eY<�   �� �Z6�@��+ l#p�:ή    �X&  ���  �F$  ���Hk�<{   �D� �� �$p�m��  �""�    �k�Z��  �F� ��� E�    C�k�Z��>}���! `O� �������tz={ 8�޻GW   �qܵ @���Ƿ�g �=�@җ/_�~�
 ez�~w   �� �XD�6{ ��  $-���3 ��D��W   ��~��Ξ Jg  	w H��Ϟ �D�   0Ʒo�ܳ �: H�@��' �{x   ����= ̡3 ��; $�� �<�   �Z[g�  �3 ��; �9x@���   pss� &�H r� ���	 �z�^   X��= ̡3 ��; �9x@-�    ����3 �A�  A� I���� �Hlp   ����= �q7{  ��; $-�b�	 ��    ��g�, 0�� ��@R�]� �\�   �� ��Z ��@��_ (��   `�eYܳ ��d 9w H��0 ��   `�; ̱,�� � ��Zs� ���   `{, ��k� ���
 y~?��K_   �1�����~8�N���������#�!�� ��˵��?��n    IEND�B`�PK
     D"BY$�3  3  /   images/7ade412b-fa94-47ea-987a-d6c9baa14438.png�PNG

   IHDR   d   �   {��n   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]�Uy�f���o�'YB�D��[��Z,� B���c�6E%�S�֧�$��XJ��Q�Z�h}
�<-�#�XD�b�f�Mv�ww��ߙ���3sw���͝9s�ݻ��/{�ܙ3��|�9�s���"��{�,W�\�r�J���[�%�2����,���"Kv���=�����F��t�X�gYǲ�����%΢��X��fy��,a�S�w!�ES�c����.I��Pﰏ��{Y�ay��Y^f�W�W@���K,og���d���_����%I��$���4�����7^����;�2K4x����7n
�1e���d|��f
z�-7��X^a��X�c����D�����3Kd؉DXַ�Ί֌���;X�IV�Hj��,��Ĝ��E:�p,�SD�Q�?G�ߨ}��BѠ�L�rEc-���s��ɸ�,+c�Ҥ����Z,
�5�_��cq�-��i\M�3l��>��Y�H��W��繐���!����(+���NQOG��QT�Ε/�\8����l�Q*&'bl���#�C��̘��g��#�� CC>A2,���d��1����"��%���Y� y�% �шF���ζ�l<�4U���<��_�9�岘�%�#`�*cj�f�}�U��S B\ځ�6�oPiq��^��J	u��{��ՃS~4��@��n�.&�0eu#k0M%��|�D9!K�(�q��5*�"3?ux@Kt�c-�%��~��2ۙ����d͈�d���E�5+���<2��)�9@>�f�X2���Y��D_���:���s4&�
�~2K������ P%��T�e��JG!�� ��5�N]�C�'���͋�'�C����E8/ЄW�)�+��!{5�Q���l�K�͖Q�[�&(Td9������;���yd8@c���k�:�J��>49+���t$��,��H��.��k�� v,H�T�ĩ����F�S�!�y��`�����&e'S�����}�(�د;!'xh5y�X�Z�E��PL'�b��?�B����W`u?VC1p�ɣ�Q�[a �e#/Q��CsB��/�۩ق�`��P����O����k�Q�΁DX���g�E1d\3�E�a�;��+�iё�zӰ!`��F+� Yy��$�p�����鲿x���Me� �`B�|����|�~�򘘩�u%E�9�C\h�k�i*:�p����h<B �eӵ��1Jƣ�4em�O��)�ȭ�lhb� �I��6ߛ��u�Đ��!d��@�������4;����!�Ў<��hV�&���E�o�v�źh�"�/��ά�Z���iJ���E�/�\伣Nh�0W�Y��U�"�@�Y��\�E�/Xl��g��!~`/�����i0��(G�f��1�ri��b�R�o��XX]O��-RO��"���DZ&�a &���ݢE�_訲�İA�4�%ur���ei�%��zb�@���U���r��t�LH�<q��]�dZb/�4[EZ@MD��]1L��J]�R�h��K���N�����7!֬FZ���*Z�@�h��Y�8��_��}b���>>�כ�t6[�Y�l�B��;z�EP��-[�;_@����}������hk>� ���I>�W��-ш�#H�Jщ�b6��du�%��Yv�-Wp�#�9/tXb��q_REK�zXC�wdŦ;hb�gjN5��l`IA3��(���!�͞�V���)t��銑�`��a�!��u�=y�H��J㿤�u!G�w��,�C7�y,#���~A	A�8�a)�Q]h�k�GE��|��tir�B�����.��{,y>�����&\u���$9�y�@l��4]�i�����]�!.s�M���G�wٰ�PGk$��(�Q"���vZ�R��zL���?���gĊu�GGZ��&&R0�J����R9/�Ē2M-�wş�|��kJ.��\O��x�J�#��D�S���l�@��I�ɫi��7�z,���C-�&̍�oT�a���)��� B"���I�&B\ځ���T|��#�TyK%�JFPs��
3�����n!{z+?í��Iu�Ι��|X���<��M���!�	�۴��w��1S:&!���G���$�Gz;��8� 6<#ܑ�;l��'@��
q��cg���1;A:�n�J��̊���}�خ ��k,�{�X�4��I�>?i�[ly������3y��Q1���4kE�u�Yʑ���$��Z\��5E �ɇ'�)�k�[-Z�(!�ЬL�Qn,�m�ܲv�A���_���y\��fnRF����:�^2X�Hv���.cy���x}��|AB*��N�����31/�ݡ���6B41�1�S���RS"m}�cڠ�XbeJ�d�:��ɚ�V&$���4� !��A��{�A�Tl�������"(��T�&��Q���8�D8�Gw��z�
Ŵ,A�$�R:��@D�m-6�J��T��ibT���I�]b��3�"�?2][^a�
�#Æ���"�����@
̗	�e��K�`��_�u��d!2>�r=*?��ۓWvS")�*]��*��C�cT��3rrh�hd8�df�.!L��,=х>
�I���>=�>I�����
B<d��e���̝��+��] d z�L©{��	���?7�" >bB�.�@E��F��,�,n4���rY��a s���h�*�T���w�B}�~�%�z^;�%���@T�}cS�i��2���oNx��1�����f�(,-I��C���$�~��t���~����D��P�㝎�=L�_�?�qoR&ģ�Y�S���S��̹�-�^����{k���g��烀�	CD�}.��d�k-q-���̖��lt�b6}y�<��#���J�.��F�¹	���` 1����4��aqf5A�>2��4�C\7�3tp"#*�6.4�-f#��1�ׅ�j���	����S�¿a��$'pWV\ �S�cV�x6]F9$�����q?��������hb��s��:��d���=����!��wy��7�+@����\��=$=�(�9N>��?�e����a9Я�Ͻ��Xu�h�WCnd9O�֍�µ2@@&_���7��$�|a��vT���
�^"�����4��$�-��h����x���&*��W�&P"����c�w�o�v������Y|��(�b�7��6Z�,���b{Y%�OY~�D��{)��E�U�A&ٟa����H׊�+*40)�"�Jk��k_gM�O<�qkȵ,g:_�@��;9��t&��G��n�ʛ�$ىN�ѨA�L��a:� 1'^�7����7�0c�3|��}��f���O��k�{�?��ڂ�l���^A�:4{·��D=1��݃[��Mz�,�x�\*F�O�^/���	�Wj� �↪q޵�)� %��^�D̿�w�޶��t�!/ź�}�t�Д*w3����0,�X�a���g�j�6g�D���ϟ�s���Y"Ok�'-σ`n�WF?W8^�q�C�5Ւ�]ۀ1Q�.r����F��!3��^��6˃��6�����k��o�lZ�A���WX"0�x���h��#٣�E�]��+�\NUa?U˥�j�Ŕ��D�wn-�K�$`��Ti��L-
����ihX(��P	�\��-\#�}i���Xb�pX�)���d��$�@:�3Q���9��v0x�b�Q�qL�����x���}�G���.Ie�,���L�	b4Y�̑!֐��"�:\N�5I����B.7�h��Q�@�yLB[����4�2�2�3n�8��d�)S�ӑ�I#i�F��-��~���/ɏK�s��Ig���7���׼	��E��i4����Q�[���e��!O�M:��pt��a�vVt��ͼeU��6�P�h���������J������"��@��r&�"�X�0��Sn2xHAO#i	�(ru%u:wu��<�>&"j�\�loG�ϟ���������W8����o���K�v�Uq���ʎj�3B�uE���������E�%�����-�5�D��JR�Yo�`��D�����bI��c���\��sڞ���7�})+�7��֚!������t������'^�S�dM2)7ιB$lxH�sN��F&��DT��xF��\�Y����Y8�(Y��T�d
�[�7S�4�tњ�s�}��i������F�g��ȣ�nWˋ3냿|j�]���V"�`-sq*:u�\*h*l�>~i��93�go�nn2��#L�Eo;9���^��$�o��(��z�^1o?|�B�B�S����dr�f��"L6�n}�B��y�
�A�>�YVd8@�W�s���W!�L����9j��j]�!+��/ [�p�]
!�
	`�'���z뭴\q�-�Ў�l&Y'��LL�B��%�V�	�ܹA	I���o��o���͉�-A�N��Du,�҂��*�!V��7J�Iʻ;�
���f&��:0�����:��[��r�ݡ��AR�`5B�@2X�w6�Aj@]�Pp�A��E�����B�@���{/e�Y��{�!ϳ\����X>��-G��"��R�� �i��RH�͏���LˉW�`sS�b�O���Hmv	|���z�<��JhZxȀ��c�I���@��X�UH��{H����>�ҡ��<��`2�mR#��i�-�of���,Pq�; %g�"Ac����Y��|_��5�-�d1�|B��"�B�X��E�;ї4)2���!%����a� Z� �8w����@���(��k�r���Mȿ���u1��R0������\@�I48/���/Q�\�}�_A���&J_`-��M����ĥ�~����� H�B�x�~��i���n����B�J.ER<��&�_1y,�~�}@�� �bї��:`������|:����6��P��S�ǂ�]_	����Ѻ��;�\2�߷o�����!�F��}ރeB<Z�U�Kɳ�[d���U�ti����r�CL�*p���x��xH���L7���V@��4�$����nr�x���B�������\^7� ���R��]O ?R�{I�邁[���ظ�$#���_	����k'--\�rb�`���5�@�FYUC<�`J�-�����I�7i�r}i�19�p�s`!����g&�k�ϊ��5`��͖�܈�uiI"(C9��b�^4L��Lb�d�Bư(�ii yU�
������X�𘁔=�``�B��TK��+I��L-�o0~��}�����빦�������@]=�炚�8 ��I�� ����F�G\� A�TGW_v>�Z� �����U^����]jl\�x=,���5����1b�D��3�zC�C�=��~�@�W�e�B�\b_�,5&�&Q��@PBT���pǼ@�	�m�b���!.��5Dp��0�G��e�B#u�}�=���B�.[P��-,�S��O�Rc�M�ףn�U^N�,˻�_G�ռ=�BB~Lj8��y\7�	I$�ϋ}�/��v881��PcktU�ˠN^
z�oB�l��t~X�R��$p4�q�h���p��nVTLn�wz%-�m5
��ur4��*�`^��DH�0Wq��)�p=�$��>B�1��U�5���P�UB�I��xP͓R����LC%�J���'��/���"��aB5OJ��?T�
V    IEND�B`�PK
     C"BYg�Ѧ�h  �h  /   images/4d53c106-8e41-4afb-b8f1-56dd58def1e6.png�PNG

   IHDR  W  '    �   sRGB ���   gAMA  ���a   	pHYs  �  ��o�d  hIDATx^��������u��B(��V�w(m�
PJ)�
Z��ۏ�P�-EkHq�K�������93swg_v�"�������k3���o�ܹ3Or]��i�m�>�,/�-�@I�4�q�<���UN��lҺX��߾ǯ�_W�������O�����깊*�kƍ��>��ݔ�=a�2�N��5f���b>��uA�'.JB��iX��8��-K�ʵ�+KA?C�n��|�#������G��(��(n�)s{�re�� <�w�gr(��I/����Mr�T�[��pZ�J�2I���}�*W	��[b;Q7�W���C�~P�i�b��ǒ,��kl[X�3����|&�G۲��{g��wPqB���%8�����#Á�ᾈ�\EZ
���R��ߟ=��跴�p����cr@Ӵ5F$r���7a�:��6���0��Q�L�f���#�wo�+mےY_�
�Π��mBQ�`m ��Z��ߗ�/�rR��4T�0����;�՟����h4�[�h�Ū9��V���0��!�l�&�P�ӓ���h�S���/�*n\Q�(���y�ȣ�$��:E��!���,i̕DX*X��`?D�-!�J��x�6F�Y�0����7�R���a�2�(�u�����_P�{��y��� ��h<�3��H	/�Q���@�b�Q�_�����\,��/��~o�%��m�C�h���}����&�G�X/-�	��_=b̊�oH�4�+�J�\f��R�^�dn3M��'�/!�/W!(�+a��\-����2�F~^�p?�ȳ�`�C9E�%�*'� �B�ıQPM� ����qP
�n��b?^��m:NZ���&�\�h꟱��U�°\f4��l���|��~�`TI)�G���DB5Ml�n.�B�hR�S"	�C���6b]P꜁2:.�_.��7�0����/Y����䄆.B�z!��Q�犦��O���\fa��K����k]ȉ�J2�h5|��h ��Z,�u�<�u����TI��}#�\
�����DmE�p[Q���MI��JкWV�
٪�� ��@?�oxQR�;��^%�2E�[�+ÌP^��3ٻ���$!2��"W(�G�p0�z$U�FD�T���Dr%��E���ʵ�F,K�$B�~-G�xq�-E]�u �&�KJ���J���5Uk3���%E��[�+Ì*���-f.&Iē�3�����/��"QJ��x�*I��2ꋒ!d%�b>k)�D���q�ܷ?�+�ؿ�+��K.h���Ɔ�n���:��r����h<�yI�^�
� ,W���Q�vwv�±,���"V�H�#?�m_��2_U��h��
�����H�BF�J�!�JeC!�&Ē����� ��D"q�D�g����U�2H��Sy�O��G�F��$��	�?,W���AI���d�ˤ��$�TK�<_(Bn�%r1�(�4��~�
�r!GJ�_�`��>|DZ��	�-��� <�A�����x>'+�U���Rن"o��<�F�y#f��Y~���re��Ɖ�l��b�0�6����@"���x�/�B��BҼ�b��"ց|!(�lQX�ئ�m�����(Q��&QFPڇH�D�X��+yW}Za�R�iY�L�,�>�v~���J��"ʙ�Dc�_+��},���m&,W��Aq�|6ws._܃nF�T$9$:�i=�x�Eӻ�')�L���@>�T��PR��a9���y�\}���uA�=���k�4K�C���/w!5�I��9gD"�?3��C}Ғ�'�.IX<I��J:�^"�ҝ^�̈́��0; x�6��;��1m:�J �'�G���DBb����u	��0 �Տ�k� �Ar%�>��%FjIm�zA����2��ئ�����/PJ"��*a{]���`�g�:$Nl�1���\HVȕ��H�Ց��Y\�o���M2�#����g��
�ր���q�˿�Q!	�4)����&R)y�hה�(QY^�7dѻdE��ԅ��^�u���G�uE;J�킉�/��"�H}�q���hIۄ�G��z���Qk��?_F����2q3��C��d��������E�#���q�\�7�=��|3�ȕav0�>#���P���mk��	b��GB���H�.�E$H�!�R��dE�U*V�R�_�ˈ��RR�/E�Gu�J4,.��.�i)�0кߎ��߀Ø��T��Q�m<�Ky�A�~�Ԇ�C�6���-��>��ȟtC���;� ˕av(��B.g>�;�"/���l�\�$A7�H&E˄\.�Eu�%��Gy��5:�<���K�0�lٗ��g�,%E�0�_D���C�u�p)�	�M���HI	��ʃ! �sǵ��$�R�^dN�B����޻BP��ȭ�T�T�?;��d��6����}���E��d��R���<��G��'!Fʧ<�A2B+M!��R���Je"���v"Q{O�����A2�D��zT��)"3D�}N���?�L��~�=�pl��̛��՘��`�2����'峙o�TT�Ek��(� �_I��mӍ	Ǔ	E��ĕh� /�1�e���o��h'2^�{�T�ߦT*E���*M�OIQ�U�m�ˁ4 `²Q��/N?G�%����>�����G���J�tŌjKɊmӲ��m�Xo��re���3��\S�I�B(E�E2 yP"�$��T��"�u��=(�ف|4���Ԩ-�&�Q
ףD�h=\N�u��'%�O�U�	�e�X/}���L�������V�c�<_��w��k��c�TW��w�{��E�Q;����q�`^��I/sa�2�O���|��la��/ J�� ��l1����O�BLzj	Ŋ��	6��`�	�(!o
uh�Ń�8t��H*h�#��� �Q�U�le5H$� ���%�����P>m�*��A��.�Ò�#Y��;=IF�)����7!��st&H*��=���C��#� �+x�ΛrE1o�)ܧj��q�D��A"٪���A���ml",W��Dr����t�t�	Em�;����Ϗ�"V��H��˯��]��De��co�nyb�>��$J�����	�	#�'Ax;\N��'��H��M�礗��lO���:�#�P�NE��a;���
�<�3�ԍY�unF�܍�re��Y4��岟@�$/Z� ��"::�ib�/����$�u@���H�6֥�Eq�ѝsJ$X�'�#�%�3 !�h�~D_�:���}T$�S���I��>I�����Z�j�C������2�&�_Bl������(.��
6�+ÌP�D��翌�"���$'Je@x�E��+f��3����A��>�������-	я \��KC��cN�}v��I��{��:�Q��~�?��Ҷ�O����0#�Zϰ-k/���?q�a�Ѐ��VJa	`$F?(�<hh���<:�?jG	�D���Lo>+n{X�o���bB-ᾱ��^�ǆ��5�(�]_�TV����E�/v��u��A��ͨ�Ǟ�as�A�"Ԟڙ��i���en�+Ì@�./�sg�(�t�]B $X!
�\)�zF<�%���_>�yT��$�������o�A*�y����>i)�G��|"�OIȕ�l�p[��-I�C�@�a���Á��F`�2�Ķ��,Ӝ&�NOَ���w�7�D��ƛ���w��0�^�G����׆ Q��0�si>��?�E�|�P|���.��W�S�H�qL"	���Hf�@D�^ɬ?)���4{ �ԟ�0�Ȕ�9�`)y�ž�4�z�����E]J��ĥ��'���� ��03��Q�'�M*����[ƿl��m�8)�I%��h|�l��:q��f�2!2"�N�:bYz�"Q�JK�'>wi�������H�v�b�(\N�
6 ˕aF�댳��#��,�0q���/�;��%���lO�^��@�BC�2c��?�9�Ҍ�h�upYX^��<?��~��G��Bn�.�yǃ��)b�mi�$ҁ��%AKO��xcƴ�z~vQV���V��2�I�8ц���c:��� ,W�aئu�cۻ�#�Au���A�����aa��D"Qن�'ʇ���v��:BV��h+�ى�#��(}7"?���w�1���߃qA��+Ì,T�hc�N���K<�iL�E	� ��
ң�4�?��j"���X^�Iw�QB�$?J���
����=A��?I$���@����PY)��U�/$J��H��C}�X��Y��/}�6��wR(�_Q#י��s����0#<qk̢9����	��蝥�ݮ$�C�zu��VC �V_Px��3�/B䕦0��C!���4a�ۊ�p��:!��q�ei�~Ñk�~D9-���7����"h[��L|(X�3�pw7�\�j��C'=���HdO�Zi6A 	��`TJI@m�C�����"<zWA�����P��n*�}o��c���}��{��]ڷ��	��P�"��_�h��7E�����?�0��v�������d��l8�*y�7�@%TJ�����E��ᾨ�ߔ���JK7�h��G��N�x���y���Nև���0#ñ�}�ĖD�4T"�%	���4��
�<e��ogP]���CDz׀�K웒']/g0�8fm����8񳄓8��䇟���Y0Ѹ�x��HT��II�%D9�Oe$X�&D�RD>-�v��hX�3B��6e���a���0�X��%4m��	����� ���E/	�ᕭ�h?��{(��,q��{�0vE���AUP��r�c�17!r��
�f$���a�2�H��jkhN�ws��@��'*���;F1����[w��P��c}�_ ��e��?�ąy^B<Q'
����[����yO^�+M�Xm�l _r��%�u�>E���������g{,�<*�y�4g����Wٟ�s�~C�~���~�Y�kga�J�\�H����y����z���{ne����U��)�`�`�7�0�v��J��БM�³�_X���c�M"I�?+��O�hN�:n�e�w`ݗ{�P~>"|�m��	H�$@��%~L��%y��-՟��c`{���7���A�zl�o�a���u�j<i#:�=� q�$�Eb)ډ(�(�;+���	A�v0b Zz�@�#}6���1P���:A��>�'Ḏ��þ!���0#<Q�l��!�8��m!�ئr!"ܞ��m7��~7��SL�����j����r�b�I�<�Gi-�����z��ayu��,W�!��Z�'�B'�H���h8T�S���]x[�F ꗶ�M�.n�*�+�X�1��&�#ܾt��]���0%�C�L����re���	qRur�/�Œ�+/��Mj#� ��'��-Oxߥ���z�{(�,\/�-�.�G)+/���A�+Ì�;Rau�S�j�5�(G�%�ۄ�"�Ē(]�È��b�z"o�~����p��q\�jS�gx̕���:���;p����zC����E`�2�ȁ^�:,B b,P$b}&\��^�M�����������D�?*��4T}�@����]I��t��\f� IrͷB Y�ҋRe<�zg��y"�<z?�V���źHա��h)�z"O��A���o�\|F�����Gi�J���h)>%�K��%nj��(�|�����D������a�2�HO�n<���FBl��|A�ϳ��wmB�����C_��,����՗��4�_�+Ì��oGA�Ý�"���X�l�P�6,�-�� !�K�u���p��>��p�i�S2	�o��Q]B,���z�	�9��!X�˕aFx������ 2�ɿ��ei��g��E�/É�/ D*(�l��KuK���6̷�J_��,W�)H��k[��do��z�耡O��)�������чX�g��1d����h���s��	�vCȊ���`s=X�3B��9+�na8��󇫳!D����u����D� "��6Eb�B���}n,?\6�`�u��1���� k=X�3r��I��=�ɿ��'օd���6�'�@Z����z��KQG��4�>D�!#Wz�6x�v(\��aas��,W�!�霑��?�e�r�r]!���[c^���XnI����hd?�I��~�o�	��1Z��9<� �+��7�kx��7�ubvo��,W�)H��Tu��X�a9
/WU�Q���P���Z�r����&}OgɘTB�*�����nB�dA�#6I>Hi~ir$�g�d����(���NA�4���Xޒ�|���$^H��#�Kw�M� �U�������m�GP�;Q�;P�;���{�-5G���H�|k����Wo-&ݛ� ��\UV�c���1tdÌ������{A�����2 $x�k8*��WfS�l_��yP�$�h�DI��G߉�^TF�����wp�u���T.��|\��Q
˕aF��,G��O���U����zX�uAXa���C�����]�k������3�H��;߉�˕MۥP������C��W8,W�A��:Z$1���R^>B'>��$!��������.$Pz��(Q�Y��*��߉&}����딆���z��yA���\f�(�JEV��&�INK!�T�r-mO�6C�C��	�.mSh($4"(�� �q��R�Nµ�����%}?4l�\�;�uZ�z��6a��`X�3���]7�tA�H#d N~�b�uZ�u�X�e8?�Gi���7���A���I����(}o}���%����{�A뚮��eW�5$,W�A�	���"�щ-Nn	�*���Wb(��0��*l����6V_@Ƕ�I@Q'��A��P����[*�����p��um\R_4�1=��<I�������zږe	TU�"W��"�^�Lo�H�4��]M7���aof,W�aD��'0n͇��p+�^ �`[V0�)O���X�� 4��I>6:ցiZ��I���;�$�)�0�1TNB���~wD�-��nRTe���X�3��u�-E���QѪ�<˰DK��%.�#0���Ԏ�i��Z���/�����S_V��(\���@x�$�OE�Bh���:��q����]XP��C"�����;���\|'����ٱjC���
�8��X��)\��*n �+Ì0��m�'bo��������'� �:IE��B>b9����vC�}l�7T�Ҳ�m��)�b_~B飜I�B�ay��.}l�{�9��778$@�\fRV^�8=�EY��?�8ܥsX8�ꖊd�<B�2����3Ty�mi�a���B�5E��Z���ȢK|����_�yr��JW"��X���	�`����u��k~Ɇa�2�$�<�D�S����Qy~��h�d��1D?b=m�}����"oC�֣?b[�����r+�ٶ�ǈ�)���K��uE�.��b_b�i�sXg���X�3�d������,�L�v�OxF[�6A�����yT/�6�ES�Gx]0T��@����-D�_��Ҷ�;\XN���R��E]Z/�\q)"Z���F*��x�@|~�/EU�n�W7�C��+ÌPR�ض�D�5��;p
��),�0B8"	JۉD�O�/K�K�R��`����ֽ���y�$�RQ
�{�ċ]P[�|"�y"?��	C��TT�`s��\f�bD���Tr.�c�����i�XE[�օ����D�>��A�Z��`���:T��=x?~�eڃ��M�hH@���~�/_��)�fN�R@�5ſa�>{�;�~=�W{��M���0#<��+���]���B���SWP�A
<�/Z�u�օlh)R)������/��IH<,r�����Oh��K���y�k��@q
y�}{7����E����`\���2/��<�KC,�������G��M���0#�D2�X�*d0��k�(T���&�q��M�q-��tI��褦w��uh��@rhz&z��ɇ.�)"�Ŭ�x��)��O
�A��t���Q�$EE�$9����DJ�C��wLtl�.�h���޷���:��_�5���۲'\��$��嵉Dt#`���~!�Q�$h���b�I��h� �G�"�x<~#��.C�re���*�bqcM���^�L�Ir$Z��?��&�')������.El4�@�a�z"Q4(֩L��*oC��	�}c��e���7�*�"Qۏ�%/a}-.T�&>�����k��KS��UU{��� �\f�������E���'1(��-J5��i,�<X���T�D��D��ԆD"�����5�KMc����)mSM���B��B�~)y����6�!ꖶ�:����w�	jn��5(�N�-֡� J�GH��g��	0#�����h�7�+Ì`�\Ë/������M�'�Y�����;�xnC�2�xuq��#$*��EY���'�'���!�cR����#��r���ۋ>�?���g�1Xo\5hC�X�G�E[���G㱧U��Q+�re�L[[�.�=�H�;o�r�w	_0�`�E�F����+F^=�/�#=��C.JɒP�L�(��z��t�����ړ��菖~Mo���MM�������[b��
D]��,o��d�G��Ǉ� ������m���a^_�r��I�F����Y/�2p�Ì8-^|��%���^z	֭[�E�I���E����t�Dp�N� ��+(�84}@,���
�	��.�u�#��}��D��vi��:"_��Y�����:��.#(�>����}ѕ@�>�����8^�>0,W��؎]��s�F�钅K�՗_���vO0$��EC?hHc���:��`]IR�B��1���,�d!+O,��v�'�B@^��h{@b�!D!��zie"�b��Cr�v��/V��\�R�?("yӭ�.�3 Q�/O���|��%�;�n���ဈy_7�?b�?~��\f�R�j�{�]�r>���+/��V��B6V��myR��K!

�CI\BS}�~$�#�S>]N�6�,,V���������E=�hh�<�+�Q�
D=q����p�J������/�'D=J�~����5��I��+ÌPZZZ�75�4�\Έn@{S���+P�酤��g�V!�B@q��1G!!:�uU��қ��I��M�>���i�,A�Ԟ�L�32"|9������~�/\��/P1>�ц�)�ť7)*K���1�J
����Y1����(Rz���+K��E�:F�_��'�s�����$�@�T�&��?(��`w�˕aF(o����t�IͲ!��q�dvw��b-È�&ʣ���(�e�2B��x�'�@Xi��H�T��D[��Q�H_��+E����X��6퓎�$(��q�H�.���'�Ŭ "��O,c��=�����!a�2��x�ɧ?N�d��\ק64���o@�{s!��N����oV �?��.,�R�v�`�ț`Oh��/_�~���Rʗ��u�`I�B�6�?�$��DCt�&�@d>T�>�n��j�gm�%E�=���?�E	��̋D������U�����0#�L:3a��9Sh�=�i��ˡ%�2w��Eh_�j#:蒍��t)<�>SJ)�QKeT��HW�^����ōJB��c�"_����"jb�2J�o:~��#"Rʧ�剈��a��M��(���9dIn��bߓdiIP�C�re�Ȫ�+�X�fM-M�Ri�/������Z��e�`��C��	*�1z5���5�2QB��������h��(il��[)��Kw��I.��@)�FIȈdFK_�$0_T"��b�)��I�H�ރ�L^�uD=t�D�t��!� �L_���U�+Q�����y�,W������Х=^�bT��Y>�J&vK��Ћ����.^�������,�Q�4	%���#���s/z�q�d�^>E}�"h)�J�P�������0��E�8nJa����:�O�,Ə)����E���ͤR�a�{��[�+Ì0��b�k���?EbF�~�դ5CM*	�+�C
�����дdq1/+OF��/k�8��D"��$C!����BB"����?_���h4��r*E�t������_%�ѥ��(b]��P��\���\8&J�.�*ޘ%�I�c�Y�s��$��.��߅�G&�H&~��n�2�0,W�a���6�yw�$/�U�b�PW��J�����]�2C���e����}C�&=�gUC�όD���R�vD�Ay��BP^X4�$ɒ�h� �!FQ����Z{��.p�z2K"�N�#�CQ�~�&�{��oqyOR�2�|�����A�|S�۫�m��9��M��uj6���T���a��i[�+Ì0�.]:�+�K�>�L���"06Y�(�����U��W���#��%GcK��y#f�����
#yǓ�����=w��^A@C �,%�).ܦ�W�J��E��<�;G����J�!���PW4����5Z�XR�#���Z�m�.�K�(y�0��p>�ß{KO�y�ND��1�-^£�U���a4O��%<~?�,�tL�$��uJ�/�/X�>;��f�2�Ǿ�b�5fm�'�7�+Ì0^{m�Q�+�0C=)�U�8�}���@T劲H�������f���*�Œ�s�eɿ�H��R�'"A����$�GB$1�!��PԉX�n�/�&���B7��}�����O�7%��~���h<T��R4J�OCtӍ.��P��A��C��)�����Ti�v�����F��n5�,W�A
���_x��BL<=鉥���A��z��`I2]�k�0qu���/�-#��|=b� ��}W��e⒙.�qŻd�B�.�1Ѻ'Az8�fඐ���Ja��D�+d+=JKc�"��_~�.��@ɑdJh���Rt��G�T�xE;!��g��ɪ�,�L|Q�5zH d��˕aF���׬\3�.O��|��Ta�h�rd����0��ߕc��~�!��U��?G�Q�O`����m�%!%Q��D�E}�"^j�T.?��E�~T�G�t#�(�#�~�M?G#d*$NK�ұbY�+%Q�?n_��y2�J}ZQ���m ˕aF��;0ۛN�����Ͷ��@�A>Q���b�`�7���&�C���0b{>���,K\�F^"�PDh/�:I���(y¢(#X?�$����x,1k�мDc���R$*o�N�^ ��@o��f ��DQ.-i�/�1��eI�4F+��%u��x"��D2~~�7��m˕aFe�/=��Q�^&�3]��x���������k � }�U�I_�n	�0��'���O%�aD��$Q�'A����dL��A]���b:F�zM�4��Zю.�EJɿ�O�~�xR�c��R^@y��I�$Q���%Rɋ4]�)6��2�!,W�!d3��7�xs/1����bQ��`vu��Öh�1s���M7IjUu���T��x2�+=b�!���h�I��C�T&=)��%?%��%n|ђ�/6�@$�rp�<*�z�F̡�%�(f4и���,Z"�uq�T��Y�����]�d�(�P��6���0#�����˗�����8�X��X*u����*P0M(�i�x��t#k���Z�E��ē�b������`f����"F�4�TD��巐$�Kv �3P.��r���KU�v��ܥ_j��c_��"_�dy�Wi;�re���ٳ>f��\�G3�D1RWU�i��/x�ۮ����v�^O�>�$Ks�h��dY�x�d�7��
�Cc���Px�nR�K�]z�,�K�D��m����N�)W$j�]�D�e)��*R�D��#B���'˦f�/&R��b��q����r^��˕aF )�_x��ch~'�)�I�)M��T�L���l�	 #
�{�T��X4��d�ѣ�%���Qɲ�ף��뚦e)ZDEz�lX�$7�G��_
�-�H�%1%�KJ4�ZZW6,V�O,�D"��S�eg%��S����^�W8`�2����wܻ�7��J��C��@M4VO4I�Ud�?h�W$M�*7hPN�]�c4�x<�:)�ߩk�J	�k�(TL�l�u�M)rDYjz�4�����'j/ʓ�Z���.E��#�F<vk<�<ՈG�������?�ȁ��0#��+V�hZ���~��1� f1�a$�hr@G�Fcf���m���iY��ף����eG`t�5�f�1t}E�$H�&Ñ�P�rm����X�J�.��>H�������#�J��(K�F/��Y�r�~�z[�re���8�ӏ?~:^CT�P�yHh
L���/Q�TUW�@Ō=������nPp+Qn7ƒ�����&��E���'�V}��*}����Do���P�B�X�~}���K�EV�s���7i��z$��&ω'��lEU��ǳ
����H�ׁa��G��o��g��̲y�'�4'��I����P���>�\5:����v֙�M�?.���3α��Es?Ǳ��H�H.�0�4���u𚟞�p�6����-�`a<Z�d9��r��ʫ�]���|�H�D���ԍ����ͅ��0ۙŋ~��OzB�҈"�mr�������Ab];��P���T�?~�M�E^��D4Lz%��&������Ҽ�%(~:�Dۣ
`���s�}��UV5<!1�S��(U�e@�GMil�f	��kA��zK��Л��x��VaZ�i��di�F�/ǴS֥ub%X�������?��q��a����e���8h���.�<	iمqG���k$$f���0ۑ����\�d�$�#�Ҡ�cAm�~u@�4��F�J����} h�� �\f;���O|��-
H��Ȗ����(%M��-A��3�ի*�����+�l'r��g�x�H�3�T���2�*�Z՜	1� W�!')0�ENM� �+�l'V�\��w�N�ezp��,�
�B�j�z�����W�7��v0X��}������*H��*��q����.���w)]�UdvX�������SO*���ݸ��u�D���$Я��<a]���4cv X���;o�a�W���5���U�q�8�Y(E��8��4KM&͘�+�lc,˪�����KQk�̃�g�n�0&�P��xL��G#�)g�zcЌ��`�2�6���}��f�6�v-��ۄ�xjtb􌨪@N����C^��3�ue6 ˕a�1�=��iͭ�	z��&K�
P�QkB� �k Qh�k����dyľR��0,W�ن�s�I���Y��A#T̀rY�ƲF�DQ�4�u��}56f�~+fG���0ې��|tޜ�SMC�A�`|*c�I����@�a��;��_�$�f�˕a��m�=p��_p�^n
�cC�։�U���G#�S�ô�Nx&6�����re�mD˺�}^~��d�����P�(��Dܦ�6I��>��ӯŨuT��og���0�����?�om팺(RՖ!�Qk}y
j�Q�(
t�-�|ʩ�hU�<C`�re�m@[k�aw�}褐� Y$Tb�
㫫�pL����=�l�p�	�M��+�leP�������͝���� 7W��X�c	�]�v��y�I�?�5J`�2�V���g����|1��HF�.�Y?*�(�l:��}>rCЄ�\f+��+/��h�zW�Ar-p
i_US���́���_�����Я�2��+�lE���7�z�Y�|���|ڛ~���q��,0sE��3�N�XЄ%�\f�!=��s�?w�xz���)�6�I�50��
��{�j���ig�~5�r&hÌX��p,�z�ҕ_����}d	t� �*B����1�� n��}�JY��3�`�2��2��UKV|���n�zŢն�@�d�+BM<	�e�����x�b�=�4cF,W�ق��Kw��x鿯|�_���̀��CTصq<�2�'cp����d�k���(���0[�L_���UMߍǓ�&N���r��r�.Q	�eU��l���cg��6>4cF!,W��B
����ڮѵȸ3f�'��4���O��{�թJ(�$�.��Sd��k����[2���c���8N�����u�v9#
�T

vZ֮��5k`�/BBV���
:턇'�?�bE�xX`��re�������U��.��Q�L	E�"�-�;�!��&&�q���"�����e�E�h���f��re�I&���ҥ����ٕQ#
�R��D�,N>�`�6T����8������U^����f��c��!�m{Rss�w��b%E�����U$W�T˶�q%pT��@F� ���c�Y,��˕a6�����L&��
�KA�ePQ��� 
�_Pdpe	�d2v��v=f<���RX���d3��֬n��e:�:�X.��[uEMB���d�Yf9&H*���#�3���tÌRX����[���y�m�5�e�$)�i����ٔ�q�qWIB��.�S�E���ϱ��UdF-,W���{z/���;��i8��Ir%��oa�6%qØ�cE�UW��HQ���LfT�re��i�3��ڿdێL"��U�N%����#�[Q�zX7ԇ�lf��re�����uY>_�L7�H�t�K�%���
������2���sr~3�a�2� �/���y
��Z��ɕ"����`�umO���Q�[^^v����j���+�l"�ƻ��/+�U�iz�e�lP��Iޝ,����gc�ȭ^&���re�M$�Μ�כ>��]Y�����S���� �^���'���<~``'���0� ������}}�����oX�rA�i�����`D4P5\T�Tݦ�*?0��re�M �Ν���̤SFUuO�4C�DK�\)��I�4<�J%����뱘�\f#�0Ƕ��}Y� dI�dJ%(ߠ��B���Z����w�,��*0;,W��==}��ә��������X^�P�*���ĪHݍ����`vJX��L�:����s��! �(�ڶ��ӈ"X��*�k�˓�K�<�u'���0ÀM��v� ��4�D�-��h�R��W]�x7�P�-���˲�̫�촰\f���g;;:��u� E��!]׽G[i=�Aee��*��U`vjX�3(���ֶK��T���~�#S�TM��-u]�h4
�N�,�F���F��evVX�3�==_I��Mw-�j���%���X<:.����V˵@V%��J�,�Ғ�f'���0%���o{{�E�k4@3�=��,1��?�e�&( Ayy��H�����0˕aB�@�--�?�d�c]���W��YeK���JS�\���H�ʊ��%Ij�*0�re��L�����㼟n�d���K�(%�\ih@�Pг�ァ�P]Q����=�� X�`[�����o�j�p �.M\�d�Li� ���obI�����<�\��H�϶d�^Ƈ��0�-?���N�aUסa �ݬ4@I�(UaMd�b�F�P�P�}EU��`�~X����A��gZ�tZ�HU	e���P@L�!J�0��
��d+k+��"ƿ�.f,Wf���Ў��+p+1`��Ve/��L�Pl<UI�V�`�ї����JY��˕���d2�����h9x�����B�TA��#�P�G!���tr}�e�P�X{��*s�.f=X��N��5�t+F?���P$��\�Ldˁ��Lw/8�	��Mz2R��=�a������twv|���c���8�(�1�`��N>��)�e�++'���g[���revZ۞���z�7 �A�$ ��i���*F�N��t,�����g�v���s�.fXX��NK_w�'��9�P5�Q�hP�bĪcY���::�5M�4�e1�bR�O�D�a�5�l�+���Y��a4w0B��Y)Z�Q���hY��(�hD�T*�c�nC���M���씸�S���}DS�pQ���-�Xs���Z��F 5@OD��+�?I�iW�&�revF�o�����ϔ��6�h�/�p%	b�2��$;y"�*˛b��Wˊ�2h�0�˕��ȯ[w��<p�[O?)=���l�*p�@$њ:P�S�V�C6�vc��'b�Mf�a�2;n6;�;�z�k���7����z�|�-�h�2�4,��&�q�5����R������h�4��XVͬ��y�+�>z��"-&������aڰ۞��{�Ǝ��O8�����%�|`8rev��Ͼxͬ9��J�Wx����3Pc:,X� ���U���1��X�˕�)ȭ\��W�z�ٮ�K���.X��	��DE�*��㏝��O�u���mA3��lX�̨�lk;��[�z�����@/�(�N�Se//�*[�����ߍ'b���C�reF5N.7~���;�=�GVW�/��k����Pcp%�l�z�E�hll�Y���ʌ^'��_���'��/k�`�'aU���t@e}-���e���w�����2̇��ʌZ�<���޾��O�uv�VSM���: 6$��c$�Z���蛑��8h�0[�+3*Y���+�y���u��e7�����µM����`�ͥ�[߼�����ǃf��`�2���5k�|��{.]�tiby_7@C-,hm��>�F��pl�:���'�|�ςf�Ea�2�
��oחn��k�/�ؔ�@t�8X��	K��@Q5�JU@&�uu5-?���W*��4e�-
˕5��Y��M7��mμ�-=���C&�e�퐳m���]� �-����UTV�4e�-˕-������/�|���˽�������k �J`D��ȵ��ο��'g̘��lX�̨`ٳ��ߢ�<���
�jY4�e�'[�`CY,�l:h�y_��W/�$)4e��˕���x�+޺뮯655iM�=�6@AWaY�:ȘH�%��U���?�?�2��+f��revh�����~�����֬ΘI���aΊ�Е�dE�P�^+W����k�"h�0[�+�Ò[��Wo��VKkU6��b<ru-,im��ZL�P��p���{�����b�,Wf������-w�v��s�,ni�^#��X�f4uuA���G\;{�a���|��/�R�徠9�luX�����׿s�_n];���-CK����wtA{6�&C��r��Ƭ��w��a˃��M`�2;�e�͹��w5���A������NP��@��â�f�L�VW��H@�4���˫j��_
�3�6����88Nd�}�g�O���
��<�{�z�`�jغ�n@W�����cڴ����Ma�2;
���}�>������`W&��.�]��ܓS�a섉��l8�ē_8�Ӿ�e�m˕�����Gn[�����u�@KW��(�˒0���0������`�]�ν⒋/V�+�a�9,Wfĳ�?�]���gf�Л��Ŷ�PU��",�h��kAEU%D�����u����~-����3�v��ʌh��}�׋���{[�a]['4�&8���&˰�����`�q�ds��~�˫��^�3�v��ʌXڞ{���n��R��z{{a�����E��~s�AY�`�Fhko�����ϧ�:��As�ٮ�\�I��7���W�]z6��n���
�u���A��OA*U�l\x�����4g��˕q�{�k޼�k
���LV�uC�&AwT�U�,4�f���j�� ��'�p\p�%ؔ`�1�\�E�+�^��u7\m�uݙ>hJ�B7F��dVvuA+F��d9D�8�sE8죇�v�%�~QQ�Π��\������[�]�c��[.�T��t@��W�fׄ�bTU�q�c@��ם>m������.�u}M�Ì$�u�U��N��������m�D�䡈iK_�C�*ʠEX��J4���!*h�������sյ�<3���\��k��ŷ������:��e�7_�&��B��zX��²���	hhh�L_j��[~��_]8f��G�nf��re��iV̽������I���"��MC&�VY��`M>9E��q��u(�{�~��_|u�ݦ�t�0#se�N�P=��ly왓z{�@*+G��SV��t��"�ї�b����:��1Hw��?���X��+��1��������g��On�s`$ˠ�X�5E:�d�(���E�f`���P�,��Uk��������9������ �M)�^u�����ƞ���-��]��1z�J& �Й.@'��q�d�&S��i|�{W�����V�Ìx8re���?���~��޹�ƫ^��=��{{!O@_$
k�&������������E����
�\�mB۫/{��w|����<ח=Q�rX����$�b�u@g��5�PWU���K�tég�p����8�\���������K����H����x5�&��t�:��E�t$HVVCcM��k�˿~�'�r��f���0�\�����6���?�����G*�"��
Ũ��X�������,��&�N��������7�|��WJ���c�
�+�U(tt������7��"�tZ6�Ĉu^�Ŋ�MƠ5��l>���A������;���;�Q�V���p�-f�ӷx�)���/�z~�~r���C^נ�q`~[;t)�5�z� �y��"Q]MM�w���G}���X��\�-J�\����]�u���k���tI:���(��f��*�ر�:��P��/��C�%vc��1̎˕�"���Xx�]��<��O�vv�!�PUV�Z�ai�:c:��QX����Ô)S�,��G���_=c��� 3j`�2��w���＾��玡���1Z-����:�:X��C�.�kS� �CMMD���֯��od��w�1̨���|(r+V�����\�5��IN.��C���P�o�X�&�q�lh/dA�G`�	P4m(��Z��o]u��q���V̨���l6M�?���w�{������f!Q� 9f`t��y�m��r 1�C�,�A�G�aL=X����ο�W}���;�U�\�����-���뺟}�}k[!�E Y^فU�ݰ�it�
d�a�B2�
r"��A&��I�ƿ���|󫕕�]2̨���| �m�3��p�-�w��׽����?�ryX����z -��n�~Ԫ�V;������u��S���ë���D">��aF',Wf��;����p�/�e+�G\W-�����ھ>���
}��:&�ZsY�TV���S��'G~��~�s_�D"+�.f��re6�kۑO=���w�s���mH�$�e�jh�����zd�Z�rMh��[֠q�dH�WC޴��G}���|��*��t�0��+�A��]߿��ۻ�z�7��r�� %�5�ih2�Ц:���:%zp[�����De%(��9�s�������s�^f��re��w��Oι�/?�-\2E�,�m��B�r���v�â�����t�j����
b�8Dc��K/���=�O�7�avX��z��bU��O�p���j��]�lR�T�6���+!�B!���������d�d�r�'cP[W���˿����nf����"�x�������{e;�A�d�į5���m�TV�SS�-^�]	fD���h&�����aϙ3f]r�W�VVV���[���`�2�e����_�5=���z{����B,���:��2��ˀ1a@u<�⋰��]ǈՄ1�L��n��W��O=��g��ɋUMm�f���+VW��y����Wg�ik7�xe%D�ʠ-��K��3��E==��/���N�P��ԍi�d0d%{ɗ��������%�?���r���{o΅o����+�g��Au](e	��S�n�������/����?(�8���N� �a@e2���_��ۓ&Mx0�avzX�;)n>߰���i�O��f������7��b�\�������{��H����qdТ1��L�}\v�:幯_�˒�?q�0!X�;!�EK�^z�߿�4����BM�8F�ɚrX��	�{�r��+{{b7���]ڻzA�PƎ���F���N9���N9�����>,ם7����G�^������h!���&*ˡ�B]�������9?|���>����̹��E����ںj�u���/}��?�sϽ�
�f���NBq��c\w���O��9������c�ڞOC�����
�u�n���䫯���8�UUU��P�]��1u�/��ʯ�T���ffX���,V6=��V���_�W�+�s&���!QS9À�|�'4�s�.[�h�Q��>�΢��HEdʪ�a\cd3�p��G<p�9�|3���gfX����ҥg,��ou����q��l�M������Lzɮ�?���k����KO=��?]��3�����H���PW� �XR�D���į9�`z? �0� �u���uMϿ��U��}K�%c���jP>#PU�6�����>�����������t�?~h/%�l� �d»i�iL�u��\������=t�0�&�re�.?}����A˫o쫡(U�����I㠩��bcü�}����I��Z���?�����Y{D�	H[������?������3�mFS�=�0��u�`��Noy�o�<��9m+������j�����"��;��G�8��߲[y��/��=k��e�=
��CeM5���CEe��.8��{���A��|@X�;:������e�n��;�+j��,D�qHUVC��Zp۞4��}/������v��q�/���<��ǋ�^����
&�2:�{`��w{���.�����_��0����ٱ߲=��u<�)=WM���H�ԁ�,���L�������N���k-Kߛ������g���~Z4�]��V�1���3>q�m��y��UU���b�C�r�q�u����~���Uuq�IrA�J�'!5 __��>���R��=Y��v���w\��>xLs[G����D`ʔ]@V%����v��WM�6�
`�-�u#�n�ы����MO={R�� d�3"P5��	�Օ+j?����IU�:Z[���~��������XW�ڪjH&b 2���v��K/�JyY�{�.���\w�LzJ�#��`�Ï��in��E$M�DM�d�i�=��Ϝ��X}�ˮ�$ޚ=�����k�Z��<����e�T�* ���*֙���_N8��琢��a�-�u �t�'V����t�4{���h���H����|Ey�ē��~���9�Og&?p�����}�~�;��t��aD���(�qc�,��y�]=u����`f�r��--��~���Z�~��\kkD5PQ�U�u ��a�Y�������Ϟ��hU�l�oY�x�	����WϚ=k��A�H��CMm�E�:��>���E7��`7�lX�#z{U�K�~��?��߷|eU��TM�~�ږ0�i�fO:��ߗO��>jS�&������]w���uk�4$�I���I���Zh��%_���3o�v�0�V��:�p]�gΜ���u�7s����f l�eI����d�Ǐm�p��׏�w�[刱����m:�?��/��5��#����XW��U��e��#����?��Ty�Кa�,����z�ڧ��t�C��)�f%͕�)������Z�{����9�x]�A3x�g/��o���u�m�{�E������Z��e�^x�N<��+�*��f�m�u;�f�SZ�����v�����x\���[�L�A嘱Ќ�쭯\����y�A�$�r���tv�}�o������G�X�,��ɓ'C�2���v�W^��	��=��a�m
�u{Q(6t���g����E�y��(G���)��m 7�u�Bn�q�<�뙧�DI��S3��e�z��/����x񢥻�(�dE%�R	�/����N8��>����/\a���u[S4k�^�˫~�3�����J��d� �յ�hͽ=`�:�}���5�Ɔ�����ٵ��t�������:d�9���1�ƂeY��EW~��o\=u�)���lgX�ې���.���������iB1���@���D҉r0�6���)'^W��w�,g���`��S�����mni�ݶ/o̘1�G��sp��{��/��U�&�0���6���z��'�����?�g�Z1�d�+�@N� /KP�(o�|�i76��=j<�$h
�������������M�͢1#��``�V�U������7M��\�r����O>vi��9�Z۔�7W��RPt�#qPkj�ψ��8��IG~�QS�R��cἹg�������9��um ]֡���j� ���>����_���dbQЄa��uK�8��uG�z��/�{���E2��Z,@kK3�5ԃ�E@.+��s�����g���h]�P�fғ�����s��g���g�P�,��uc���'b�|鋿?�c��_Єa��uK�jfŊS�<��W��{��q˒��N(t���	���j2�"�r�w9��_�ǎ�/H���b�����?���Y�@/��A�H�*�)��u�QO~��}����b�0#���4�2˗�晧�o~��'���,��QÀ$F�z"iU�����V�񣮯����$Y�=xd�ғx����������m0�﷬�Q�ģ�����şp���03�a�n&N.;���w�Y��c����;{(�<��V� ��C����B�q ����O:������t�5袟w�~��?_w�7�~�����7�nX%S)�-=��W.���˫�*��03�a�~@���i/�zQۓϜ�^���I�Aql��R]]5��ޯ�Y� ����S�<��ݦ>(1����g���t�������/�WB�&�aL#h(XI��Ͽ��7|��]#�03�a�n
�c���5�-O>{rz�1�i�c�`�Eb��2p�������秞|�-e�NyTu�Q۶�x���?sǍ�ڼ9���F��T�5��L.���_��W�WYY�vЌa���p����ҥǶ>���=��ang��0�te�7���xl��k*�������O�!5i�� K���A,[���?�����ˇ�E�0T��RP^YF9F����/}��=sƭA�av@X����fvv�����|����yw��e�a;��6���k� ���(��������}{b���"�=���w��n�����靝՚�QD5��PU�cÁ���]pe<��0;&,� '�����;�h}��S��7��ݝr�yP"x��H2�qp1B�AǺc�,��ß{�AD���.��"m�N�zm֧~���|m���z
����Äq��f5q�ą|�k��c�;�f�����ru����U�����	�^y�����������@Ѷ0J�@��#/	{��I�{G��iO�����Z�b�Q7���+^y��#�z��x$�|ǎ��;
�9��N<鄟������q���jY�Bs�o�}J��/�7wޮn>r�T׆h��T�[L��S`1(�c}�]��z�ɷ$�N��l�|�_GGǌ���k���?N��������&��Jږ�?p�W�p�.�����0���C��cX�=�;�����={fۛ��S�Ks�PD����P��H(�(���$+r�3�}'1c�˦����P�
/�����)����s��Oϟ�pz��P5(O����Fl�~�s��þ��;I�0<ff42z�j�U���};�z��η�:<�`���/�d���&D4���-U4 ���*"SvY2<ظ�>�Dkk�7��0�\n̳/<w�q.Juozתc�w�_UY	��j��'{�)��|5n�/�2�(gT���e'֭;���wNhz���:�̙�d����UQP��(@4yY��$�Q�О�{��G|�_e�LzF�FV]n۶������~��/����j@!o��jMM����eY�����̹W�`�} ������M�wɮXqp�/����έ^Sc� �.�X��ѩ&�`b(��PmM�&���3�˔����CU����Z^�V��Fq'�x��cn�������+���uU둨���:������f�5c�K�s�/Ǐ���)�0;	;�\]W��z��-Xpl�o����M�j�	N���"%�L��Q�#K���`i2�OY�p�!��=��{��7�ސ����+uႅ���[����7����T�c���@��j�x�����=�ӿ�g��o�2���C�����5��|督���;�k���fKKJ1x�oct*]�ێ�`�Os�
��eY�l���W��s�������]P�Π�Mfђ%'�����ƒy���lk�A���H�@}T��B$�\~�������>v��imAS�avBF�\1B��{v�,Z|l׻s�zo�^���&�fT��.��㧮C�Q�HL5n4ReEG|�������R�N}/��P;��?KW,?�ο�u��O?s(�nu�/��B]uTT�y7�j��7q���9��cͿ��012��8Q7��]�j�ܒ%w�����w5;:n��uJ���J�*^�LM��*`�lu�cǵ�������z�l�ė�dr^�g�=|`V�\y����sɳ/�tPsS�M�@ST(K�P�U��*=n�t�AO�z�פR�9AS�a��&W������f�-\���7�9�oѢ)���r9��{��S�X�ŦDt�[8)�%����)�VT�=�՚3��66�#'����`���z媣��/=��Ӈ��w4����������FO��D,w�!�<u��'\[]U5+h�0�϶���*n�XkvuNͭ\yP�o��3w�G���UN!2F���}�q�_���$f�Vޢ_�� �r�ƌY��m�����Zb��7��w$�X���C�8��|ɒ��/�>��}W�Z]����?K@eM5TUU��쁇��ɧ�����J�*�0ò��2�/vv�޳`ѱ��_X�z���c�\VS�"
�D���h�S��>1�����K~WS@�E!5m��U͜�r�n��kh�+Gc��r��D���S��~����O�I��eY�Q��|O��a@yYy~��g>s�������Š9�0̰l9��f���3��z�A]�\ﲥ�gW��`��T��/at�������4UWrPpx�����h����R1m꼊�L�l������w$U��w�7Ɗe�O��O�}�������Q�:����V�@*��h,��9c�N?���V�T�4e��(J�VO���\f��}{�,/u���{�t�hz���e��Ro�n�˪
6�/�B-����T�Y;}����{�N͘�VQ�H�E):�~[���pӃ��ϧ��
����uKƼH5fD
���gO?�������V1��|�:Nb�{������U��<tg[AQ�LP,#R���2%��"�ՙ�n�,�����]�����#'P�}�K2��.���K~�%#&��=x iR�a=�c�:��ʊ��AU�a��f�ձ̺�E��_�����׬�d��8^��:i0e�ԧ�|�B*R]ۑ?yq|�y53g>�VV.V��%h�ޠ�m~�H�Ph��t5��
���y��=��)�Xy�����I����d"�S����l�\%˶�[Z��\�r�!-K�LM�v���c?kͺ(�w�d�P��M���)VW۔�8q~��?m�C�DW�$� �6�X(����|R.���7���x���\vʢ�����ǣ��� �a�C�!��]]ݧ�kj�x����eٔ%7S�L.;f�4U�6�;g��п�)�P3yʜԴ=�0*+���Ț3��Â���r{-X�𢞮��I�ƿ1v츿��>?��0�U$W۶��r�=���|>_m�vY"��H�R�u]/�׻�w,�VV�^�6�([�q�zzz�;w�'��{�N��Ɣ)S��(JKP�af� e2��Q���P������X���b,�"�I�6�\�p�֬Y�'F��	��u�]�lƻA�a�m��Q�1�kG��G/я��P?=���q�{�wawww=
u��ɓo�F�|��a����O�!����������71R�9�Ìvx�2ÌD�`�0�lAX��0[�+�0�V���0�`�2�lX��0[�+�0�V���0�`�2�lX��0[�+�0���j��K�J�K    IEND�B`�PK
     C"BYw��V�e  �e  /   images/d004afae-d6a3-4a65-a5d4-4f8d37106046.png�PNG

   IHDR  W  '    �   gAMA  ���a   	pHYs  �  ��o�d  eOIDATx���\U����O=����"E�\>�EA���  
H���#�E��h*�*�� =$9�O��[k�f�̙s�@ʜ���g����>y�?�z�R=�A��c;ﴊ�َm&I��.�����&D����+��!׼��^�W/(��s*�G����r���y�*=e�U���ʖǰ�QA�.�v�4�h
��\�3�>�J������C�&��U�1j�g���\���N�k����Yt2��]��7��(�_��v$���h�B6���Y|��y���5j�F_b����%�m��F���9�潅�疎�e�V�m�s�e�P,a���̊�]7�/K��;W���a���l��m��%9r#b��p�U���T��BX�^�_�I%��߁���(	uDXk��Ί�Ip/���N�,�#�N�ԫٶM؁����	�q�l���i�L#J�����J5��%Q�#�E����_CXK�گZ`�;����w�����>[6Ms�mۗ��vR<���(7�]�������ˑ�z�V.6��p�4�*���P��ȕ�O�G�3z��,M�6+>���W�b<�{��JW���y.���/3����8]��c���!q%�9��z����+m�ڿ�0��sg�!��Va/�����wf���
���G�=�B,�/^�����{��k��Z��/#�^M����Z�b[�=�ǲ���8�w\c����$K�b;B�Js&.���:�}������R���K�k�b�\��#�|�m;�X���X�
���e�g�W������C}�|�
�a"�ڥ�JA5�!p/\|�J�;��"�b[�*`�\�E1S8�):��'c�+��l�W��Kx^�����iZ��}�r�.��y��!.�����B�Q��IauV[����	-�t�rTS�-r�|��<;�G��{�@d+���QH�5��|3o~]��R4�[lSe��6�ĕ ��e�V��M�B)_U�p�Z��W�k�^ڏ���q��J��i]�>��{���V�>I��nE�*��nP7㧍�s�g�<̺� ���ɪ��Ɛ������̢�	�Q�W�,6�P�i����B�Z�Btk	k���~�i��uHJ�f��<@�ľ\��cT�20yV��S}?��4���W��1!)��؆���ܠ�P(�c���e�J�޹SD*��P�D�˶\�ZU��ul.bV��*�L�
�����i�B11Y�jQ
Ѭz���K���"�ַf]����u�kh�V
nE�_�Y�����nν<�Ll�d�>l#H\	b�#3q�P>�{�F�}�J_k�D5� �s���uܒ�֪8���rQ�+�vD�ղ�+��-\/N`y�ݯ͞����~bA��3��6�E�x�7Na��6�ĕ f9L$ߓ��/dBi��
�4�j+V3V��-f}rk5�f�hI�y��d%H�BI���Vʔ?wj7f)��~.�y��$�l����*���Np_.�;�D�Pp���t��Rv�+��q2[�+�ĕ f1L4���_�M�ӏ��C�Z�ay؍��T�|+�[�b1�^�m�F�J���˳�
�Z�Q+��V�p=TG���T���
4]������u�wLg1�}��˶�Um�EU.b��W�C�J��u�,���4�n\Px�]�BdhY�ǲ%��`Z��rQ�F�Q(�}kYx�P �K@��=I�d��h�V�#"+�+�T�kY4Q����<6</�1�$n�zH�_L�������}b�����U,Y�Ѣ��8�o/���'��J���W��C�J�&��¼�h������Vq��H>l����BW�1�ζE��T}���z��Z�nh	��b?~���L�-PN����Ԋ�-�RV��嫹����a��0������Xq?��U�I�e�
y�+�������������Cc��9�l�����(��π ���""��b�>J.��%WYtP+���.*�~l�|��O+�8��� ��\�>���,Yד���y��<�G,W��z�3�gb����Mpq��u�EW�H-�/.��ٛZ[Jֶ��ÿ��'�c6�e@�J�f!��]?�DC�O²��"�}�^P ��r��^
���*Z�/��Q���d:q-���!���zn�
˳ҝ��nI��������bu����3����Z�?G�n��P,�(������VB�J�
��2�O{��X`L,������~d����Xg�j�p��$��`���WJrZ�RY�Ċ��\��r��E-����U�"vC��+���EVrP��ߗ�R
c������资Hih�;�Q�J>_x����`����)W��=0K���Y��T�7��5�[�j�
|�\:�z�
���(�,�6TYb=ǭ2���v�V.�s�8q�6+����,��\n�r���x�� ����d��r��n�U��`$��]s�
H\	b���[���P�����})���=��:��6	+ζ�e�s��U���+/t�
a�$�,�r��%H��J�䒏�SJ��f�M��m�V7w�#�-M?�����P�UJQ~E"���5�o���?*|=ߏ���[@�q�ߦ`���e�~-�~��hoR��[��E�J���?��^f̞��/y�6&�~ Bq����Ä��Yy����D==85|9��*7_)�JJU�����Qw�t=�US��D��*����z�?,�kWD�%E�ŝ����/���_-�]N��l)o�W��+U���e�I�h��$���U�[�_F�Ju��f�xi!W|u�
*}�WTވZ8����n0�R�2�X��U_{7/h�58�( P� U(��f�aT_�+'1�"Ss�J�r��5�~�W�>�)c��5x�h��ԥ�9���X�Găn��?YLq�w��e2O7���|�-+~��\O]&�1%��F�G�5D�y���dE�ݖ����D}�狗䳹�~�3���-��r�+��XPD X"�շ4
���\Y��J�U�OU]��Qe��ͻ�D��b���Z�BY�(R�)i�bs�,�`��1��]��(|�B�V��_L
v�ro앰-�ú�߁-���ĕ �˴ޛ���Ŭ4�iS�-���貥���� [g�~V����Z��5�Dzn
q�xa�RV�T-~�,Ay��rө�"Ǆ��}k���*VJ����� \�")i�Q�Y`��,\]��07�	a蓍޿8��gY��5C۟m�ǖ�ߑ�D����B�SL[��ך"RQDi'�}�L�7n�(9*+�D�w%�B&JOE�߶^�(N].��ks:˵fqj�v�g-ϰ �D)��r�r9� ��ҽK7���)W5���7?��ű�STM!q%���Z����J�`
�ZX�/�4��+ש�(k��4��\,y�ʏ���K
�YO	R��@�����Da!�
R�"�_齴5hS��\ ���r��U�T���1��	�R.m��V�b=�7P�d�L���.[޴�g$q%�:�}�������*�ˑ�N������iu DR0�]�ª���W9p�,�5��3�eThkeԼ�*��� Q�U-��b8/���6��h��8VX�"�V����7H��]�u�=�����+A�!�cn[�R�i��kF矒��1�g�k�+��j$n��6za�@��������W��h�ٽ�P�ZT��V;���o�"���d�f� ���������9ܥ�T�3+Dj1.e<� WvK3��$_��rU:XՏ����'3q��-1$�Q�LX����E���m�zK��͠�HS��R�����9s陨%����U��x���:/V�,Uv�ݮ��UQ�%*ʢVy�k�_�������i�������H\	��`���i#�=1��5T�Ay�㿸/1X����N�zP�N}����p�U�+2��(}�_Y誃@�����ܣ�_Kt�%���y��T��Q�n���g�- Dϯ޲y�`��z�Ϫ�ݿ���{/H^9p�~��l�{%��a�A{�~�H\	b6�X�����u̄�֢Өp_��c�4�����3�Ol��:[j�nn�-	|պ�Z�8��:�I�O��F�(��0e��#���鸭��'q%��B�M����&�0��g�K�I����\Sx���j,? �[�N$K@��-��V5���-�Ћ;U��d!\��k�ŖfD�7�[�:{��CUJ����wJ��-VY+�Vq^ޞ��e+�a�Դ~(|=�^f�I��n_W��#���2��kRJ�k��o��x��R��&�g������*p��FE�PS��DDk��t�l����>r�o�T�,��b�T���z�/f<���,xs���^-�3�+A�<�ۛ�F]�A�r��"�3�(�QN���˅���V7��Z!p������o�z��EEu�a[j������+h��WE��[�^ɷu�T�D�S�M[��;�}� �Z���鞇ĕ ��qr\�yK�CK��xE�I`}�Wbq���2��_�ؙn��t�{�u���?��X9�[���
�4:�v�81�������ͻ��`������t;��D�`����Ŗj͘:5K|.gp+���\X�rG�Ն@e}�SbG��=�_TD�B+V�f�iJ^ke떭�V>��L�>"M������`?U�udښhޫ�Њ�Ķ`*nA���6��-;�p&��@�W��ؗ����WUg	L�/�^��b�_����3厊u�~'p�ҭD ,��{S���ט晶"�U��Z]d0�\W.�@�S�T�V��:"��Z�����L��#t]Oa��$�Q/pq��v����y�a٫&T�\Qn_���xA���p.�le�Þ�b
?����d�����S)��R�j��!���)]���3	�tC����/ɲ�!X_��V[��JU�����^ÃyG0U�B�V�U���R�5��\�u�+��pF�^��"�ئ��ŽvmW��g����	\��F�oHR���"�?K���ħ��!�_]t0U �ȻW���mQ���^x-�xvQm��ն�y��`:�k��u�nb��uE�{���S���$��nv͚So��D��yn���J���q�FQ���+��ҍP=���U! ��n���\�0���E��-Q��K������,S1�c��I�^�s�/Q�Q���z���{�i�n$�Q'�/j+#�\!�e�jy�e!���Z����j��V3�V��υ����|�z^��n���\i�I-˵Zt�6�{�?�M{���m�=/�+A�	��ľ�J��>MPE�o�*l��	H�K ���f�vKu&a����"���c��@*����6z�ZV�L�=Iz�� q%�:�}aSg���&,����Z������߷����m�����T��5�����7��F�J���6��VK�?�@(��06�KS�c-��od]��	�l)ӥ0��(���)Q�5pL~�����D3��k�9�v��\EA���������e,A�J��=�F! .o��ږ�6�w�e� �[k1G-�Z���EP�J���k���֏B�:�@�Ju��&��H�J$7����)O�Wd_��T���u�]�}׀fE��A����
��`O�e��a&?��^]m%*���X,6��봑~7*�~�E���<5͊[���~�l������``ы1��ޮ[�uA�J����y�"H�6������YZ_~ْ@F��`h?�?�rߩ�g��%s�-$�Q'�/�˱kIJ)�jT�r#��#Q[��VL�G���j�qf� ���"(<p�+(�Pk��E����������cM;��+A�	���}�yg{#\�n��כh��n��m�s֪8�e�5m�Tጺ���[�Ƕ�.5K_9$�Q/H�3����Jnj���௓��l�-II�^m-��U�5�<���Q�����չ�e�,��{~YQ�!5�&���}�s���"���珊J� S�ն�6ڄ����j��7�2�vMD�MiiX5r�(��|��OwO$�Q?dٗ6]��ӡj	k)����L��?�t�\mu֪���lb}u`�O^B+c������g;�Mw�$�Q'��sVV�Aϳv�{�r�!��$D(���d��<Y�ˢ�u�����km�sc�iS�iZ��6���c��J3�K���a�'�;�ĕ �	9IU7���Z.��� Y�a�&w��y�\fy[=�"��ۆb���sH�X0c��BP�����K��[V�Z�'o^�����ӫ�ƇݰD��(��2�sx�*�7�Q~�*��D,CS��`��A[B~�~�+�ֶ��R�A��u,;�!޳�i~cm~���Xöd�{^W��LUQ��9*�K�/�r %^�ʪ����LA�jf�V�ߎtl=�L<�	+��y�V���Z���q����4.yjs�꿥�㤪��Gk��"q%�:BQ��!l0]�떧��֩MX��E��k	M�@��t��!Z���V��5 ař����F����jB\]�j���V��w��S3��+A���>��d �iF8~�P�D-�@�k
��be��\���Z9����`��S�����{J�]Q@��iX�`��<匁h���r��t�*�av�	�zn�{%q%�:�	�:EV�L���n�hpɭ
ֈ��QKL��)���IG8��Z�k�j-v�ІS�T�D���)���gt����љ�?@��E�f�x�����Vl��I\	��`_�!����fG�~��P�iL�B���=�������ԙR���Vz6w}1e6�{h�V���= �?@��ea��ZK|�t�Q�>:�=��D����x"���x��Ұ�[h���)�`���E�93Y������b��	�T�^�^d����6U���`�,��<�}`=�&gˎk��ʻ�qq�%Y��Z��EU�r�d	�l�rA�@؝�OW��=M7���,�+A��x�&�b�jLf�ܯ�
����Fk&�OS�T���^���HP*?�L����X��XY���Vx��g�V/�t��ĺWQ�G7w$�Qg���"�k��
�����U�O�d:�H�A+��4Y�
�ް�s����/m-��/҈�_#�ו�2���rDT_����2�4�5����j-���a���Vk(��o�g��*�O{��U����߃��8V<�nw����{NW��3�w0�J<>6<�*���p}t/?k�^���[�Q���9�%�t.���\�l��V�<�f;p)t��N���	��!G2���S�"���j�;6����D���x�`���Hh�Z�ᗼ�nmMIi�T#)�-֪Κ.�us��Y��������g
�C_��Ӻ<��X��E�D������y}qU�㸯��b���¿qx'rl����l$�Q��㱻��&�U9��f$rؒJ�W��[�����ۢ���
6g�V[Ե����\S�]>�/Uu��h�+����+�O���0(�t�<�����}�a q%�:D����������$x��L�0�-R����T[��V[j�Nwl��7�O���kԾ�r�o��)d�i�Z"P`��E�!�R�oG���b)�3���U-h��klf"I�+A�)�����0If*�nW.ő��1*�Q����A�ZV�����$T_�������v!���Jn9��	&:Ը��	�,מ��dq���X�K��1�o"��е�U�[�+A�)F�x,ݐ^f��J�F����S�� _=c��:0#��bx<S *��NX�}ݩ=+��j7 {4*���Mi�"��]��\׆V����	����9D��gN��Y�l|�Ӯuߥ{���c�k��8�W��Sx�Vsk��z7l�߂YDL�-3M�~A����9r�z��@k���W��癄x�u[�~���D��D���P4R	��`��Œ�Y2<��K���Ԕ0�����1���u��>�D�O�
H\	��I�����e�d*��S0�`ȡ����]��{
Ȟ�Wr��O�V���y��v�����刨x��T
���:e��`F6��B!�j��*<x'~Y�S��Ue��ﺁ�Ye�d��g��˺a�Bʃ^���9�ld�Z=�7,d+~���w��^" �L&�b���ҥ$�Q�(��)�46d&�{���~n@8��G�7�O&Aߚ�Z_�J.��H��FЅ�[����[���r�j寊mS�Hɭi	<���:�c��G�P�E�XJ9��5/��Q�vT�5U{RU�;����D�ݧ#�����u��ޣ6����-������a};�;��a�ʢ�	(Y�"g4ղ�X]��7=���|��{�QP�$_�ڥ|.w��f@T�;��%�88�	�_�����T��V=�Kľƞq[	�+A�1�|������~�Fc��Y�:l���"�BaZ�5��u�H�Cj�$:�UUJb=_U�A >WW5m� z�����S)�r�8�
l�6a��%+a��R*	���V���WN<�����[m�rH\	�����?���7��hn����$KU��������S�?��[��5B����o
�_��>L92��No2]:T4à�#u�s������E@��Z��o�ʒT�XѨ�$ڒ���,~Nk�؆V+w�U/��0�`4��m��e@�Jű+V�r�
��~���/f��\�0�U�^��r�R���Aʆ�VI�%n�TY�U-�Q��$�{�u�;5�E:]D�<,�+�Wq�j�u���\0P�xU�"%��~��$��|�T�:�w|/W��S�i��{��^ҕ/���>��T�]at>L�w�09dM	���o����f�u��V��<�V1���O
ߧ*,���QĝU��췚-7H�n��yK6����1\/���R��E~���2�¢b������ұ�?��p	w@̈=�� ��/W��S��b�=�ܳ�f�Y<���8`�}ѐN�.�����@�?������b���������\.��l�(�v��T'�G��Tq/�Q˲�;8V�zaY��!��*,Z�\Z���J��|6���+ޣ3@*��'�I[�C`:H\	�N��X�����}�1]�Po?���CX2>���a�f��tH��xD��eTgCa���Y*�De��1^����)u|Q�<��L�h@�<����%����Z�\��0�/(]��sQ9��W)̀t���
`M3J���F ���~$�r�,>��y',��g ��R���U�-^!$�Q�<�ēG��ŷ6Tՠ��{YccP�q4�0a[�ŉ���e&�������+�Z\�DSm�aV��g����C��@�T_lu@�-��m��lْ.�]�S��+@�D���ʖyE&{O$7F�����D�5u��\ l��>���{v�`�c�DKK�}�!�e&�0ˌ늢�|���^q�-��\�W,��V</V�pA,=�FKAa�q�� \e~���s�n����VIg�ߞ�G����ӷJ� �a��o]ן��◱G��6�ĕ �l&�h��g��V�&5��45��	F߲����w��������+�V\�g�]��x�
�\d,�w����y,�7�~�V�,ܪ�
�-7G���T�DbY�C�⌦��a�k.�~ +�ZP�6�`�Z�|;�*;�H|Q����F��D�~��}7l����V&�l��՘B�P���f.���݋��6t��&'�g�z�+�]
�� ��^
+��0�3���0��g���:�a;N�����4���=8'J��ꔫ--�>W��ݮ���a�ֲ%]��n!�"���rf���בUe4Ր>O��?`B�Ju�����F>��u2;�G��C�f�����Y��W㱿��n駯inmm5�^o�ng�At���H)Z��l\5`ZA�J��֚��f�?*-�����u��3��*�L��/�V0-�F}�\X�ӻx�E[:�\~��d��~IӴ���!q%�:�4��G���~�I�`f
�Q3��Z�L06�D��fAV�L�u=ړl:n�o�rf�Ώ6�.�XY���r�~��
�+��8�.ZA��)e
��eDq��U�%�~�
xM]�ϲ.�b�/�Z���"��n��������������G&�L%��	돰 q%�:crr��٧�-v,qEc�㠳�-�2�&Ǡ:E4&pty��O�v<̈́�WO&�ڭ�'�'/�t[<��;�O�L�ԃ@
:e����`uMg�.�X{9��y\9(�����Q�AuV�2W����J(*T�U+��)o��GH,7@E6A���Ml�_���D�����J��F��D��jժ���|�9Xi-���&41��G2Ƭ<��LQ�����O�
-	�������|� ����S����e)�� ]>?<�d�3�ab����r�.��^<��j#��Z��%�D��~OĊ���,iUb�����E��K��K� Sc�=m�}Q���[������.�^)(�M&��v%�`���+A��<��q�����e���O���Z��6����?�U�gU�e"�|Jӵ���S�5��S��b�\=|V�H�LÅOgtyz��S��Elۮ�W�:����X��E ��㢤��+���PJ97�\iVI�$�,�[4�Q��D2�&����uK q%�:�X,�?x�CG�R���;B%�I�֐Bar��Kl����v{�yɒj����1�b&�O��s,�Z"�;��3��J~^��'�sKX����m1��o�"��ͼ��.��^[�*NP�@�W�aˢ� ��U��Fg1(u���թT�\EU� �+A�#CCK6�۰Pa_M�Y��TlkL�5�34F�8��������4��$0A��XJZ&��ّ�z�s#C��o3XU�F�{l]�O�F���dM�ŵ|�GF��J��VقrYqmE*�2,����^D%U� Y��D�#vg"�����8v$�QG<��s��&2)b����V�x[�Bq���2���=���-X�eU�7��?��[̂�Y�h*��}�ޫ�Ɗ�x�ޕ��
>k�V�8����׊,WY�eʩV�m���̟�W�����f4AMne�Y����X2��.���`;�bB�Ju��{�=�X��G�2�i]{2	�P@�hB��U�������\�(�bo����4C_1�?�2�=+"��B`�5�����rcl/���!;�;l��֫��^�:[�����\�ʜݪ9�h(P5��D2q��������9$�Q'�������p�!�ˬ��D�	��(�PpIAρ�Pb�����$���=EK��.��U,�k�����Z.3-�=�ʢ _lÔ*��K"m�:'Ve�A�E[Ρ�=̥m�e��֩���C��Q!�y]7~m��oJ��,v$�Q'.\�z�"=f��<
hjnF�n��݄F6/ZLCF��偬�m�1Z�Ŵ����*?](Ov,�ӫ�ܯZ(E%T�k���>�����:��jt��`�_Y��4qJ��oWUOU�q���j�[��N�ĕ ��{�?,=b��ڈ�!���V��P�j�=ns�p��ܹ.�I�������O���	�`�ղ����?����(�K	=�*���֬딬_��Xj�y����p�,ј[�%�+�Ze�2���4��x2�&���uC�H\	�`V`���#/9�3E�D����!or:2��,=��X��6��/�E��z\?�Y��v-��h�߶����J��Vǭ��Om�g �*�-]ě���"�k��Vji��,�߯���Y���`u�+A������{�A������1�6"&ɰ���{�ڇ$M�.�o&Zk]�A\W�:�!�i~�,��l{�Im&��y�;���fOF�`U0�W��
2"���kص���������dEy/sv���+A��֮=�wæN^B�Z&$+��T3̒�E����3��'��#�I�Y����{���ȵ�㋅�I�}/&wm�rMDS��ݳ����Z���4�%�VQ6i��0�������;<`k q%�����_o��D�}u�w�ʢQS����d:�`:m5���_���|fG��u��]�дk��531��΁�i��X0����kړg�&-�.8�A��h�k���h�*)/�������3A}4���de{@�J;�l6�s�=�*;�_k/�Z�qt����b��,�u�}����d�|�!0Rd��L�~f�c���.p�PӴq]{��y�$ܲ5�5��!������H2l�)�rA��1I�_R$o=;�r6��]c#{�a'G�_	$�����ݴd��5�|"BMZ����P��QzSSf�뎸���qI�Ǚ@>�ԟ�5{̺����	�Z�:�R�[�E�bj�w3\�S���N枿�}�gC�U�]@LU�l�P�Yh.O�gƟGہ<kmۖY����b�����N`8� q%��H�P��/��ٕ5=�䠑OF�HB��^F:�Qf�x�Q�I�6bV@�J;�ލ��_�r�b�S>o�l��H6��[�V���ab+���퇾��\Č���N���xw1W4��ג'A�t%�p�Q���0	�������Y�+A�$�ܢ��qױ~#h�񛠴��heV�����x��<����E΀�5���Nbݺu�?�Բ=t݀[(B�,,jkA+T-�A2�@��nb���[9�\�W��9ȷ�򖏛�xV�q���	i�yAb}�^}�[%%�k@�*H\	b'06:���w��:IWa{.С�h���"҆��֚^�hS��G�b�A�J;�e�-;j�K��S�ӆj�X�؈FۆbZ��������TM�^1� q%��m�Ϳ����q��`� ��xUV�D#{�d�`�r{����@�JH\	b344��#�=r���H�Prڒq���<$UA^���#�ϛ�0�Y	�+A�`���w��xM����joBJ���5�F��i��~�\��J��C�J;�B>���[n9Y���J_�&YFOc�F<�Of�w��N̛�Y�+A�@^x���?���=M����sX�І��4b�<Y��a���G�	I*�������u��[o��c|�S.T�A�Y��5�"-)H�c/���w�-1��o f5$����������Pّ y�?�`g�	=�4��װp��>'�x9�Z�\�]W��x����?h``$ΧC�<q�jj@{<���`8[��'��OZke�H\	b080xԍ7��v��W����dca[��3�@�w��Eo{�� �$����<ϸ�oO��p��Ȉ��|=��J� gr�8��ć��1�ƚ#���vfr|�տ���(�yf�&��.�V=�ߵ�Ryg=��tǫ���9�+Alg|���_\��˓H������N���gdN,��>�ѯBQ�@�H\	b;2��|͵מ�)�����2��� z�F&ob���t[|���@�)H\	b�!�}�=�|f��&C�8Xܱ�[Z1�7��=�,=��K �Ys
W����Ӷa݆w�x�/N�,��6 Yy��:����@��k>���+�O��s���6ƶ����享�?}�k�˅�Y~;��dz�190����t�A��Ĝ�ĕ �!��%2c�w>���>���u�"֞�I�ګg!��Y������[2� �$$���Nf��[�{a2��X��M�!���3Ղ��V&x�ێ,1��� �,$���(����^�k�x b���˞_�ї֡IR��򊌮��';�1g!q%�m��]�×g2�}��aq����d߽пqF7l���ݏ�����&�б�����[`�B�J�}xx�����cbLT��jB����:Ҋ���.;[`44,�l���u�B�J��l6{Joo�l˅#{�-��LD��,p�>�H66�H���� Sq�5�{�Xl-�9�+A��Y���w�i�-��l�o{�+�	��^�$����eA�$8L��䣒$�������G��L6��_���,�`���e�	�-�NX[g���:&���q�9�+A�Lr��[7���!�v�ˬTG�Ud֩�AgV��,XY�b��v�z��c�S����S �4$��2�\�ehx��q�m�a�@�4�r�H��p=f�z�5�C2�~��1�u��1�!q%������''�'_�?s���J���n(����ʳEͷ�6}IQ�g@�yH\	b+�,�����rW.	��Ŕ�+շTC�g.����� v	H\	b��FFF�*�%�i����꾸r��>�
$׷Z	}]�!�M�&b��ĕ ��B�x����	��j۶�NӸ��Z���-Y̒d�h1��kjj�����Zp�ĕ �f�&GG��*��<; ��<�*�N�+�
Xn��V�hjl�;��]b��ĕ ��L&{��D�M\Xy�U,��[�
�R��'���2�nL��
v=H\	b`����?����l��V��wx2V�T�l4]�Y�O[{�Ou]���]W��������������SN����Ŕ/۶�nhH=�LƯ���f`�9���S�l YR!)�� ��V+>k����ʲ��.	�+Al����33��~�ju7P��-V%dq���_'����p#�A첐��X�}�@��]��U`��m]��WAO�y��������R�Ӻ�C�J���3500|q6���<	�_k`�jp�v�\\u]�S�\��~�����eYZb��ĕ �!��~`dx���3��s!�V���. .��sLO����:E� ��C�J5`"�140x��8�*+����,ڡUG,��se�nW�e#K���5^,����!q%�L��:3>��ǧ�<hL`^}��{�k#)��ڮŋ���ZZ��ei%$�1˲^344�I�s�� ���pC�@P���&�
b%�ō� BH\	"�x�З���|������|�VE񅕋�����+��� BH\	"B>�?uld���L�2ܰg��U�^PV�K
�$�g#���hkn�ӈ�ԧ���ĕ B�Y4�7��h����島r?+/`b�3�|�LXm����t:���9ͧmɂ "��D�P��œ㹥A�������'l��*��LX�a�b�x����"EU�	���ĕ �����G�'N����\N���������H0$��.�p��W--7i1� ����<l�=ׅ��JAY��D��$ǅ���Pً��ˬV۴`4�W%�R�a�lQWb�'�;cb|�x�e�}��X�~�|ZlCS�PUL��Ab���,l���=K��U�Y�4���4���� V²�t-����j��xS�d)-�v��oc���wƚRׁ f�ĕإ>mbt�`>�������X�r5�Ⱥ�R�,n� ޺U�%��ֵ�6�\д-�f q%vY\�Y4<0�a.���@S�v�Z�Yf�ż�B��;_u�t�4/�>KR�e ��@�J�L�M��.XKU�� ��5����a�rИE���H6&���]���bAl$�Į�f
G�
+156��[���	n����������:~ʄ�z[�+�K�nG&;����pl�7���Wy6@�Y��c#�J!7��bO�-�A�(��bH\�]�����c<��A�����`*l����3�Ј֎N4�w5�M��]"+�:�V@�J�r6m:��[o=�g��F�q��b��ݡĀx��b>�D5������k���J�	�����^.w��_ɲGm]���x�'������?�}^�w0�@*��cm�����DC�*�ˀĕ�u����~v�w�~�����=�ް��z䮻p �_��|˛�����u#���2!q%v�����G���LUAQ5�g�#o�P:�_�<�{�Y\��/>�5�듲"� ^$��.A~ݺw?��N����4��nd�G��H5'����k���?C�JlH\�9�58x�?~r�%׭m����狫�ЈXc9� IS��.���d*�4b@�J�i�|~���������}s��b*�e7`u�_ �I
���Ϟsگ{z�)+��f��s׍����������X�i��Ob��0Z�:`��g�8��ß{߻O�?�� q%�,�r��>y����6�k\+F����Φ$����^s�}�K��b�
�6�ĕ��l�ǣ����_}xt2#{�p���ף73���6�����rٗ������!q%��6���7��fժ�P&��}���6�ot�t	�@>��q���[����� �$�Ĝ��끫��W�֛ɢa�"����A(��ֆfd3�������K�Ue� q%��e5>r��?|�������66!�Lb��U�;:;: K�sE|��_�RsK�C ���+1W���r�U/����k�oR�Hv��_/�G��`��3˵o` ��G�<���؎��s��w�������'��P�m���q2ˬT��!�b.��?��N?�LI�� ���+1�~��s���ӆz{���q$.ANW�z�Zd-MMM�<�mmC_�����(����܋/|�����/f^\�Ȼp�-F.�ĳkWa4�A���d֬��_z�7:��� A� H\�YK~Ӧ��ꪋ����\&��j[^|iƙŪ%t(�
Y�p�;�����Z���a���{bb�'~r�w6=�l���L14tw����QX
��Ս��au��O~��?W��I��ĕ�u��B׿����ǁ�#���"6��G1����d$����lt/����/:�0�5 ��+1��l���k�:|h�&�:��yVu���Zd\�-��	�d&p�7�yAG[� ��+1{p���_��uw�����qL
�Zڑ�cXɆ��a�q,H����$�=�s?�w��@;Wb� ���׭���7'&106��v[#���o<9�c���021���}'����A;	W���<e��|틷�����8���J�QhLㅁ>Z2lEAsC�3��{�=��s�g>�*�(b'A�J�=k�|ە+~��[�&
6�Jk'6Y&VBO����q�`�����~��T*��!q%ꚾ���֊�~��!��`\��vt`D��rh�d�6�̒�f�������mm��� v2$�D�2x�_~��δ��NLL`�U��ъ�����zQ����a����_�����k�_� � W�.z��,���s��a=��c̱൷bHW�n|������jB&7����7�GQ'��uǦ���kz�2<bLd3x)��4�c���OL�o"���v�1aeV�[�y����G� M0H�$�D]���×<~ŏ.��yy2;��y5��ȧSX7:��L�t3bZ����^��G�<��O(�2��#H\��a�m�}w��o��7>!��"6�3a�1ٜ��ka�4��:t���+,]��3�_t�'u]� ��3H\�����/���o?����e0�E�?9�A	(6�1/A����g!8hmi\�%_8#�LP�Q���;�q�+����޻�:��X��̈́�,`#T�g>6�sX=<��	��g�k45���rz[G�\u�+���,�y�u?�a�>>�Ԏ�8�A6�@!�b�k��`����U�3��/}�K��[0�/ �:�ĕ�)��b۲������������؄���LZ.�T�#�0]�{������/_���KoA�9$���|��?����0��aڈ�|L�X���od��r]�}���X�~���/}��|%b@�J�P̗����߻j|��U�A�u0��c�^'�)d4#�"F�&�b�lܰ��o}�Q_A�H\�Ff��<{ŕ_���BF�k&&�K�1�cS���|v[�x����8缳��淼���
Wb�0���_Xu��7�5��F��xat��4�2a�b$o����&ള>������� f$����u�շ��ʕ��������mې���cº*�A��ò��Ą+�����شi���g~����l�,�ĕ�n8�\��?��#}�X�h�ST��$֛E<?���*�����0�X�^��mm����g��������J,�,�ĕ�.�G��W�t�����X�#���&�X��İf�L'0��"g�X�p7�Z��׻�w���q�1�H�d� f)$��6grŪ�]y��ǟzf��� �
��a����!�6�����~b\=�w/@s�	�����������A�Wb��w�C<s�O/��c��X:�ۯ��L��X�8�3�0]��/DKC�b��ŋ.���_w�7As Wb���vꅟ����;�~Jad��"�܂L�Ƌ}X���HBG&�ॱx��W���	˳G?w�9����@��3���{|b�����ʡ��y#��:�����LX��cMvㆆ1CE������	��#�n��yga����bA�J�"�k׾eŏ~|���,F>�dLG��	��<�\��L�t
����\�t�/�i9hjm]}��/8k�Ԅ��s��/��{�h��n>������rH57@N���s��s]�Rq��H�5�B�.�&z�_~�y����ybB�Jl5N>׹�����S
�bh잏��b����݄1UA!��`�����hnA���2�v�ݟ����Nkii�b�B�Jl�����芟d�Zv���A���7��^�K��ȧҘ�M�XE�	��cϽ�F��0��s��/��O�R�gAsWb�]��=O��o:��.�y2�Z�1!]71����xat��b��((*F�9�ZZ�Ǟ{bdho<���?�����ւ �8$��f�'����.]q�M�H#c��-@M7�����Y<��Zd�1����\���g�%H7��P,����������EA���3b�������\7�ēG���E��J,��}��L��jl#��q��44�����F�2����ǿ~�Q�����A�"���2���S����_Ͽ�rն�8�{�#k{d˙t��sxqd����L�hjnE<��n$����g��w�}nA�b��S��fk��w^���_�V�$�E�Y��=X�nr�?���a���Pd]��=H54!�J���c��g���A삐��V�z���tY�e�F��H2�;ڡ��xf�F(��0������/���$F*���`ll{���g�y�鍍��A좐�>�m7n��W���/���Y�!�H���Y�ډb{������ߏ��p����y�n0aǉo��N~�)�Q5u�C�J�;�_�=��ǎ�@N��������Y�%,9�0�8>���v;֎���u$c1�6o	��Pe%w�θ���^�vJ��C⺋3����'?��\�na�o�:ۡ4��45�I�lt��U��;x��_0U��Vd]��:Z�����_X�x��A���.�W(t����?���;ORsLa�n�1a�<�Œ���s��~�ǖk��Udh1���W-E�s������3N?+�NQ�AD q�ɿ���U7����G�q�T,B�4�/\ ��	k�F0l(8褓�Y71�����w���Pt-�:��Ӄ���]'�p�	o?�b* �����Bx�ܒ���%�p�{01W&�R-M0���02��}��<�����o��57޼{ޓ�w��T�m�uE+���?{���p��	��.���7=���7�[�T���y�{��75`����k��Ϝ~-�:�����ʝ?ܕWcp%�]�����)�������9���m�� �i!q�㸖���׻.~�7����nS����llB��y���l�%�z�����Z�����s��޿_|!kn�,�hnmÂ�n�x���������X,����9Lvժw���/??��G$���Y{:!57c��b��G��{�k�w�������?|�h�S�v��z��n�q$b��G>��=��#.A[���-:{�������c��V�p!�:-DNU0h��x���8��/�W��;W]��?�� �!��$!�L�A+MӰ�������]]��� �-��u��_���5���������,�AK��=бxz�9�]�Ͻ����a���֯X�~�����Ƙ�Nd'��^{��Y���o<�'��_0�Al$�sgbb��;��|�m}����!iP���f�ۚ�*���|��i�SO���:�}��~�?���ϯZ��hHBf��6���斦��G.��}�A/�َ穓O<y�s�\w��vm���!O�����v��屶�y�ٗ��ܑ���o~������g��yЪ!�%���q�x��g�u���M�t� ^$��kd��տ���7���w�y�.AgVh��r��3�����s��/�t���Ͻ������G�x�-��☾o5�002:����z�I'~AU�� q����>��cg���s�5�;,��@nJ�57P�jy��:�ↅ�4������|�7�����;UM��z�{ϥ�U	Ɇ�����K�.�� ��F���2
�6�a�o~v�]w�5Vtf�zF-�0fHȵ��m?���|ӛ�GR��၁�}�k_�߿���#�$�Ⱥ�i�n����U�|��3>����4��f����lf��?������l�`R58��Լh�z��.�����򥉮�=�M=�����������}}����笶64#O@U��w���oy�~QU�1�M!q�V�|��_�x�����p�(К���ҟ�*��Է�[�|�⣏�.9[�d��zӍ���/o~�X.ע0�Mqt��"ńu��y+>��_���{�� �$�u����K�����������j��S�v�Bnh�:�������?p�E�֖�<ϋ�}q�;�{��.y��GVb:]A۷���9�ux�>�i���@�v�ĵ�ݫ�x���?��#�kֵ&ƠjL$�u���*:�==��������{��c��~�ߞw�7�k����t|��Y�m̠E��>w�et�� b���ۻ���{࿳ϙ=�d�CB��	�}�5���
ZYĽ����>���io������WE���
Z���@ +$a�3��d��̙sNߙ�}���@���y��3ɜ���������pH4�����Y��[ߕ��5_ @��h�g5�����H;7�/���x��	�c��;�1��'��Ŗ={GGT*���h6C����aË6}{��V6�F�2�p ��g6T}���n�|AJ�(��0:�qX�K�P2lK�m�=ap��~r����>��g;�}.#�B��I���Iڒ���f��� �k��e��z�i�`v��m���w��;�%%��l9C�3O��%o��ͨ�2E�}��O��Ͼ��?���Z�u������S�ɮ�G}��A�k !t�a�^)�Hrϡ��O�Z�4p�>�#��*K�3=4Q�RPJ�aښ�n��	c4���4Mسc���~������h
��]�FH�$����3߿s��{��
BW�������s���������Qd�DW2SR��B��c�\��>%��C{==��>��}�J��!�������i�F�׋�O?���9�ٸ�
�+��2
o�l}s�}���dT�\l@��F#���qڎ-��9WQ�
���'�6��|��?~���;_/��+��N ��ӦN^�dɢI�zBW��e9�=�̺�v�Y{qt02� ����K���kgֿ��R�ue+Y���c~��/����Se�Or�%� ��p GQ`���<��។��B�k�����1����MgE�tc��tz3��� �����/y��ՙS'�Np:�_x��cGoz��������\S x����Tp�P�$	�F��[xϒ�0��M�P0\�j����=;����������L�H��n0''��q�X� qz�QZUqS�Ӣ+q˅��2�X��V�aŭ��b3,&+��RAST�ȡ��_�l��q?�Ѐ���U�46��Vyz��{;7o����|��^/�F2eA��A�	`=jS���gi雀��O���z�Ϟ��{��	440�JN�O�
�"0e����=Kv�Bh �p�T�l���rzc��ε�f�a��� xI�� ��t��z�c0��nw��S^H����i����}Yo��������oyz|ɂ��o���J!K�v8����~6r��e��0\�$U
��ԇY��QM!#���j���p<��\ ���
�윆��7,w�(x����9t���>��ÇjjG���� �Xk@�9~ou��q;�,Y���n; ������|y����[��־�SԾ>0�J|�T��ALv�J��H��o|�:4g5�O&��{�C~��s����ߟ
G,�Q`3%@rj
p$`)��]x�_�~��'�O�>@l�CS�HG�Ϟ���Z_=���D*'GA�e�*�u:�-6�,F���a[J��~Œ��!��?4�VŸk�����������r͖���Հ��a��������B誃��9�H�!?>���j����4�G0p5���� ��	
���c�/+�X2o���̵@S�v��[�=��s��kˎqJDV�3Xmv�&���G�~�g%�ůB誅��i��ɞ��s�o߰�ޚ�|s4
��T|*�*�@� ��{P�I���[0m�r㐬����vZ�ϗ��ko<����y<n�q :�V8�v��
�����h�G,"@]�0\?�Y�5��ޱo��#��f5���ư �4pFh�B�)$��R��M��1mt�ۺ$�f���~JT1�ٽ�[���W�7�/�y(�&�	�g@l�}Pz��w>UX��: ����p��!�t���Cg�ݹkR��1Ӡ1��j�Iu|�)/�
Syy
���Θ��� om0|�ʨSm�S^~��Gv��9���7"P4Y�3�T�I������3���E��z]{�����<���ܲu���\-:�T��(�F���03D=D�074�X�s^1�d�G���s��ūV���w��ά�_J�IM˓s�;SHN�ʕ(.*ܵx���Vk ��v��pUU!��-�9r���7�;�Q�@��*�T(�4R]�� cJ����5����,����ĝ�q��������7U߶b��[��c���f�R�R@�#���r�;n�M�������( ������*�v����}�����Mٌ�oPA0*2�8���,�����F�"�.{HK��1�S��>?��T�$)�z���o���|�%�^�,�Ǉ�v���:������V�y��ǝW���Z��&�Ϟ鮭�ٱ��8O]]6�.��a(R���(�:��(W�ysI��Qǿk���u'/��)�b:r�ȌW�������'�,	i�����tƗ�F�Qm����,��}�Պ� �F\����	����޶���ã�S���PhE�D��T�2# GU���b�ytC���&�_c:���Z^��TUUlnh������ߵ}g����t"��
��鐔��p�l������H�3 ��)W_�j��}��������jkG*giI5]l6*M��T!_��ˣ>�C~vS��1�G�|�w��M��"i��664�}�_�����A��[�j�`�X!1%��V��i��[������k�U�Z(�$�>;�SS3������,�����a`U�T�4Ć�
G�R���D^�ؽN�%d)̯O(�9���ό�Z,�������2gٯ�=�r���s���L�e(0�L�Lr�͙:��uڌi�M�2�)���B�50ÕT��^o~��yzO��q=��K�'�X9���|���5��S�d2ԗYh�([��V���cD�fsn�V2�o ���2�r��u���6�YsH����Wp�!!�X�LK�8a��i3�?�;�"�bF�������ɓeRK�h��ڱ}�����mԂa`Hu*ƺ�R�,���T�0�@T�u�bALK?o(*�M��xߒ5x;c25�!��^R{{��+W>X�m{EgGG*Gs�1,�R]�r���x�௨�����|�l6�B}�J�+�IRZ��\���yr灚)���l�v��$(*p4:���Llk�hdR)Ɔ�
yo��lK.)��,.�SRjh���$p���:�~r�[+W޽~Æ��λ�5M��r��-���x�Q/U�S5{�̧v�@�O�<�i��$�=�����s��,���a��N���&�i�)
�����EB�T�d�����"p��'-C��g+�m<x���P�p�R/OUU���e�7޼k��}�m'O%q�ެ����t��n'�OG���2g�l6U��g�p%a����{���64���hoK�� ���2�j4R����BѠ	z���w���1@�EH����^Z����V}r�QZԷ����T���oS��z��U�֏�IV���b��ǃU�Z����o���_:�� !����.\eٮx���S�+z��w�x~�ԩA�_b�6�_*�T��v{/��T 4����.=�+1/�X°�����ͼ�QC��~�����h�|���{��Ѣn�۪��-���T��f�	D�(��l�w�:��]�B��5�����hj-��4fP�]i���W"20��O4��N� �=m4��i$��e�xtV��X��XP����x�`k��b�:��mX�~qu���,��X�&&�@o��+U��O?�z޼�~d�Zp�*�����UU�-Z���j�$͂^	Ao�V��a(��
ȱ~����>U��0Қ^��Ϝ��Ct��h�����.����T�|k��I7(kH|��Q=�Ə�:mʔ�l	���B_җ
W5*��M��ZZ&�<t8ˀH��2�B$6��hPt��nsFV�a�c���*�fkfL���>��4MӅ��dR���u�*,*zỏ=2js���՝?�`���Y�0M8�
!t�.6\���$uuwN:�~bLWKK�QQ�V�A��1p�AE���*�I�zWb�i��z[a�:19i?�ہ��"�������R `HKO��t��?�\��Ӧ�8=#cwNn�ZQ�?!���pe{zz+�vt\�h��iJ8])'J�F���\���)�]���t�Y�u��u�-��u�/e���4$I��и��ӓ����?3k�
���/��NԷ/){B�+�w�(�TI
��A�Pȡ(�%��h3�ͫx��!����9�sm�K������UU]^�����c�����rr��=�0L ��eĒ �@B�{i�Fq<�f��fY����_�'�Y����F566.>}�t���A�1�_
�P!t���=�9O�tɥXP^U[����[>����7)77wOVV�+�(�~��Œ ZW1��<yyy"���O�"���������RU�H��pE���!���+B�W���!�0\B�`�"�P?�pE�~��B� �!���+B�����?*�9�	    IEND�B`�PK
     D"BYW���  /   images/19f08d4b-a68c-4e36-96dd-32682874608f.png�PNG

   IHDR  �  	�   yT�   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{��w]����g&�6�|h9h+G+���.�x�TtE���E]+M&PquGݥb���tfR��b@)��ߺ��˅��Ρm&iB���4��=������A�=$�{�s����������H�E^���                                                                                                                   ��J�`zz���{�����3K�  �������kKw  ��f��?��?����,�;E�޽��F��w�y�ו�   ��p�رۏ9��7�7��na��Jпv��Q����HD���-    ��r�[GGG�t+��N1g�y�_��m�    X%���G��ǿ�t+��N����J)�N�    XerΟ{~����Ϊ���|sD��t    rFD\��~�ɥCh/�;�jbb��"�C��    ��e�cǎ��!��ѓU399����U��t    t��:t�������Uq���?-"���g�n   �������t�apg�]s�5k����(�    �O����Z:��3���r�iÆ�9���-    СR�������t�cpgEMMM�?"~�t    t�����^z�//��3��b���~3"6��    �.�Z����۷?�t'��Ί����ɜ�%�;    ��|{UU�����O)3��v���ߛR���(�    ]��F�ov��Q/1��V�]w�s#�Sqj�    �b?u��!'Ht�;ms�uם600puD<�t    �s����Q:��gp�-&''�6"��t    ��?����;˖sN�=��#�[    ���RJ=::���!<1�;�6555�V�    zԺ�ҕ�����t���βLLL�RD�a�    �qOO)}���ꯞQ:��fp�MLL���#"�n   �>������ݺu��!<:�;'ezz��)�OF���    �JRJ?044t��Ȉm��I�MNN�^U�����-    �oRJg�~��Z��oep�LNN���+"��J�    @{����o����9n;v�G�G#��J�    @��9o����3�;��/x��G�ϔ�     ""��R��������k�����w��c�    �l�9�K.y^������7��.(�    <�3>��~�ɥC�����511�}��k    :���nǎC�C����411qVJ����t    ��^���m�#����Gu���?-��وxf�    ����666������η��k�\�Q�    8a�e||���#����o�sN6l�@��_�n    NJ�9_6::�oJ���;�`jj�}�˥;    �eJ)��^���!����?������.�    �œj�ڕ۷oV�~ap'""&&&~"���    �[ά���/����!���NLNN~oJiGD�n    ��ǎ�؎;�Cz�����t�Mω�OEĩ�[    ���Rz�C�����u�>v�uם���tuD<�t    ���1>>�{�#z���OMNN|""��t    �:r�����\�^ep�C9��#��[    �UUK)�����kJ��"�{������k�;    �"֥�����^X:��������/����t    P��[�֧/�첧��%�>r�7�PJ��J�     Žxii銭[��)�+�}bzz���Z��7    )�X�f͇~�#�dp�����WUuuD<�t    �q~q||�OKG��{����\���o+�    t�?��������v��Q���F���n    :�����+���=�/x��G�ϔ�     ��@�������S:�[�{������,�    t�9��\r�%�+ҍ�=hbb�r��-�    t�3�{R�ncp�17�pëRJ?�    ��{y��oFFFJ�t�l���8�V�]�K�     �-��cg�q�h�nbp��_��RJ���g�n    zC��m���_��[�{�5�\��^�*"��t    �[r��u||���;������ӆ.��זn    zR�9_�}��.���]nrr��w�;    ��6TU�Ƿm����!����Ŧ��~#���t    ��Z��?�}��g��T�.511�9�m�;    ��rfUUW]~�委�D�.499��)�1P�    �;�<v���v��Q/�i�]榛nzND|*"N-�    ����:�������E���Ӗ������n    ��yccc疎�$�.1999800������-     �x||�gKGt
�{�9����7�n    x�Z��#۷ou�N`p������t    ��XWUէ/���)����&&&ޒs�ϥ;     ��[�֧�m����!%�;�7��C)�ED*�    �^\�ׯغu��!��;����Kj��'#�oq    ]�׬Y���K�w��nxv������~    t�_ܾ}����(���a����u�Z튈���-     '#���FGG�^�c��;Ȏ;�CCC���/�    �)��ccc?Z�c5�;�Yg�uqD��t    @F�'FGG��t�j1�w��������     m�!�t�%�\��!����&&&~!".,�    ���zll�I�CV����n��U)���    �w�<">6222P:d%y���8�V�]�K�     ��?�3FKG�$�{!�_��RJWG�3K�     ���������/ݱR�\s�5k�����-     ��=����R:b%�WY�9mذᲈx]�    �RJ�ccc�/�n�U6==�ވ�w�;     
��Ol۶��N1������_�9��t    @xj�^����۟U:�]�dbb�'"���     �̪������O)��U099��)���[     :�+�;��;v�K�,��}��t�Mω��#�I�[     :QJ鍇~_��2���뮻���D�sK�     t���Ʊ��sKw,��}�LNN|""��t    @��xll�M�#N��}�l��7��     �"�������_]:�d�W����E��Kw     t�uUU]y�e���tȉ2������["b�t    @{F�պr۶mO)r"�m4==��)�ED*�    ��^R�ׯغu��!����&SSS/��ꊈ蚟|    ���k֬�Pι+r6������3r�WFDW}{    @x������8�e���k�UUueDt��     ]�GGG�^:�ܗ!�\�hD��t    @/K)m������SSSo*�    �#�����]:��O����ƈ���     }dCJ�3�\r��J�<��I�����x_�    �>��������ƞT:��O�7����"�^�    �O�<">6222P:��'���?�V�}:"֗n    �s?~��_Z:�����k�}j�^�lD<�t     �룣��*�u��{���ODċJ�     ��RJ����J����9�cǎ} "^_�    �o�RJ+��ܟ����)����     �PD||۶mEO)1�?�����EDǜ�    �czZ�^�쥗^��R��055��)���     �3k��Uccc�K����(&&&^�s�XD�n    ���*">�cǎ�j����M����H)]O*�    �I��C�]��75�?��?��UU]�+�    ��l��ռ���a����k׮�DD|w�     �/���cccoZ�����ֈ���     �M-">�}��W��������F��Kw     �v몪�rll�+}���'&&�\�    �����m۞��7���}zz�SJ��T�    ���z�~�֭[׬��vp���zIUUWDĊ��    @G��5k�|(�"a���>==�������>     @�y�����J\���k��v]UUWF�K�     ��RJ4>>���}ݾ�sε����DīK�     PN�y|tt��f_�SSSG�ϖ�     �����'�o��]�`���EĹ�;     ��UUu���۟ێ����>55�Ɣ��Kw     �q�SUՕ�\rɩ˽P����ӯ�9,"�[     �H�r```�����r.�Ӄ���_fUUWE�)�[     �h?q��_�����~��>�^�6"�U�    ����ccc�<�/���}���CCCC���n    ���w||�ߝ�����sNǎ�@D�p�     �N�9_v饗��D����������~�t     ]km�V�Զm�N����'&&���     ��=�^�_}饗>�x��g����O)���     �g�U�ծ[<��������s�����-     ��W��><22�{z�����g�����'�n    ������~��O�y]=����PU����-     ���������>��VL�MNNF�U�[X�V�7�|�RJɑ@    ��z�������~�&��s������z�v��-"~�t˷k׮8x�`�    XQ�֭��Ϝ��c���s������<Rfrr�?���'�߿��   @_����V�U:��[W\v�e�����}jj�#�OJw�|w�}w�s�=�3    `U�c~~>rΥSX�g�Z���m���G�`W�SSS?�s�pt�Q8|�<��v[�    XUUUűcǌ���z��[�n]����}rr��9�+"b�~2mvv6����T    �KUUE�Ѱ���Z�v�s�)"�^��xLNN>="�WD<�t�3??7�|s,--�N   �brΑs����SSSq�UW��?���k�]744����-,���bLOOG��(�    a͚5144T:���)����G��kCCC	c{׫�*fff��    ��f3Kg�|)�<�у������;X�}��ő#GJg    @�i6��j�Jg�|�;�OMM�#"�-����z�q����    Бr��h4����),SG�4ujj�9翊����Ͻ����~{�    �xKKK188)u��7y7�OOO�2�|UD�)���<����gϞ�    �5��ݭ��믿�̔�?D�SJ��<���133��`    �䜣��,��I�#[���ڧ����#�Y�[X�f��v��    8	KKK1??_:���O��޽{(����xU����j��7��F�t
    t���"��zGL���O������e�å[X��s�ڵ+�=Z:    �^�ٌ������������9��t˷o߾8t�P�    ��F���]���>11������w����    �9�F#��*��q(v ���ԏE�G���gy������Kg    @�j�Z188)��)<�"��7���g#b}���>��ݻwGιt
    ���sTU����Sx�>�OOO��;"���������b�Νΐ   �UPUU�c``�t
�aU�s���?�����D��V����B���xK2    �����h6��3x�6�_s�5k׮�xD|�jݓ��j�bff&���K�    @�YXX�����<�U�7lذ5"~l����ٳgO��Ζ�    ���l6�>сVep��������ո+k���q����    �����_�ì�KS���~1".�����be�}��q�w��     �j�b`` R2�v�ܧ��~ ��wᵹ]��/~�3    �G�9G�Պ��A�{X�#e���^�s�ۈX�R�`u����޽{#�\:    �&UUE�Ѱ�u�y�}rr��qMD<o%��ꙟ���o��    ���#�)��O�_{��r�WF��}mV���b�|�ͱ��P:    x�������>�mI)����euUU333�h4J�     ǩ�l���b錾�g����d��۷/�9R:    8A����j�Jg��{i*���[o���     NR�ш��Jg��;���{ﾻt    �9�8v�X�K���;���������     � ��F�辊�DD���l�޽�o>    �!�V+���Kg��;�l6c׮]^�     =hii��J�}��j���L4���)    �
Y\\�����=����rαk׮8z�h�    `�5��XZZ*����}l߾}q�С�    �*i4��^A�>u�w����_:    Xe�F#��*�ѓ�}�+_�J�q��3    �r��h4"�\:������Çc�޽�3    ���������=���G���b׮]�]    ���%�{������B���x1    �O��l����>�j�bff��V    �baa!Jg��{سgO��Ζ�     :T��t:F�{���������3    �7??�V�tFW3�����;���    @�9���|TUU:�k�{�<��v[�    ��TU�F#rΥS��������޽{��     N�����{L�ш��g-    '��jE��,��u�=dqq1v���S    �.���hk<A�QUU���D��(�    �f�����3����G�۷/�9R:    �1���>N�p뭷ƁJg     =��hDUU�3:�����{�q��w��     zX�9�;9��)����|��ؿ�    �䜣�h����K�����ݻ��    VM�Պ������ޅ��f�ڵˋ
    �U���dt�.�j�b�Ν�l6K�     }jqq1Jgt�{�9Ǯ]�bnn�t
    ���f,--���(�.�o߾8t�P�    ���h4��~�{���;����/�    ��FTUU:�#ܻ���;�(�    �-r��h4"�\:�8�{�;|�p�۷�t    �c��*���Kggp�`sss�k�.ߎ    t�������jaa!fff��    �������P:��{j�Z133��    t�f�ٷ�����ٳ'fggKg     ��f�ٗ�w�;���������3     �e~~>Z�V�Uep� w�}w�s�=�3     �-����QUU�Ucp�<�@�v�m�3     ڦ��h4�s.��*�`vv6����7��    ���O�����F�333}w�    �?Z�V4���+��^���b�ܹ3J�     ����Ş�B�TU333�h4J�     ��f�����3V����}��ő#GJg     ������=b��^����(�    PD�ш��Jg���}��{�q��w��     (&�ǎ��s锶2���|0���_:    ���s4����dvv6v���S�x     ���j���|錶1���f��v���     ��������+��j�Ν;��l�N    �H������P:c��+(��v특���)     ��l���R�e1���}��šC�Jg     t�F���Gs�W�w����    ���h4����'��8w�qG�    ���s�F�9��)'���f��}����     �ZUU���|׍��6����]�vu�;     t����h6��3N���Mbff��ߢ    �)caa�t�q3��A�Պ������/�    �S��f׌��6سgO��Ζ�     �I�f�+N1�/���������3     z���|�Z�����w�uW�s�=�3     z^�9��磪��)���~�x������Kg     􍪪��hDιtʣ2������ػwo���    ��N��'��h���Lǟ    ЫZ�V4������~c�Ν���P:    ��-..v�Vkp?NUU���L4��)     DD�ٌ�����d�t@7�9�-��G�)�  �u$"y>�)1T��n^�    IDAT  �m~~>j�Z����)��q�m����Kg  �{�"b6"G�lJi���ٔ�lJ�pUU�1[�Վ朏���f��FDDJi�V��~��9�f��<��o6�s###��}�[�n=mnn��f͚�Rz��?VU�@�y�#�����P��6�O�9o��jO�9o�9����o���DĆ�8����  �F�F#֯_�Z�C]R�/899�ɈxS��[�=�����/� @wX���Dā���q "�O)=�s>P���_ZZz```ࡍ7��y�\p�S�Ϯ�jϨ��Y�Z��9�gDĳ"��9�g���O-[ @7��j�~��H���q3�?��Ʈ]�Jg  P^�F�q{D���~UUj�����~���P��5222t�i�=#��̈8=�����3k��ss�gFķ?��'� �\�^�u����avv6n��h�ZO��  �Cq[DܖR�-�|[����ҽG��322r�.@Y\p�S֬YsF��:=�tVJ鬜�YqVD� "���  �ĺu�����(���czz:���K  :_+�6��{s�_�9�Q���8r��]'r�9��=�y����V�}{D��RzQ��%�xZ�:  �ipp0֮]���5��V����177W: ���wG�-)��qK�y���y<\p�S�J)�,"^�s~YD�4"Ό�s  +o͚5144���4�?BUU�s��8|�p�  ��lD썯�{j�ڞ��-�}�so?�쳝H[����}���ЋZ���RJ/����/���u  <��k���������{���￿t  �j6��3"�"b*�4u�ȑ=###U�0��%�\rj�����xED�4�����"bu� �	�_�>����������o�=����  DI)̈́q�.3222t�i�����+�kC�+��  奔b���Q���7(�#����gϞ�  �ȸNO�����o�_k
� ��Z��ׯ��V��<}?�>|8v��U��t  �ྈ�|D|!">�������������z���_�Rz]D�."�\� ���ڵkWtt���}nn.n���XZZ*� Ыn��ϥ��PU��ټy�����ر���/��UU�6"~$���SJ�(� Ћc�ڵ+v���bzz:���K�  􊥈�9���|����w���_-���/>�����__{����  zŚ5kbhhe^�ӗ�{�Պo�1�=Z: ��-F�RJ�k�Z�x�ر���O3�
�袋��j�~ "�uJ�G#���M  �l�ڵ188������>33_����  N�׏������ߟ����~t����j�~$"~$"~4"�T8	 ��[�.�z;������sO� �n1���s)�O�R:�F;v��u�]ߓs��Z���9��DD�t @�K)źu�^���m���:yp�뮻��n+� �ɪ��1�����>777��###����e˖���^�s����Ɉxn�& �NU��bݺuQ���y��ܿ�Ğ={"�\: ���9�V�]�l6?�E��;r�颋.���󏥔���� �U�^���׷�Z�=��C���ƾ}���  �9?�R��r������b�ޔR�q�������2���xCD�) �Z�V;v,֭[)-���½�h���t,..�N (���ҧs�?z��###U� ��������rʿI)�9"~&"N+� P���`�]�vY����}qq1�����h�N (喜��~��T��3����=�S^��KWώ�g�n (a͚5144t�_߳�{UUq��7�C=T: `5�"�s�W�Z�+�?���J�eǎ�/�˯�9�)�������M  �i�ڵ188xR_ۓ�{�9v��,� ��n�9_�s��;����K� �c˖-�H)�j��-���=  �a���Q��O��zrp�җ�_��K&  ���SJ]ZZ�����}�c�޶cǎ��w����үF��E�)��  VJJ)֯_�Z�ľ��!��{�7���/��= �J;W�/�_)�\:�?]tѺ��sο?��  �-���rJ�t�3zO�>�`���D���	 �����\J�����O���,���/���z���қsί-� �N�z=֭[wܣ{��q�M7E��Z�[ ��*"�w���׬Y��{��A O䢋.zYUU��R����K�  ����@�[��>�'���������{ ]�@J�C�Zm���λ�t����r�)?�R���ڟK7 ,���`�]��	?���V����177�Z� h���"�/N=��+�9���= �r��������)��Gķ�� 8Yk֬���������sαs��8t��j� ��E��k��֍7�.������/Z �кu�b`��oLW�{���ƭ  �i*"�k��۸qc�t�j���Ϩ�joM)�VD|[� ��~���������o������;W�6  �r8"v��r��ͻJ� tO� �(��ׯ�Z���k��Vcp���b߾}+y �v�)�t����ߜ{���1 ���/������I)�FD<�t ���j�~��H�'���>;w�V�  ˖R�BUU_�Rʥ{ �Ņ^��^����8/7 t����X�v�7��]5����ō7�KKK+qy ��Z����9�ϱ1 ���q3?�R���xM� �G388k׮����}aa!���c~~�ݗ X��)����r�ƍ����5[�lyED�^D�rD<��  
Y�fMED��V+n���8z�h;/ �\�F�_=zt���ȱ�1 ��}�{�����9�E�)�{  ���{W�333�կ~��� 8i)�/D�_<�y�����>�U��߼���}����������9  �nݺ�������w_�. ��M)�ɦM��+@�֭[�,,,�-"Ώ��� �[J�����+n��v\
 `9>�s�O�7o��t �jdddhÆo�9�QD��t п:vp���[n��s�  N��j��lܸ��! <������G���� (�#��z(n��横�MU  '����1��aD��t �?:npo41==���m� 8.���wO�`�� �j��}qq1n���8v�X��  ��������1�{UUq��7�C=��$ �G�R���8ӦM7�n`卍�����?1�� zPG�9�ؽ{w<x��9  �斔һ6m�tU� V�����SN9�wSJ�J�  ��#�/}�K��/��)  �있���?��8��[�c (k˖-OO)�a���#b�t ������{o|�_lw �#M)]�v����;��;GK� �Y.������?��7�n �[���������9�;  "b1">800�G�x�;��������M�V{����[ ��Tlp�����n�)Z-�� �����ۼy��! t��s�袋~!�|AD��t �]��Q7??333�v `%\WU��;���/�����rD||�֭W.,,�ǈxwD<�p �%j�}�V�333����ڷ zۃ�G�����r�{�����?[\\|aJikDT�� �η�G��c�Νq�Сv� �_UD|$"6,@oڲe�+"b[D|_� �s���{��5� m�R��9�����_5��������=���8'"*� t�U{����o�;Ｓݷ ���y�����}��^
��z�����Z������X�?W �kU���/�����[ �'G�_眇7o����1 ��-[��`D\//� t��>;w�~ `YvVU��^�
@'������ӈ�P� (kE�p����]�v����9��ѣG_el�Ӝs�9�����j�^��t P֊=ᾰ����1??��[  ����~cӦMw����g�g?�s���n Vߊ<��j�b�Ν�v �d��s6m���v �ɦM�����/����- ��k��W�ڵ�g��կ��� @H)�}D����n�iw �?m�?�������� zޑ�شiӦ��r� h����=O�ˈ���- ��k��}��{z���}] �w���~qq�7�?���J� �Jx����S)��8�t �rV�w ��t$"�ٸq���e�7o�L�^Y8� z�� (�.--}����#d ��w�����sr�o��{K�  �gp V[#"~kӦM?�v ���͛?ߝR�d� ��� ���9��9�zxxx�S� ����მ6m���ү����� ��� ����ڼy���! �)6m�ty��U1S� X>�; �ҎD�/���͛�J� @���V�}Jik� `y� ���9OVU�������t t��766m��{��8\� 89w `%��ֹ��׾�Ｕt t����O���וn N�� h���)�7nڴ��FFFJ� @�9���8z����8"��= ��K������}衇No�u����V��z׻�- �`˖-o���#�٥[ �'�	w �����ѣG�`l�����V�U� �
�p ��HD������C �Wmݺu�����r��n �'�����ol��u��67m��{)������� �� 8Y�9�rxxxo� ��6m��x]D�^� �Vw �D�RJ����i���s�c ��lڴ�ơ���O)���- �72� '�h���7mڴ�t ��s�=�������KJ�  ��KS��u[�V��7n�]: �g[�l�����>P� ��'��'�R�B��5�v �<����UU�TD.� ��� <��:��S_�ٻ�(�ϻ���g�=3��v;7M�p)q(�J遐BI�S)�$P�q���43����L�M
N�`zh���.�Pc�#M-�P�Ĳ_%ۺے�����?,%�"ٺ��Ͼ�^ky9�e���3��G�off�`� �̮����z�u�a� P�� 8��s�<==�cW_}u�t ��6n�x����7����t �*�; p&�)�����T�C �s��?��O?~����t �"�; p�#9�255�;�C ��WU�������n-� ��� �jwD�nff棥C ��R�SSS7DĦ�ȥ{ `T�����9ߛR������J�  kczz��r�?�� =`p ""�*��-SSS�� �����I)}gD/� ��� ̶��7NOO. t���Ԏ������ ��� #,��;�^z�?����x�!7==���x�t +�; ����m?|��W�� F������x}D<T� ��� F�6m�tuUU��! @oMOO������n�acp��R�uzz���R.� ��q��}�F��"ⓥ[ `��`���n�����t P�;����f�G�_�n�aap��s��� ��]�zבf����- 0� 0�=33sk� ����]�:R���]� �� �\J�=���?[� �_7n<Z��ߔs��t 2�; ��R555us� ��mܸ�h��zS�^ .�� �׿����\: �z׻�D�wD�=�[ `�`8�����# ��3==}8���q� 4w >�=??m� `p���l�ZoJ)�)� ��� ��������N� `��p�{"��#�@� w )�����?PUU�t 0���>S����J� � 0���9߽nݺ���kWJ�  �eӦMw眿'"|� ��� ��ᱱ�7_s�5�C ��433�є�G�k� �Y�`�N)}�;��Nw� ]555�{q]� �gw P)�Ŝ�wOMM}�t 0���!"~�t �+�; �vD|����/ �������p� �Gw L���n/ ����:���o���Q� ��� �oLOO��t 0���Z�t:�gJiO� �'w  )�����?Q� ��۟R���t� �w 9�{k�ڿ���U�  "bӦM�DĿ�g�/ #�� ��F���7- p����?���.� ��� ��?�q�ƇK�  ������"��Jw @iw �s9�>qr �/��r�V��)��)� %������pzz��Kw  <�M�6-�j�å[ ��; ��O�[��m)�\: �\lܸ�ш���U F�� ��|�^�5�\3_: �|LOOo�9�l� (�� }(��7n��t ��XXX�w�� �^3�@�������) p�����("��n�^2�@�d�V�T: �b�����j?�s`�����j߷iӦ��!  kaӦMK)m.� �bp����6m��`� ��t����F�GKw @/���zz��Kw  ����:�v��q�t t�� �{�^���t @�\������.� �fp��:9�޴i�S�C  �ijj��)��R� ��� e�������#  z��l�dD�.� �bp�r����  �r�7<�s�шȥ[ �� PF�V��pUU˥C  z���t t�� �xߦM���t @	9�M�p� Xkw �����7��  (efff!��o��2 �; �V'��#�� F����Δ�o�� ��dp�J)}`ff�/Kw  �f�9�Jw �Z1�@���j�. �/n�ᆧ#b�t ��; �HJ�ڍ7-� �O���?�s��t ��; �@��������  �G�F㚈X(� �� ݷ?Y: �_mܸ�є�ϕ� ��ep��{����#�#  �������� ��ap��z<���#  �]UU�q]� �w 袜���̌�H �����EĶ� p�� �=wMOO{P* �y���#�Y� .�� ����tޑRʥC  �ƍ�M)}�t \�; t�o_w�u[: `�7Gı� p�� ���[��{JG  ������� p�� ����7�) 0�j��/D��; �|�`m��j���  t�6mZ�9o)� ��� k��6m��T� �a����q_� 8Ww X;�ׯ_���  â��V���� p�� �FRJ?w�5�̗�  &�5">]� ΅� ����Ǐ�Z� �aSUU'���� p.� �rηVU�X� `-,,l��O�� ��bp����^��t ������Rr���gp���K�6mZ* 0̎?��x�t <�; \�c�z��KG  ����t <�; \�_۸q���  �`ll�?Eľ� pVw �p+�v��KG  ��k��v%���� p6w �p�{����- 0J�Ư��Kw �������|�t ��ٸq��<��O�� �31��h���l6�t ���ضm�ʗ����; �L� pVWW#"���-[��t �(���S�&&�]zi� �w 8O9�h����t�+� 02fgg�����x�^T6 ��� �����������*� 0Jj?""�w�e111Q� >�� �S��:�����.� 02�m۶!E�ĩ?��+�(� gdp���j�"�|��`UU� �Ec�����S��/��R�" �Bw 8��n?i,"n�q
 ����G>2�"���9�F#�w�e%� ��� p�r�g�#"~��o��^�  ��K&'2"^r��{�ke �#w 8G�f��~��n��ի �Q�m۶)癳��e�^ccc�L��2��9�9?��񶪪��=  �b�V�����|J)�x�z� gep�s�s>��ROW����  `$�u�]��Z��O�µ2 �	�; ��s8�~�nٲ��l ͕��"�=ׯ[71�׭�E <+�; ��gyX��R��y_7[  F������y����]+@0��sh���r�̩�����ԭ �Q�i4���p����@?0��s8���z_UU�� \��;w�����{���c��d�� �� �9�������[׺ `�N�ֈh���{��߅ 8ww x�v��o���[n��yk� 0�vn��m�=�{��<�zP�� ��^'s�K���z�Z  ����\#�j�t��bb"֭[��I p^�e�n�    IDAT �,.rp��x��7���֢ `���D�߿��p���� p�N'r��2��v�֢ `��q��GĻ/�u� �dp��X���'}WUUo^� F�cc�D��:&'clll� ����,�pp������.Y� ;w���������.�ķ] �ap���t:k�r/����� ����F�t>��p�x�e���K�y1�����n���-[�|]7^ ``u:�G�׬�K^v�k�r p�� pk|��I�N����[�ֻ��  �fnn�����u�FL�_��/ ��� gХ�="�v��uM�^ `P�S�۷EĆn���N�P�� N�s��s7���n���/��  ��������xc�^�2N� �; ��K���j��n����| FҎ;^���{l�Е�� �|����`p��x]J��2 ���9�Z������R��c�{��1�; ��G�{�o����z�f  }��U2���u�S� ��� N��tz�V��[�n��� J�ضm7E�|����@����:�~���{�7��M z���Z����qY���N��� p��{䜫-[�|c�� �������)r~C/�s|l,���z�� �8�; ����ɜ���t>t뭷v��a  ��m���)����� ��� NQ��	_����� �[�m۶!�j��"G�7��!�; ��s��sɄ߼y�*  ���j�_�_Q��'''K�5 #�� '�N�������,� ��v����[K6L:�@���~�#⒈������> mn۶�J9�r������3 w 8������ǎ��JG  \����K�^ߚ#��>���֕N `D����������s Un�>�*�q���^1�@<3��ɕ2��s����ה�  8���w����tw z�� '��	�����UU��t ��رc��"��P��tN��+w ��y`꙼<"~w�֭�� ����qǕ����1^��t�� �� �����7�ڵ뽥#  �fnnn]�������t˙���EJ�t #�� ї�ɜ�͛7���  g�n�j���3�&E��x��`� ���{DD�9�����a� �S}��;g"�GJw<�	�; =`p���="b]D�aUU/+ �s���S������@/� �J��^��r�-�+ ����ۿ6u:��pwW� �w ���#"^�����[�n�� �𙛛{i�j��n9Wccc� w Fހ��'}�]�~�t 0z�m۶!��?���S��|���; #o@���k����t 0:�n�Z��?�P��|�5� w Fހ<0�lnټy���  �_�9����="��t˅p��^0��`K9�۪�zS� `���ر9G�h�Uo4"�T:�!gp`��2'�Eć�l��u�C ��sv��)�ݥ;.F���ke �2�; #o����:�ζ�o��U�C ��27;��)�WJw��z�@w�J����="�E�v{{UU�( ����7F����8^w��.3�0�hp����������� �ܝw�È�È�(ݲV�p��|����e�����K�  �ivv��#��#��-k�fp��|�`��	���~D�^U�e�C ���;�|U#�ΈxA閵桩 t����7��{D�7F�Fw �\���~ENi6G��tK78�@��J ��Eğ�z뭗� ��Ƕo��F�\����-ݒR*� ��3���{����Fw �l>�}��wj���#"jw ��� ��uKKKRU�P=� �xsss_֩��"�K�t���.3�0����}KD쬪���! @�۶�+���h�������� 0Z�!"ꅥC ��fgg��z}g���ap��� 0z^��j��h �n�Ν��G|<"�,� ��� ��U1WU՗� zk��;__�tvF��[znt���; ������n���W: 荹������n)a���@!w m/o���e˖T: 讝w�������tK)�; ]fp .�t:wn޼��� �cnǎ)�vD��n)�	w �����K)�N�r�\U�� ��܎�G��O6 w��u�� '�Gć����t p����s���9�R��_�R�n3�0�p�<���媪~��*�' ������$��?��+��O��v� ��� ��\�_U�d� ��|��;�L���"�J���v�S:�!gp`�9�~V�s�}�{_R: 87s۶}U���9�5�[�Q�	w �����3�?��l6���o~U� ��}tv�ۣ^�+G��tK�r��n3� ���v�/�����! ��휝}{��o��-��� t����W��rx.��?ؼy���C �ϙ��k�ܱ��N����=���j�N `�Y �sU�9�RUՇ��ZW: F�w�qyj�����Q�e䜝p��� �<'���Fĝ�
 ��m��U�����Z�eP4���	 �  #�CS/�����lٲ���Q�s���>�p�W�n$���� �<����N��q��@olݺ�>7;{K�t�(<���:�@4J @i���8q��WE��UU-��a4;;{E=�w#��K�*'��'� ��k��"��UU��t ���ۿ��7al�(���� w ��ymD��͛7� 9�47;�SQ�ݕ#^V�gЭ��5_n��O?���k�� �M+++�t��Z���xGUU>�����{a�ۿo.�2,����_X(���s� �	�.x{D�yUU�, �f���o�v�o�ؾ��p�� ��/�]����UU}o� UU��v�>�j;"�K������@O4J @?0�w���UU���~bff����3���}I#���9��t�0r��^�. @�R�޺��p��-[��t �����~{=�osJ��.Y^^.� ��p� ��=�9��)��+;��_VU��#bKUU��A P���\#Z��:�N�uՒ��� Np�LO�E��Dğ������) ��m����n��H�g����; ��: �`p�7�Z�OWU���p� #������ٷG�~w<�qz�	w zŕ2 p����.��VU�}�o���S: �iǎ_Z�����R�eԬ���N `DX ��{1o��O9���:y�����2�����rt:@o8� '܋r����T{y��� !� 8!�dt/�iw ��S��c��@9� ���j��qyN�0Мj�/KK� !���)��z�>�M�ɪ�~<�v` lݺ�>�c�t-�O��ǒ��2��)\)�w��UU�W[�l���1 p6;v�x͋^��?����K���%L��\) �p½o}}������>ﮪ�X�  ����?���WV���5��o$����B� F�c| p���V#"������z[�f��r�i�w����r_~�등���ϗN `Ĭ���n�m��O?}�Z�. ����j������}�V�]�����! ���;w~Mj�%R���-<�O�sO�6��3 !���ӸVf`�����Ϫ�~5"n���6 �j۶m���wG�3)�<��VWW�� ���3 �q��@�Ͽf ��;v���z�ވ�>^�o��$ �iRJQ�բ��N��}qD�窪�שׁ���A ���y�rJ�O��[K�p~�?^:�dp�3������]񦪪~sll�=7�x��A ����+�3��wF�D���q�; xh* �A�ݎ����\������.���M�6�_& ��#���%����+�ÅY^^�{t #�%� p�z=RZ�?���.���9v��g��z�֭[=�������;�����o	c�@{�ر�	 �(�; �����/���ڵ듛7o���1 �����7�����D�ykD��t���|� F�;��,�F�������r�RU�lD�TU���� (kvv��zĭ���-��N��w 
1��Y4�XYY)���{cD|���ߏ�몪z�p =677�%��~w����p�ؐ9>?�N�t #�CS�Y,..��6�#�����:\:������t��S��tݱ�����O�� `D��Y������j��o!"�cD�\UU�K� ��fgg�����H�"���{����h6��S Qw x�N'Kg�;����n��������2��3"�W���_X��x�t #�� �aaa!rΥ3�-�;� 3�������� `���9�Vf�-F�oDĭUU�-��3��]�|�@Qw x��!"V"�?G�f�;@�1�1??�?�`� F�� ����bt:������h4~�nz�t��۶mۋ'����qI������q���� �8�; ���p�ND�ﭪ���5sss_���wDď���=����OG��*���3��9�9���B��ӟ��~�U�z���-oi��fsw���H�ڈ��Q/�C�8v�X<��å3 �� �jii)�m{*g�PJ��9�۪�r�?������~�{s�3)}c���#�w�SG���  �; ��f�+++�3��#�?6���t�MO��T��~�e����u�ؔ#^V����n�����y; ��; ������	�Ո�������>]:`P��ͽ"��WG��K���>{�t D�� ����qq�rD��ꪫ��=� g�~v.Խ���KK�3  "� p^��v,�@ǅ���h4~���n�]:���o���u��?�"~2"��t�giy9v�w_� �,�; ���s,..Fιt
��;SJ��s�ê���	`��ܹ�N��9�_EĆ�=�Ǟx":T: >�� �iuu5VWWKg0<���߉�TU��t@��r���F�ו�a�u:���=�D��6 ��� �S�9Jg0|�1�R��W��U�w`X�r��#��=K������D��,���z8"n��7�x��1 �knnn]n��RK�r�kJ�0�v�w_,-/�� ��cp���tbqq�tï�="~+"�kUU�
� �UUU�7|�7�.����/#���M�����,� _�� hiiɝ���rD̦�~+���WU�A@_عs�S��ֈx[D�,HO<��q���� �� p�Z�V,�k̔q$"�$"~����� #�c۶��N���#�G"�k�0bVWW�S�v�� �32���9���Rt:��)��=��z�7���w�_:^sss�ϭ�w����]�<	�b�c���'�,� gdp����;}�"�C�F��o��'J� �onnn]�t�Y��_����㥛m�V+>�k� �-�; \�����ٍ��]���ZU��w���|�#��NN~[����ZJߓ#.+�'=�wo�?x�t ��� .���j��z~%}��x���WU����w�4���W�r�����GķG�D�&8]�ݎO���� �5�; \��s,..:�Πx,"�4��'/}�K��ꫛ���2v����Z��o����E���<O��[: ��� �@�ٌ����p������R�H��O���/t�Ν;_�r~st:�,Rz]x�)���ħ�'ZN���� �F��΀����="�WU�`�`��ͭK��7���)}Y�&���'��+� ��� k�)w���1�R��9�YU���A�����}e-�)��qi�&�N�0H� ���rgH�#�o#b6"f���ʏ����������5r~cD|G�xY�&XKN�0H� ���rgD<;#b��hl�馛v��Q�u���_�¯M9�������+���n��S�vE��v �� ֘S{#��RJw�����GK�0ٺuk�%/x�W�S���#�[#�y���'�ػ7�<X: Ι� �X�Պ����PҾ��DJ鮔�l����UUuJG�����ǎ;��'N��>"�)"^P�z��lƧ�7:_B w Xc9�XZZ��>�xD�eD�yD�wUU�O����������7Fί���)"^�JwAi���O>�T� 8/w �v�KKK�3�_-G�_�3���E��UU�/�277�%����ZJߔS����U)�V�����r��� p�� �%����j�Jg�����g���'���=�y�=���bm߾�������N絑�k#���<�z(�?^: Λ� �������b�dG"bW��k��'����3��_/-�����O�C�<R: .�� �hee%��f�&�s'��6�|ϕW^���W_����;v�<u:�M�����s~Q�.t9���bee�t
 \�; tQ�9#�\:�Y+"��3���#b׆�����B�2���ۿh�V�*"^�"������Ƹ�q���x|��� p�� �e�V+���Kg���ό�񟬪�`�*����\��n���ҫs�U)�W�_)}mDl(����jŧ�7��v� �`w �����t:�3���Eģ��S��w���Ǫ�Z-�F7�~�����/O)���鼼���M_)�:r�҈+���ݻ�#GJg �E1�@x�*�#��i����RڗRڻ~���\U��n�:~��I=�9�/J�ڕ)�W�W��W戗GD�t'pf�q��� ��fp�� U�x檚}q "Eā�ҁ���_��t:�CW]uա���-�F�[�n�����^��h����Z�ŝ�_�r�2G|qJ���T�9v�w_,{P* C�� =�j9�xf�?ό��O��OE�|J���M)��j��f�xUU�Ū����;|��F���N���KR��̀��S������9�%)�E9�Eх�-@�ػ�ۿ�t �	�; �����HD����>GO���_�9��n������WsΧ^��RZ��h4�����ͭk4�O�����KSJ���������D-�Ɉ�NJ�z��rΗEJ���/��K"��9Ⲉ�4R��ď��"&��4�0XYY�]���@ C�Q:  FI�шF��V�t
0^p�s�s>����/�ҿ���}M���j�֛FJ���g�9���:��?��ǩ������?��I���3�0Tj� `�LLLDJnG  FۡC����Pޞ�3�@���bb
 ��ZY]�'��+� k�� ��Z `��xt�nW� 0�� P��e �Qt�С�_Xx�_ �� ��Z 5+++��`����F�ccc�3  �.�����* ��� 
w� 0������`�����R�[��t @����}�� ��3�@���1>>^: `͵��xtϞ� �w ����Q��Kg  ��ݏ=����3 �'� �G֭[�>w `h<|8�=Z: z�� }�}� ��X\Z�ǟx�t ��� �����A�n��G��s� �)�; �!�� ���={���H2�@�r�; 0��8G�~�t ap�>�R���ח�  8gǎ�'��+� �����j����(� �VWW�ݻKg @Qw �sccc166V: �:�N<���j�J� @Qw  Q��� ��G������ P�O� 0 ֯_�!� @�ٷ9z�t ��; ��Q5� ���ѣ�w��� �7� 0@j�Z�[��t @,..ƣ{��� ��bp�S��cbb�t 0�f<��#��tJ� @_1�� ����� �j�����G��,� }�� jbb"�F� `����G�����) З� 0�֭[�z�t 0"v?�X;~�t �-�; ����G��K: �]�=�D<��S�3 ���t C`����R*� ����C�Jg @�3��H)���x�ȑx��'Jg �@0�����jFw `M=�����=�3 ``�`��j�X�n]� `?~<޽;rΥS ``�`����X�~}� `�-,,ă�<�N�t
 �; �z��; pA��⁇6��0���j4Fw �,--�=�v�t
 $�; 1�; p��WV�3=�V�t
 ,�; 9�; �Db    IDAT�\�WV�3>hl��dp�`t �fyy9���h6��S `��`D���-.-��<�d; ��; ��F��ׯ/� ����xࡇ��� �f� 0b���� F���B���v Xsw AFw ]���ぇ�N�S: ��� FT�^����� @9z4|�ac; t�� FX�V����H)�N ��ɧ��Gv�6�@�`��`��?p ݳ'rΥS `���H)���d�j�5 �a��޽�ľ}�3 `$�T D�3�����^��N �@�9ٽ;<X: FF�t  �?N��+++�l6K�  ��j�C�<��S `���/011�Z-VVVJ�  �ieu5|�X�u z�� ����X��byy�t
 p�����V�U: F�;���j4�~��H)�N ��ѧ���<��� 
2� Ϫ^����d�j�m �~u�Сx�G���N���J �9��brr2�����n�� N�9ǣ{��SG��N �� ��������J4���) 0�V<��#���P: 8�� �������j���R: F���R<��#���Z: 8�� 8occcQ��cii)rΥs `�<u�H�~�1��@2� �V����d,//�� z �{����N ��� \���{����f<���k�>gp .���D���XYYq� �����xx�n� �� ��F��Z-����) k��C��޽�@ �� X3'�uw� \�V����ǎ/� ��; ��N^1���\: α����={��5  �; ��F#6l�KKK���s�s�}ľ��K�  �� tMJ)&''cuu5VWWK� @�Z]]��w���) �E0� ]7>>��+f<� >�ѧ��ݏ=�V�t
 p�� @O����������h�ۥs ��N�O��*� ��; �3)�X�n]4�MW� 0����ݻ=` ��� 詔R�����ؘ�� ���s8x0����5 Bw ���R�_�>��f�������[Z^�G������) @������Ƣ�h8���r� F�� (�iw ��S� 0Z� @�p��a�T; �&�; �W�v`�9� ��� �������뱼��N�t <��s�;p �8�T; �(�; зj�ZLNNF�Պ��� }k~~>v?�x,//�N 
2� }��hD�^����h6��s ೚�f<�o_<��S�S �>`p BJ)&&&bll�53 �#��'�������o �� �@9y�L�ٌ��U�� �s�������c�CQ�����466�F�53 �L�Պ}��C�J�  }�� ����4�XYYq� ]�ԑ#���G��1 ��0� �^����d������j� ����b�y�XXX(�  �; 04���cll�53 \�f�{���O>Y:  w `���f����j�J'0@:�N�?x0<�2 ����T��bݺu�n����s�9ǓO=O���k�fp �����[�V�����G�~:�ػ7�WVJ�  �� ��F��F#��f�T �g���޽q|~�t
 0$� �H����XYY�`U����{��#G��N ��� I�
0z��f�?x0>9��9 �2� #��U;�N4�M'��T�Պ���C�<� �*�; 0�j��gO����� �5�; �	�w��`h J1� ���0�� @iw ��0�C; �/�  ����}uu5Z�V�$ "buu5�<��|2rΥs  �  �V�źu�"��f3VWWK'��ť�8x�P<u䈡 �+w ��R�������n��Ǐ�����ǎ�� 8#�; �E����h�Z�l6��n�N*9�8r�h�;p ���K�  <+�; �h4�h4����`�Z�8x�p:|��O �� `�z����j4���I eye%>��|2:�N� ��bp 肔RLLL|���f��w��p?; 0,�  ]t�V��v4�MW# ��j���Oơ'������9  �� �#�z=��z䜣�j���S��o��^��4=��KJ�ؤI���l1EcOu�A��A���1�_J�ďd
�-�zw�ۦ~� D��뷰U�z�|�&-nn���{7../} ^� ���f���d����zތ�z=�/.�_߽����� �*w �2��v�����������CP�WOp x��ާi��j���C_��L�4���ǻ��M� o�� ������ǩ��je*x������������- �M� ������f�����؎1nnn����8;?�<
 ��� ^��|>NOO����c|_�V���F-��qvq1ޟ�����C_ ��� ^���>M���kZ�V���b�_\���͡� �,	�  /�}��״^�����xv6��C_ ��� ^��}��>M�X�ׇ���L�4������������ ��@p xe����zm��Y���r\^]���Bd �B�; �+6���Ό1��=pX.����Nv ��� ���������l6c�Z�i�L���\.����8??���C_ ��� ި�|>NOO�����ڙ�z���l6�qyu5�����Օ�n ��w  ����8::c�ǽ�o�^�����v\]_����>v �oLp ��{�w�g�'���e��q�X|�b��+H 8� �Ϛ��c>�����1ư~l�ٌ���cd���=��  �Hp �7�~���f3nno���Ⱦ����. �gJp ��=]?��M�×�M�/nn��Ǐ�/ ��;  �� ?Ƈ	������j��0���a�V�  �\�;  _�l6�d��w�iz�����,����b�az}����  � �oj>���������]��l6"<��nz���n�~�b����� �+� 8���}"</�Ӹ����F	 ��� xv~-�o6�O�ϡl��q?n��>���݃M � x������7���
�_��v�V�q{w7���X�ߏ��r,�K��  �U�;  /���O_��nb�n�|껏  �[�  �J���� ������u[�����a��ߏ��j<�ߏ���X.������� ��� xS�V��y⭩y�i�4}���q}���K �w  �� ��n�v����q"~B~����l�j����էi�i���qb]P �9� �4���l6������k�ݴ�~�+�i��fl��ދ黈>}��~�  ��Dp ��.��V��O'柾��3O�����x��l��i��_[o6c����7=����z��vg��<��f3���z���� �k&� �3��K���/���_���  o��     ���     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �<�����O}&     <wyp_.���g    �sg�     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     ����O�urr�����nGGG�6���C� �����������C� �X,�y�\����������c��>     �3+e       �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �����|||���     �;c��+�     ϖ�2     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     y(�    IDAT�      �    @�>��~��4M��� ��_�V�}�K  /�l6�~������ ��*�����l6��� ���OOO��З   ���J     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �     �;     w     �     �      �    @@p    ���     �    ��c�ο�.���_{�<ABB�$ SA�T����Ӟ�o�u�����*CeRE�d
3	!@ $��CƝ����� ��~>�ޯ�\]������\���Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q@�       @P�       �        D�;        Q�=     ��������g��_�xQ�`0��&�˥��Ledd(55Un�[>�O�G^�W^�?G"��a?����A���+
Y�� ֤��+++K�x<�~_�|�G����G�`PCCC�������� &P��,^�X��@kii�ٳg�d/]�T�ƍ3����}��7F3����jݺu�ǈy�{X$<
�522�@ �P(����̄Q�W���ɓ��������8����	&���P�ƍSNN�233������L����!�H$���~���>����G�{��O�"�x�^���H&LP~~���������b}����~��~��߿���ݹsG===Q� �$
w x���rM�4��H`CCCֲ���URRb4�޽{F�7��r�����Iedd��-���>*�E��gQQQ�\e;b���QII����4a�)77W.��X���RVV����T\\���.������s��޽�;w��oP">x�^M�4I�������������IMMUQQ����~�������ڪ��������+��  3(�  `���Snn�rss������K�w��޽���NJ,<���Ҳe�l�rssUYY���JM�4I����Gz��ri���?~�f̘!������z��nܸa��v����4���hڴi*++{�f��,UUU������'��ب;w�(�X� �t�   �i����ɧ������ޮ��VݺuK�oߦ��#s���ĉm��(����/��3fh�������4��֪��V�pX�o�VCC�.]�ħwb�����ɓ5s�LUUUY-ٟ&''G,Ђ���u��9�?^�G �Ll�I   <EJJ�***=3�ƍ�z���^�J���233�t�R�c�9y�^UUU�^��ɓ���q���֤I�4i�$���jhhP}}�:::l����^�^x����KO��U,���Ӳe˴x�b]�rEǎc� �
w   Ľ��TUWW���Z###�v�.]��k׮q�=�,_�\iii���3JKK����5o޼��:���h��ٚ={����u��i544���>�Os�����󕕕e{����z5c���֪��QG�Ugg��  �Q�   ��|�G���t��9�;wN����G�aUUU�vg#����?*�ci/�����~�z-\�P�}���^�j{��USS�+V�}��s.�K555�>}�.\��C��g XD�  ������W^yE�-ҹs�t��q����dddh�ڵ������h�IY��\AA��y�ݾ}[�~��Z[[m��0���j�*�����(�ۭٳg���ZG�թS��� X@�  ����zUWW�9s���ٳ:r�m��(z��ו��a{�AUU�V�Z���lۣĔ��R��w�SSS����ϛ����vkѢEZ�h�<��q�����˗���Z{��e� 8��   I��񨮮N3g��ѣGu��i�B!�c�9���i�ԩ���(eeei�ʕ�>}��Qbڴi�T^^�o��VgϞU$�=R\��������V��k˖-:t�N�<��! p�;   �������ڻw�:::l��gTZZ��˗��4k�,�X�"��ǌVjj�V�^��S�jϞ=�=R\���Ժu��ԋ~������UVV�ݻw+�	 ���    �-EEEڲe�/^,���ko233��[o%ժ�x��z������_�lS�L���GM�4��(1��_Ի�K��3UUU������o{ Hx�T  ���v��d�m޼�]�q���護��k�������k֬Y�G�k���ڼy��͛g{���r��b�
���kr�\�ǉIyyy�����kv �	�   ����rmٲE%%%�G��p�\Z�v-�}�@yy�>���%!x<�Z�J�V��T��׫7�|S��Ϸ=J�KKK�{ｧ��ۣ @¢p   �Off�~�ߨ����(x�E�i�̙��������{��j�͛���~[^/�e{�i
���x<Z�~�jkkm� 	��   ��ϧ��zK�g϶=
���VK�,�=~Emm��|�M��4}�tmܸ1�_c�ۭu�֩����(q��kG� �G�   ����Қ5kTWWg{�HEE�^�uViĸ��Z�[��;���Ro��VR��.�K�W��f�s� 0#��T   F��r��^ӌ3l�Ieeez�wX���Ν����'el˴i���o$�Q˖-�HQ�v��~�zM�8��( �0�A   ��\.���모��=JR+,,ԦM����l����>}:�dƌZ�fMҼ�3f��K/�d{������M�6);;��( ��   <���ц�׿�U��ݶ�I:�����o~���Tۣ�)JJJ�nݺ�.|{{{��ӣ���G}}}

��
�D"����T��n���)##C������Q^^�rrr,�*�l������ѱc�l�bTqq�֮]k{�����Ugg�:;;���kddDCCC����4���(55UYYY*,,TQQ����,O�o���ڰa�>��c�A�� @\�p   ~Ejj�6nܨ���/�=N�(,,�o�ۘ*��K��X�B$Q[[�nݺ���v�������������ĉU\\�ɓ'k�ĉ1�&Ò%K��ޮ��ۣ�����7Z_-544�k׮���Y7n�xT��UNN����U]]���
��-..������W_Y� ��;   0
���Z�v�v��i{��0q�Dm޼��=ƹ�n���[��ʲ=�"��nܸ��W����)*��������Y���:t萲��TUU���M�4)�yc���������ǉ*�˥7�x���7n��ɓjiiQ8~��<x�.�JMMUUU��ϟ����(L�l�͛�[�n����� �(�  �Q���Uss�._�l{��VVV�M�6�F&���K֋�@ �.��������f����̙3:s�&L����:���Z�ퟞ����~;�V����i��Ɏ�F"]�|Y'N�PGG���@ ��/�ҥK�2e�-Z���cyO�z�j���y�
 ��; <�_|����cX�r��e��9W�\I�=�O388h{X���D���"����������x��������z�JIIQff������������Z��kV�Z�[�n�����(	���2�֓��Ə��_~�Z���?�S�Nixx��ݻwO_|�:�%K�h֬Y������b-[�L��mZ�l�����Ӿ}�t��m�2#�ȣOQTUUiժU�?�4==]k׮�֭[��DA� Op��}�#X����{��#Y@,���Oy<eddh���*,,|�0�����d����իWk۶m�GI8555Z�n��=��u�{�إ�Dt��E}��w1��W����K�>}Z+V��r+[�a5ȥK�t��+����x�n�:G��A:tH�N����gu��UݺuK˗/׬Y��3q�ԩ����] �(�  `U(Roo�z{{�Xۍ�cUUU�������m��0�͛��+W��,����:+�.<x�ݻw�֭[�g�Ugg�>��S͝;W������p��Z�f���׿Z-��W]]��������ӎ;����X��}��jhh�[o����tǲW�X�k׮)8�	 �����   �_�p7���?��Ϫ����}�+W��&v��n���kZ�je{�����ҥKϽr�����qQ�?�DT__����/�w���EEE���s<7Z���][��֦���/1S��XKK���׿���۱���L+��@��p  @�����W_}����������Dl��q��i�ܹ�ǈk>�O7nԋ/�h{���ŋ���D���jǎr,7������G�ƍ�g/Y������ꫯ:���7n���GL�)z����o������Ν�	&8� ���   q���W{���G}���.��h�<��egg�w����N�j{�A^^�^x�������ݫ��ޱLS����u�V]�x��ܔ����K�fFCEE�jkkɺy�m�S��z���!mݺUW�^u$��r��W_u$ �;   �N[[�>��C�>}�������~�&MҖ-[�ˌ�X�d�cW�Bھ}�.\��H�B����٣3g�8�;{�leee9��<\.��-[�HVkk��n�e�C�PH���c7�+++�=� ��;   �R0�����k�.�E������z��Ǜ��:m޼Y����G���竦�Ƒ�H$�={����ّ<'E"}��W��t�z�qu˽��J'N4����m߾]###Ƴ�-j���}��#y˖-�9 0J�   �k�.]�֭[5<<l%?==������j���<l6����ˎ�n?x�._��H��HD{��USS�c��g�VFF�cy���riɒ%�s���v�ء��A�Y������>s�A�EEE� �Q�p  @�kiiѧ�~j�t_�`�cEd<*((Ж-[4c�ۣ�eddh���d�;wN'N�p$˦p8�ݻw;�<
�ϧy��9��<���yH�t���9��رÑ?�^~�en��(�S   ��۷���+;�����~�'�3g���?�C�G�sx��dBww�8`<'Vk���
��͘1#�S�˥ŋϹr�Ξ=k<�)������/��L�8Q����s  �Q�   a\�vM��﷒=k�,+��*55Uo���֬Y#��g{<�˥9s��	�Bڹsg\��~N�ɐ�����RG����ɓ���o4#X�s¤˗/;� ����� �xG�  ��r��]�t��ܩS���~d'TTT������m��((//W^^��'N��ݻ�sb�ŋ����HV,�vz���g|�����3�c�����(���Paa�� �w�   H8_~���~����G555�f��ϧU�Vi�����ɱ=�d����3�������ωU�HD���S04�U]]-��k<g��������ҹs�f���_(��q� �g�   H8###ڻw�����M��h^,)++���G͛7/�wDcl�^��N�j<�����z+�߿��^�4M�4�x�X�������w�Yy·�n߾�.ͨ��Qzz�� �g�   HH�n�ҙ3g�,++K�"--Mk֬������8kҤI�w�߿_�ϟ7�/N�8��-���r�c���b|��ݻw���d4#V>|���^oL�& �(�  ���9�@ �X���֔)S˳���V��_��9s�p�=A9�����>�o�Voo�#o>����ӧ+%%�h���Ǎ�Kz{{����Ī) �W�   HX��,���0n�8���{z��7���i{d�p6��"�8�c�����'�b�̙F�����r�ьXs��)�B!c������� �(�  ��N�>��-�X�9M���Z�|����?�����80,??�����/:��g<���н{��fx<���������7ϝ;�t�����UCC���� ��Q�   �;�:''G�����9��ri�������o-X�@���H
����=FBsb�Lcc��xt��E��r;y�̙FWR�B���E}}��󫫫c�� �5�   Hx����D"��M�8ѱ,�&O��-[�h�ڵ1�>fhhH�|��޽k{��f�����n߾m4#^]�~�x����g�Fmm��󛛛���o4#V�����DFFFR�Q���p  @�����s�cyEEE�e�R\\�����ڼysL�zzzz����M����GIx���׮]K�5���ե������v���|��/_6z~�3�	/�o� @<�p  @Rp�t),,t,+�


�q�F��Pyy��q~��ݻ�������nۣ$���L����hnn6z~<�D"�u�ьq��=4�����t��5�������'�*++�vS-��ym    8���ʪ���0a�^~�eM�>��>�g��ܬ�?�\###�GI
N|�����xF<���Puu�����Ҕ�����Ac�f�ԩF�onnV04��������flETzz����Y ?B�  ����ݭ��>eee���ɑ�덋����P�/VUUUL��pXG�ѱc��ß�L?����W}}}F3������g���Y+����TVVf4��������ʕ+F��PYYI� ?��~   �4L�hx��r_����4mڴ�,��駟��ѣ��+..6z���T�WN�iii�3���*�P(���c���뛦L�b�| �7�   H���s,+
w���E��ú�?�����k��޽k��D����)))�3���3"n߾�@ `4#^ܿ_===��/,,Tvv��� �P�   i8Y�gdd8��H"��N�:��?�X�����IJn��xy�������x^���3��$�&M2z��7��oL�.�K������xC�  ������XVzz�cY������Ot���B!��$���Ly<�����B����@�*�3335n�8�����7o=��2 �o<4   I���_�Hđ5*�p��/j������yyy�3L��H$###�z���nk�����P���L{{��������xx� D�  �$544���s����������K555�����������f$
�u��')--5z~GG��Oě��{3855UEEEjkk3r> �V�    �:�c�Ȋ'W�\џ��g�����k������a����r��n��PVVf�|J��3}���) /�)    Iũ[�&�@Ļ��mݺU;v������q�3��ݺ|��Z[[������M>����+�?�^�


�fP�?��ׅ� ~�O   H*N��p��P(��'O�ȑ#�{�ajhh���KKKSVV����������edd(''G������h~�S���ρ��(((0����>��=�r�\�D"Fs  �Q�   �8U;�/Z[[�o�>uvv��`hhHCCCO���\.eff>*ೳ��������p�����pj�֏=���W���F3�՝;w�>8��p<@��p  @Rq�a������࠾��]�x�[�	.����O}}}�{���9>�1:�Z�=����x644�������(,,�p�/��R    IDAT�(�  �T�*ܓ�o(R}}��9�@ `{��::N�6n�������m��x���e�p�0a���(�  �T�z�i2�pojj���u��}ۣ q��(���<x`4���n���vuu=?ޙ��l� (�  �4\.�����J�����u��Mۣ q-##C���F3�~��6���1�)#n�?���}	F��x@�  �������J�dZ���۫Ç��i�����؃-�q|ܸq�3(ܟ�tល�+�כԟ� 
w   $���\ǲ�^�`�������{�9s�r��)S�ϰQL�.��������ga���r�4n�8ݻw�h �2
w   $���ǲzzz�rZ Љ't��)�H(�GӦM3����;��]__�FFF�~ڋ�@��p  @�pj�l(R__�#YNѹs�t��1�HH�<k�����3~�t��:�_�D���c��N��XF�  ��QRR�HNoo��#4ippP�������h���5�����|
��=6twwS��A�   H
n�['Nt$+Q�������ɓ:��FFFl�$���M�>�xέ[��g����1��+���_''�� ���   I���P)))�d��-ˎ��8qB	uS�us�̑�k���7n�����L��n����˄��~��;�� �E�   H
N<�𡶶6ǲ�%���YgϞUKK��q����x4g��9�H�����l��c�p��ʒ��R$1� ���   I���Ʊ���vǲ�WWW�Ξ=��/jhh��8@Ҫ��q���w����qL��"�Ϙ%�_�׫��t� ��;   ^aa��������w$�yuvv���m�$=�ǣŋ;�u��eGr~.++������
�BF3�o�deeQ�HZf�   1`�ܹ�e���������ĆY�f9�`8֥K���<��='
w'>� ���   	-++K3g�t,/��� ����jѢE�d���X+�M�p��&'^�5##��� �(�  ��^|�Ey��mRlnnv,@�{饗�|��EGr�t����sb�=�;�dF�  �������:�߯���� ķ��<-\�Б�@ ���&G��tK�>6�?���n�| �e�   HX+W�TJJ�cyW�^u,@�[�r�c���t钂��#Y����f�|Vʌ7��
w   $��S�jڴi�f^�r��< �k���2e�#Y�pX'O�t$�q\.���==?ј~��� �Q�   �deei͚5�f��������L �)##C�V�r,���I~�߱��KII��m�~6z~�1z>�;�dF�  ����x���o@��]�tI�H��L �i͚5���t$+���ѣ�d=������X�~�RSS�� ���   	e�ʕ*--u43�����L �i�̙���jhhн{��{'n;�RflL�^N>? b�;   Ɗ+4g��s�������x.�������+W:��u�������J
w Ɍ�   	aŊ�?���ӧO[�?�^�6n��認3gΨ��۱�'�p�=�_/��g|o? �*��   ����z�v�Z͘1�J~GG�n޼i%@�X�v�
���Ç�{��|��J��1]��\.�|>�. ��;   �����a�X���￷� >���9���C�444�h��|>��B!�A��ƉO���P�HJ�   �;�Gs��Ւ%K]��s���jll�� �UTTh���f�����ٳ�f>��u2cgz����'  ��   q���B�����[�}��w�D"�� �������o���8�
���_���&Ӆ;���Ή׌� ��;   b���VUU����4i�$��H�������b{ 1*++K���#��cǎ������_��J�����o4@,�p  @�����̙35g������p8���@���|ڴi��߷���t��1G3G��j�p8l��D��k�w Ɋ�   1���@UUU����ĉ�r�l��'O�TWW��1 � �ǣ6������@ ��;w�d����b��X�5�:'^3n�HV�   �������H���*..VIIIL�d���N>|�� b���ֺu�TYY�x��_~����sG�t�J�>v�p s(�  `���Vzz���Ҕ���q������ܸ�
��k�.�Aۣ �1.�Kk֬QMM����ϟWCC�㹣e��J�cG� �P�  8���\k֬�=�ss�ݏ��|�G?X���*55U�?,д#G������ bЊ+4k�,�s�����~�s��t�J�>v�H�xF<�� �D�  �	&h	����������� �^y���⋎玌����?��Ȉ��c����w 0��~   �����Վ;(u ���/���_~���H$��{��ŧn��{xh* �C�   <��Ȉv�ء��>ۣ �1.�+��b%����1���Ǹ�{�x�L� VQ�   O��i{{��Q Ę�jٲeV�u��1+�ς� `;�  �'8r�H�� ��%K�h���V��ܹ�ݻw;���h�{�q��;�$+
w   �1Ν;��G��@�Y�t�-Zd%���ںu������ge�p��7b��7�$+
w   �gΞ=�}��Q� x��ri���?���@ �m۶����J��0���]�c��k�' $+
w   �GN�8��R�x��vk͚5�5k���`0��۷����J��2����%cG� �P�   ��8p�����m� �x<�_�^���V�C�������͛V��=�8��7�$+
w   $���^�ڵK�nݲ=
�����a�UVVZ���ڽ{������G�{��; �C�  ��v��U�ݻW����GC��Ҵi�&���ZɏD"ڷo���G;�c�oRp�@��p  @R��_�K�.�@�����{ｧ	&X��o�ѹs��G����p;'^3n�HV�   H*�pX.\���544d{ 1f���z�����km�Ç��ɓ���=�8� n�HV�   HW�^շ�~���.ۣ �A%%%ڴi���ӭ�p��	9r�Z�	�`����c�w 0��   	-��ʕ+:~���ܹc{ 1���Jo���|>���;����Z�)�wv������; �*
w   $�@ ��/�ԩS�������̙�U�VY�)}��!=z�Z�I###F����9���@��p  @D"�u�Ο?�+W�p���Z�x��,Ybu������Vg0��2��� `�;   �Z8Vkk���Ԥ��~�#��Gk֬�/�`m�H$���������N0]�z�Tc�����a� ��S	   q����ƍjiiQKK���� đ��TmذA�f�D"���/u��9k38�tធ�b��D�D��w Ɋ�   1mxxX���jkkS[[�n߾���>�c�S���z��w���om�p8�={��ҥK�fp���6t��x��� ��;   bB ���������ݭ��Nutt���+��@(..�;Ｃ��Lk3�B!�ڵK����fp��А��}>��n���ќDB� �P�  ����!�B!ippPCCCRoo������۫��>=x�@�����O��u��Y�=22��?�\����f���w��%���z�10]��A� ��(�  v��e�8q��Q�)��ÊD"
��mS,X�W_}U.���CCCڶm�Z[[��`�ExJJ
���.��Z Hf�   �ݻwm� 	��vkŊ����:G__�>��3uttX��'�W������}pp��� �(�    	'==]6lФI�����եO>�D���V�ɩ�=�oP��� ���    �Pƍ�M�6i���V�hoo�֭[��N�v�p���4��s�@2�p    $�ɓ'���Vjj��9nܸ�;v`h<�
F�&�cc��;�;�dF�    H/����/_.��mu�.�/�P8�:G,0Z��~�%ޘ~�X) �Q�    �Z�<U�N�:����Z�H��(1���_�ƍ3v~ff���QVV���� �Q�    �VZZ�6lؠ��r�sD"8p@�O��:G�2��>##���������- ��(�    qi���ڴi�ћӣ�g�544X�#����=����x�?4������ �(�    q���L7nTzz��9����}�vݺu����t������Ȑ��2����g�| �e�    ��2{�l�Z�J���~�_�}�������zzz�����s��;�dF�    �n�[���.\h{���i۶m�%�7�)�G��k4<<l4 b�;     ��|>��曪���=��{�n�Aۣ��7�����v����$Ӆ;�d $;
w    @L����;Ｃ��"ۣ�ԩS����Dl�W����D��w�\��Ƞ�Ӆ;�d $;
w    @�*))�ƍ��	�Bڷo�Ο?ou�x
���ק��lc�C� fQ�    bRuu�֭['���@@;v�PKK��9���7Z���婣�����"//������7z> �:��     ��y��魷޲^������?�l��E��"9Q�7������F��X�w    @LY�p��-[f{utth�֭�Ȉ�E��"9x<������;�dG�    �	n�[k֬ѬY�l����&�ܹS�`��(	��ݾ��\���D"��~c�@<�p    X��z�n�:UWW�E�N���_�H$b{��b��3���3�=x��7� $=
w    �Uiiiڴi�JKK��
���W_�ܹsV�HT~�_�`��^���L�|>���9?�� �㡩     k�������[/ۇ����g�Q�����e�|���-�_a�����4z> �
w    ��������	&X����룏>RKK��9���{���O��t�_��w�= �+e     �+,,�o~����[��֭[ڱc��Α,:::�����o��xg��-�o� @<�p    8*V��˗/k�޽<��A����b��ǳ��\edd;dd��  
w    ��&N��͛7+--���HD�ұcǬ͐�:::�D�r���?q�D#�&�oFtvv*� �x�w    �#�������`P�v�l�dhh��-茌���;?��.��� ?�p    WZZ�����V����}��Ǻ|��� ���=��2�g�u�s��� ^P�    �*++ӻﾫ��Tk3��~}��Gjoo�6~`�pg��/y<�hmm5z> �v�    �yX����X����M۶m������o����ϗ��3v~��߿o�| �'�     #JJJ���ڳg������S]]]2�^���Hn��x�HII���oݺe�| �'��    D]~~�6m�d�l?u�v��I�c"��n޼i���������ɓ��O� �F�    ����l���JOO�����W_����D"Vf�ӵ��=���������v����h����(�    Q����͛7+77�J���o߮��z+�Ӆ���񤤤���������e�| �7�    ���z�z�w���o%hhH�~�������c��߿���c痔�(33���񤪪������|� ~��    ��<�6nܨ��R+�<�G}�۷o[��ؙ���r�4u�Tc�ǓiӦ=�ڵkF��xC�    x..�K����*++��wuu飏>b�E�ijj2z���Ӎ�
���g������  �P�    ��5c�+�����������^+�xv7o�T 0v~EEEү��9s���oݺ���� o(�    �l�ԩz�W�d_�~]���?488h%�'�ƍ��w�����������իF��xD�    x&���Z�~�\.���ڶm�k��2/�����cYUU�222�����h�| �W�    �1��|ڰa�RSS�nllԮ]�
��Ft]�zU�����/((Pyy���cً/�h����f� �xD�    �իW+??��܆��ܹS�p��lD��Ȉ�$���7z~,�8q�JKK�f\�t��� �(�    c2k�,�c|�K�.i׮]��	�tq;e�͈5/�����t��u� �(�    �6n�8�\���܆��ٳ��=���������.�KK�.5v~�)--UUU�ь˗/��	 ���    0*n�[�ׯ���s4�ƍڽ{7e{�
�úp�ь��*���͈.�K����ьH$���z� �(�    ��h�";���ޮ�۷s�6����Ce͚5�x<F3l�5k����׮]�����f @<�p    ����B�{������>��Ȉ��p^oo�����fL�0!�������˗�9u�� �g�    ��r�\Z�z��n�~�ڶm�˄]N�)Y�d���6��n���JMM5���٩�7o� �xG�    x���:G�_��a}������t,�ݼyS���3���x��o*##�h�Ӗ.]�ɓ'�9y�"��� �g�    �'����+���h�w�}��ׯ;�	�"���;f<'''Go������0iڴiZ�`���߯�/��x��     �X�l�RRR�knn։'�ClillTww�񜊊
-[��x�i���z�7�r��g>|���m P�    ���D��������jϞ=��HbN�r��hѢE�d�����w�}���vI����� @"�p    �����k�����Y釽�;w��!���˗�߿t�R���9�M���z�������HޡC��� �D�    ��iӦ���ر��'O���ձ<Įp8�o��Ʊ��^{M�f�r,�y���k������s$���U����d@"�p    ������ŋ˻��>�Xb����{p����ڵk�l�2�>���������^&Lp$/k����y�1�p    �DMM�c�^$�޽{�C�8x�ckL\.�.\�������:�9V���ڲe�Ə�Xf}}�:::��D��     �p�\�?H�w�q4?hooק�~j{�'�w�N�8��:�Y[[���<}������q,�i\.��Ν�+V���8�����'O �P�    �2e�


�s�\JKKs,����b{�_u��M�6��[�����ӟ���G��ĉV�����_]�g�߿_�@��\ �w��    <�`��# ��A�۷���>�O˖-�����z��x<�7o����?Y)�ϟ?σR�q�     I*,,ԤI�l���͛7u��)͟?�����R�������t��Q���=�f͚��^zI���F�����k���V� P�    $Is�̱=�X�~��JKKU\\�x�������5m�4]�~].\PsssT�������͙3G999Q;w���v�ڥ��k3 @��p    ��󩶶���c�B!�ܹS|��RSS���r�4e�M�2E��úv횚��t�����i���ӄ	TVV���jM�8�����7ߨ���� �(�    ����Vd�����{�nmܸQ.���,)))���QMM�$)�޽{����������B��RRR������4edd���P�ƍ��[�ջp�N�:e{ �{�    �G�!ˮ^��o��V�����Q~"55Ueee*++�=�3ikkӾ}�l� 	!��N    8.55U���� F����:w��1������ۣ�� ��;    $�iӦ�����}�������q���W���?���o{ H�    ��N�j{`L��v�ޭ�ׯ�%n�������zzzl� 	��    �\ii���1�Bھ}����m�w��'������( �p(�    ����(33���3	�ڱc�eƠ��G���u��=ۣ @B�p   �$VRRb{ไB!�ܹS��=J��������wuuu� ���      {&N�h{�E"9rD���Z�z5~����رC�@��( ��(�    �����]��    IDAT����ϫ��Co������l�"��N�>��*
� +e     �egg����w���?Tcc��Q�����'�|�P��C��    I,''��@���_�Ruu�V�\��njjҾ}����o{ H*�    ��<�222l���ب�7oj�ҥ�5k�������������u��5ۣ @R�p   �$��z�r�l�588�/��RgΜ����UQQa{$#FFFt��	}���
�����E�    I*n�utt���������K/i�ԩ�G����a�?^ǏW__��q  �Q�   @��pG2jmmUkk�JJJ4o�<UWW����k����t���>}Z�@��8 ��C� x,��o<cpp�x�����׸�����&D"~�q����迳�p��ٱĉ�{�M�~���Mmmm��o4s�L��֪����XO��ܬ.�ƍI�}
 �Iԗ�M�<�mxx�8��     �TPP�iӦiʔ)*..��g���E7n�Е+W444d{$ �SP�     �Lzz���?{w��ƶjtV�Vn�	� 7����>@��ɶe�bW������F�"��${o��6E����������������;�ꙇ������������_���?��$;��   ~�(�����������/�?~��������c�\�|>��i�6��u�V�xxx��j��*����������f�9���S��   �7���?��3������,�b6��l6�����eUUE۶q8������cpf�;   �u]��Ύu����      �@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H@p    �w     H yp��C��	     ��'܋|N     �hV�     @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @e�O8���'�ɼ�o~�g?����}     ���h�6}p��9Uo����1���     ^��h�&ڶ}|����M:yp?�<Ͽy�3O���7{|�4�9F    ���q]׏��o޿�U��ʲ,�,����(��ߟ����D8    0,ǀ���)g2���1�������    ���4M����s��Q�_���/!���4��     ��1�?}��f+�?C�e��i����ӕ4O��    �N۶QU�cX���b[���J�_EL&���g�o���    ��k�&��z|;}��l�{BO#����.�    |����}�������*���    �E۶�q�����3{����6Mu]��    � UU��.���U��y)��GY�EY�Q�e�f��S�u];�    \��i�~�M��/��KX�~    ��1�o�ۨ���qz!�_��~��Z|    .F]ױ�nc��F]�}��;��JO�O��ǵ3�;    pnUU�v���n7�OSܯL�e����w    ��d���==��4M�    of'��	��t�{�uQ��c|    x���O�����ǹ:�� eY��$&���3    �o�u��&6��C�o ���}����w     "��f��v��l�fODp��O���G    ��i���G��E��S���    ���v�xxxp�		�#�eYL�ӘN�Q�uTU�-    ��ژ�ju]�=��	�DDDY�Q�e4M���    \��mc�^�z�v���w�q\7�u]TUe�;    \���c�^�f��F��;?�eY�f��L&�{�   ��t8b�Z�n��{�Q���<�c6��`    .��p�����n�}�B�<��է'ޅw    ��~�w^Dx   ���Mp�U��w��   �i�u���v�_8��7yz�jUUQ�u�#   �`�m�^�m���;I�y��<ڶ��~M��=    \���b�^���C�m��8<��NRy��b���ib��y�    ^h������C�WHp�$������8QU��    �QUU��ݹ/�	��d2��,]�
    ?Ѷm����f��{�Hp����e����)    ���vwww��@�MQ�\.O�[3   �X����������w�n:��d2�f   ��i�6V�U���G�wz�t��n�s�   ����vqwwM��=
'"�ӫ�(���&�����    �KQ�Cp�"8�   �9�>.�;��KU   �Z9�>N�;�۽(����N�   puv�]|��%ڶ�{�Lp�"�e����{    �������>��uߣ�����eY���*���{    �������֪�ܹx����BU߆   ���n�����ܹy��r���ng�    �����Kl�۾G�B�\��|��!��}ߣ    0b��!noo��;Wg2�DQ��n}�    gg�?��= ��q�LQ}�   ����������9���ʲ,��yTU��g    N�m۸����_ܹjY��l6�<�=�   p��!>�M��=
Npg&��cto۶�q    ��y	;���(b>�G�{X   �v��ʾv^D�dP�<��b�2U    ����.V�U�cpew'˲X,Q�6&   �2]���ϟc�^�=
WHpg���yL&���    �J�m�>}��n��(\)G���lY�EUU}�   �k�&>}�u]�=
WLpg��i�y���    ���p�O�>E۶}��R�Q(�2f�Y�c    pa�vR���,c�X�=    Bl'5��Q)�Bt   @l�$wF�(����}�   @O���?��Sl'9��Q*�Rt   ����ӧO�u]ߣ0@�;�%�   ���Ω	�   0u]��ϟ�vNJpg�ʲ��l��    �H�4.H�,w���d���1    H�m����S4M��(����0�Nc2��=    �t]�>}���������leY�=    o�u]|��9�Cߣ0"�;|g>�GQ}�   �|��%��}�c02�;��|>�<��   p�V�Ul�۾�`�E��,�b>�G�e}�   ��v�X�V}��H	��y��l6�{    ���븽��{FLp�_(�2��i�c    �m���ϟ�뺾Ga�w���teY�=    ?�u]���F]�}���	�����%�    ���>��}�c���q�D   �˲��b�^�=D����U   ���4M|���1���/0�L�s   ����Ѷm�c�#�^h>���   г�jUU�=|C5�W��f�eY�c    �RUU�Z���Bp�W(�"&�I�c    �N۶q{{���C�;��d2�Z   �����i��ǀRᕲ,��|��    ����c���=���o���2    g�u]|���1��wx#�   �����U2\<��Z   �t����z���[�;$P��2    '`��Dp�D�ө�2    ������1�YwH$˲�N�}�   0m����C�c��	�PY��羬    R�����m��M���r   H����l6}�/"�CbeYFQ}�   p�����^Lp���f}�    p�v�]����ǀ���<��,�   �*����=���'2�N#˲��    �*��6��{x�N�)w   ��{xx�{x5�Nh2��=   ����vq8�^Mp�r�   ��V�U�#���pb���    .�~�w���'�É�yEQ�=   �Es��!���r   ��������ǀ7�����<��   �#���� 	�d2��=   ��i�6v�]�c@�;�IY��eY�c    \��f]��=$!�ÙdYeY�=   �E�l6}� ��pF��    ��~���������<��(�   �"�,����̬�   ���e���g6��]�
   �^�4}� �	�pf���.w   ��	���ጲ,��,c�X�=
   @o����mc>��=
$%��M&�Ȳ,f���2   �hu]��08�;��q�LQ1�N{�   ����ǃ�0�;�IQ������-S   �O�i$��g��E��1   ƨ�o�{Y�.Oe0w8�,����<��	   0:m����Ld(w8���k��   ���l��*^�V�pbY��4��   �k?Y,}�o&�É}�J�)'�  �1������|�;W�#N�W��#��q�U�   �_�,��r��	�pBeYF�e���r   Ƣ�_���b�ۖ�Lp�zΎv'�  �1����.w���'2�L�����   ���b��|>wʝ�%�É<�t{�׵3.   ��W�۟���)w���'0��^�JlY�'�   �,�J��X�e/�Up   ��+e"������N�!�Cb�]%�=�   ��=�����f3̈́�#�CBEQ���x    ��S�\�z������   `��{a��ʲ|uo�>�HY���y���   �`�t��S��2�,K8���	dY���M����    UE,�˾ǀgQ� ��l��WZ�p   ���b�<���o�ڋR��;   0ToY)s���;�e�x
�A�U2GN�   C�"�E��"�4p:�;��l6Kv2]p   �(El?Z.�
Mp�WJ�J���   ���="����I?�$��+�Z%sd   ��e���1��wx��b���S�   �y��e�����/4�L�,��7u�   ��W���^O��xD��y���$��	w   ����<޽{����^`>��,��   ���yL��X,'���R�;<�l6��(N�k��   �Мj���r�<��_x���,˘N�}�   �w�,�ϝ��Q�Q�پ5�	w   ��+�"޿�� �ï�y���l�ީ��
   ����;&��KT���0�����H�;   04�����|~�Ó�=�~b>����T    �z��]L&���`�w���tz�'f��   ���Ⴣ��Bp��e���쿮�   �9W�<�5?|��˯͸	��DQ1��{y2�   �)�">~�(�sV�;�C��\.{{�   �*��Iw�Jp��gl��   Q߱{2�Ļw�z�����,�b�X����4M��>   �P�f3ѝ���cl����w   `��>�x4��{�p���_�'��^EߣD��   pj��Rt�wF��b{DD۶}�    p�r�=Bt�wF�c{��   �p]Rp��9��ѹ���;   0\��#�F������``ʾ�s�����R��u]�u��    'q��=���̈��z��$���(�y���"c{�u2    }�I�2�#$��y,�ˋ���t;   0h��e"�F�w���=pُtx��(b�\^�-��G    8�K�3��<>~�x�sr�w�,�X,W�$)�   �o2��Ǐ/�D>��#�A�L&W�#��   ��Z"vY�����(���Q�B��(��N�1����ٺ�si*   �)�"���(˲�Q�2�;�2��c6��=ƋX'   ���l"8ʲ,>~����Q�"�;��eY,�˘L&}��bUU�=   ��][p��:�����Q��;W�(�X.�W�WKp   � ˲������b>|��8��|��?�e���j��#w   `<�9XO����?���'�q���ћ�f�X,������躮�1    ��MF��2U{����~�3J�}�Cxbs�   �k>8yt��X,��$�sU�������|��~��{   ��Bt�������?^��}��h�jL��X.��yR�.�C�c    �Ր�d2�b�o���`�y��2f�Yߣ$e;   0FC
�_?>|�����G��} �R�e�����jj���=   ��eYY�� �b���d��*���{z2����,�b>��b�dl���   ���r?*�2����mj������E��2&�Iߣ��n���m�   �C�_���>>|�0��'?�o���eY�f�X.��2r�   ��Z�!�N����i���Ý�PE��������n��    ����O�O��X��6���N��,��t���Q�f��{r   F�(��4��l��$���'�ӛ�,c6���T��v��{   �������Q��N������w��Rԟi��:   �(�"��{����f1�Nc���f��{�9�����_��3��v4��   ��XQ�e�\.c6����C��G"���ۥ�?�UK   �ʲ,�<�z��(��Ǐ��ﭙ�������UU5�o�   ��1��㚙�zm��9�,�b2��z}����u�#    \�<�Guy��dY�޽��b��&��}�#�
�;ɕe��\h�i�N   ��/O���(����1��c�^�s�2�;ɔe��4���{��cw;   �ύ�޿�L&���~���fM��=� ��fy��l6���p���m��   ���(D�8�w��v��lF�z��)�����<�   ~�(�h�VG��,�b�X�l6��v��ΟӅRJy�<�c:��d2�{���u���    ϔ�S�y����b���n��Vx�0�;�&���f���m�   �*�ϓ�y,�˘�������-����   �jdYf���Gp秊���deYF�e}�su�n   x9�����N����_�e��y��m�n   x%��u��}�XDUU��l�9���ʣ�d��4�<�{���^�=�   �RQѶ��(��eY�f���fQUUl��8}�5
���eY�ڭ�I�i�X��}�   pՊ�������M�ӘN�Q�ul�����}�4h��HE���ژX�V^}   x�<�#�2�%��,����qssc��	��#�eY�eim�	��n�}�   0N��w��\.�p8�n�s�=!�}�<��t�ɤ�Q�����    #�����I��L&1�L���&��}l�[�o$������n�����    ����N��X,b�X�~���~�s���> Y�EQ1�L�f?��m�n   8�c�j���QFa6��l6������p�{������ȞeY������WZ   N�x����eY������4�c|��ǯ	�W�(�(�2&���޳�n�T   �+�2��{P�7�W�8��W�����1���~��   8�,�"�s'�{v�h5"�p8DUUQU����/��Iĺ�˵Z�<�    ���2���onn��TUu]�Z�    IDAT�=Zo�s��,K���UU�ͦ�1    F�,K�x^��kg�����b�ߏ.���*�ڹ|]����]�c    ��������(�X,�X,��oV�}ﻺۃ<�#�S�����nt��   \��(�����!Ȳ,��iL�ӈ�h�&��c��z �����O�����m6��n�}�   0j��>�`;t�N:�ϣ뺨��1��u}����	�y���9~�0�u���}�   0z�C��\�,�/^=:��������FY�}�"�(
+b�뺸����/r   ��:v9�e�㸆����o"�����_��u�������+�    �,�8I�1�����54O�.)��?q|u�i\ϲ�����l6��l�   �(�r�������>�7MM���x}p?�z:��㏅u�����    ,˲Ǔ�Ϗ"|DD۶��i���D���S�O�����gڶ��   �
�^�z�ul¿
�Ǐ�����y��彠N*]���ϟ=I   \��(��:���K?�G���4·m���:~�#���	�c����ՅtN���η!   \��>wѝ�*�"�����s���G���}6�����?O������:���������1    x��>wk�9��
��%�EQ��3\��n�ժ�1    x��҇����TU���}�   �eYe��FmFFp�8b;   ���y.�sV�;�כ�ooo]�   00y���LHEpg�ڶ�O�>E�4}�   �	E�;g!�3j]׉�    #�;� �3Z]���ϟ���G   ����9)��Q:�l����Q    8��("�eQN�#��9������(    ��,Kѝ��bTڶ�?��Sl   9ѝS��b4ڶ�O�>��   @D|��v�����(��    ���TI��{ 8��i�ӧO�4Mߣ    p����,���͜pg��C���b;    ���y���ɼ���`�v����S�m��(    \ѝ����f_�|����   �+��yL&�Ȳ��Q�B�;��Z����Nl   �U�,��,Ew^Lpg0���/_����Cߣ    p�Dw^�B"�m����s��G   ` �,��dM�D�4}��ܹzUUŗ/_<�   pEQD�eQ�uߣp�w��f�������    `����ڰ���\���b�Z�z��{    F�銙�m��$�suڶ���ۨ���Q    �,ˢ(��ѝ�ܹ*��>����k   �7Y�EY�Ѷm4M]��=Bp�*t]�����(    _��/S݉ܹM����)    �8O���ʀ��E�n�qww�B    .ZQ�e�3#'�s�ڶ��j�ͦ�Q    �Y�<�<ϣ�k�����ũ�*�|��[p    �J.T/����bT    ��i�qܹN�   0DN����N��j   `�v���������s�   �Q8�v���Q8���k�6V�Ul6��G   ����<&�I4M�� 	��z���je_    ��eY�e]�	�#�s��>V�U��G   ��p������I�m�����n�    .R��1�N]�: �;'�u]���X�מ$    ����~�;�m�۸����     /�t�L�4�B�2�;��������o
    �(����\x�2�;ov8���>���{    �cxo�&���{~Cp��꺎���   ��EEQ�X��	�X]ױ^�c���V    8����t�x�L�;�&�   �e8�x�/���o	�    p����"��S��!b���=
    �O�{۶��Dp�/��}������}�    ��1��mM��g&��h�����C�u��(    ��yy�G۶�o���>rM��f���f�    �޻�{<����#���c���v��{    �Ĳ,��(�9�n�Lz���t]��6�뵵1    0B��~��n�LZ����l6��n�j    D�_��8��v��@�m��2�p8�=    p�����.���_Ip��뢪��l6����    �"Y�E�e��]|9�} ����v��ξ%    �;��V�<��~������    8����{�4}�u��+r8b���n�����    ��w'��Ip�`]�=Fv'�   �K"����~a����~��.����    \<��+��g]�E]ױ�����}�    �jO�{D<��1.�{�4M�Ǔ�cx�    ��y�y��㧧߇v^p?��m�����.<    �������6��ɂ�	�u���1��     �ʲ,�,�����k���u]����~�    ��#�q�� +h�8�����9�    @z?
�������h�曰~8�i����    ��
��>"���O����>��m�ͩ��i�p8X    p%�������\�>�w]u]G۶�A��q]�N�    ����O���1Ŀ�_up?���?~ԏ    @�?��?U�7?~��F����=��m�8��=;�||;�Q?�w     H�G+j~�� �<�����W�_%�~7�P    �����|���4���pH�i    �=�\<     �K�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    @�;     $ �    ��o��$�����?3kc��)%uҘ|EJi@B"��R"��Ui0D6>ggg����N�&������>��*L�*7(�"��ׄ��$�0pk�w������"�������>�������>��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �e��/��/�������0k.���k"��z0������m=����׼�����״�̾|p�Gy���Υ�^z�%�\��[� f�c�=v��?���; [i= v��h�DD<��`���~����G��F��]�o[� f_��g��'[�`�F�WD��n���S���w�G@6'e      ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     ��N/">�z0�J)/����;�z���#�#���̬��Z�cD|�����ӧ*��_o��Y�#�N��_[��PZ��l8v.���+J)�"�u�� 3a#"���:��z�����?�v���Z��z0>�����{8~��Ο�x���d򆍍�K)���`&���RVj=���Sbuu�j�qeD\�z�휌�{"��~����chk<���ɓWo���?j��~J)�Eđݻw߻gϞӭ����#�זR����z�-}��z��������?�zl5����Ç_����w3�<��`�}��z{)�~����c�.g^'�Z���{��7��߫�����z��#!�\�R>G���?�w��I�=p��0��=:�ĉ�"b1".k��:F��N��_z�މ�c�~�����W�π�?��R�]1Z\\|�������J)o+�\�k��*��Z��`��c��l��;s���,�Z_�z�V)徍����~�J)��L�����ϖR����l�h�o#b\k}�`0x�����	�"�'[��z<"�����_�-	�F�WD���ƈ�k<8NF�=����`���c�+++/��k6���[�ΫJ)�ݻw��}v2�y$�y�u�� �՗j��&�ɭ�Z�10w؆VVV^��t��Z�F�sZ��F���N����������Z�a6�u�})"~��`˜�����?i=�����\[[{�p8|���&�;lc���٧N�zs)�Wk}I�=@�����kkk���n=��a�u�kK)ׇ;�0K��R����k=�������xcc�m	�L���Z�؉K���"3ଯp��W��<5�3-������="���<%�Zo���;������cع<����^��� O�Ɉ�'"n����j=���3f4�:"�E��#��x�����E�J�߿��8����J)o+�\�k���<PJ?~���p��z�q�#���/Z�~(_�����r[���j�1�]�0����_��v��Z���|�o�R~w}}}eii�����s����'N\O�N���{��p�>���`��c�9���U�L��"❝N�^�w���nw�q7�|�����FD�#���">��Z�3o=��Y��E��Z�b-"�>}�������n=���Ç������	�tp�r�C��w���k��~D�R�=�ӔR#�w�wϞ=�[kyy�;��oEĕqA�=��|��z���{���[���k<?�ԩSo��ň��z�0�"⃵���`���c`�m�y_��+��NG��R~{qq�c���V8|�������n�zn�=0����r�������;i=�;v삵��_��.F�?o�fY���N���Rʭ�^��[�Y"��v�С���^o��>���!�*��5�LVo��ƿk=·���v�o�'_'^�z̐����Z�x0�~�1p�l>��w�!ӧ#ⶵ��w��o��Hpb<���ɓW�R���K[�m쳵�csss���z�p��{��Y�������NF�=�n������l=Z�Hr8q	���?�wޯ��"����6�@)e|�����z�10-F��+"���xcD�5��ŗk��O&�[8��c`Z�F���Z����S�N�3��z�z��;�]��?�FD|��r������lee奝Ngo�uoD<���RF�ѵ�����'Z��iu�#�~D�L�=0��UJ�+"F�����;��|_����Eĵ��ߌ�g��S�x)��N�sxaa���c`;���>u�ԛK)�Z�KZ�iPJ�occ�`����RJm�����;�mD�k����;��������#�Rʵ���{��/�Z�X__?����Z����̝�Rʁ�xe�=��Ɉ������z�zlw	��'.w���~�١=�8'�������֥����{`��R>G�g����:q_D�>"�������>��t޻��>^ZZ�B�=0k<b�و��Zg0�I�1��'�O����זR�_�d����zd0|���	���_��v��Z�����&"�v:�;z�މ�c`֝�H膈���Hv��rg��P���\�1�wȀ�myy��;���#�MqQ�=�4�E��q����U�1��|��?277�я�k<��١�Zk�F��3��Z��sss���z���H�����R��J)�E��Z�s�Z��dr���z1/ܵkׯ�Z��K���98�������� OZ]]��Z�5��������}�@��G�Ο8q⪈X���j���ODĻ����7�h=���yg��f)�w���W���>�z���r�-?:�L�^JyGD\�z|N\�6&�[f�����}��{`S����ZǾ��ˡC�~��z]D������{`�g"��Z�{���� ?��pxѮ]���Z��GBL�������Ӈ���82��  
(IDAT����܁�byy�;��oE�#b��v��qOD����?�z�ԍ���<y���f�����TJ�/"��޽��={��n�xj<bJ|��z���{���[���8�>�������h��z;�Wj��*�������z�g������AD���v�ID�^)������Z�r����B�u!"���Z�aG��R�-���ػw�� ��4q���]�n��x�������Lz("���t���z'Z��������"|�%߷J)wM&��o���Z���GBl1��a��eh꬯p���z�_)徍�����δ��zYD\[k�͈xf�=l{������;������c����ѣ�'N��*"#��{��NF�=�n������l=�:�;05F��+"��p�sw*">Xk]�l=hoee�qM)�ڈx~�=l;�R�Ǐ�{8���u�P��Y�������/�Zo�L&�8p�k�� [Op�����K;���Z�ވxN�=L�Z룝N罥�[{��߷�L��x���d�Z�qy�=L����p)����?n=�N	q�<"޹�����p�D�1��#�Sk<?�ԩSo.��j�/i����鈸mmm�����ۭ� ӯ�ZF�ѯ�R�w�����R����k=�<�{���Z�؉Kع��L�cǎ]������^D����)��Gv��}�={N��lO���?Wk�&"���C3_��ޱ��~d�����lO	��dD���t�z��h=hKp���h������n�9��"�C�Ng������`v�r�-?:�L�^JyGD\�z�G)��q�}v ә;凜��N�Rʝ���㥥�/�L�ؖ���_��v?Qk�o��-��R�//..>�z0����E����Fį���W�~���̶��իk�����V���w�����N��L�N� O�7��Z�7[�`�=$�[m8>Qk������?[o f��ӧ?�z[���?�v��     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ��;     $�     ��     	w     H �    @�     �     �@p    ���|�c%��    IEND�B`�PK
     D"BY��Ed  d  /   images/5779bcfa-264f-4061-b24b-5c8b50561781.png�PNG

   IHDR   d   �   �K�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  �IDATx��]	�U�>3sY��a+e���-V�e��ڠ!l�Mi�V�m ���mZ������ԘVA,({�"# ��00�f��Y���w��g�ܷ�{��{Η�y����������X"
<(���+�.JJJD}}��u�l�>_Iuu�"##C��7o^��"2�����ׯO�����p��iii��u=WZzz�u��)Oaߚ5kģ�>�༰�0@�N��WTT�]VV�/m�t@o��T�����|����k׮�<�H�<WBT2����N���AB��\G?É���w*I�m�sr��u����/H6�8��?$YM�0v�^�:Ԟ4 ����Ba��d`pې�-~Ar�d	6���8��5�	� �x�$�d6@J�G��'���T�ak�{ؐ�8�X@�0����$�I[2f��
w�z�;���#	,�)j�]��ng�����K1����nY�쩻�[$�2!�6C�γpq^^���믅A�ˤm۶�z�n�1!�%��<
2
ŉ'�юāj���B�▟LHK�0gbNN�4�ޡ��6D�LH��d��/��N�p�e'P�kjjd�iӦ�1��d�sG���册$���۪U��~�y��cǎ��*�5�0PFr����<4�]{�v$ږ(�7j ���/�4��ɓ�!ה�3$�~�'9Jr����\��0!hAHWa���H�"A�%4CUU�Ԕ-Z� ;`���Ռ��尰�!*H��O��� ���H��'\�|�PYY)5E��
:}�O�֩�8N�"��HJ�NX�hQ��Z�J��

�r�9�ycȮ��l[�}���ҥ�N?h�H�,�H>,�n�|2v7�l�X�B�<M�ɫ$�#�+|�lC


Dqqq����+�A�c�Φ�	�Q˗/W����I�	����GXh/�������K�J��J�L�CcP��P�� �,�֑<��Hni(ĠݚB��`�t $[ؚB*�p����O2�dI�b�M�ea�Q���6�^�A
���I�N�s�M��\�A;�j�pB%���n#=�OI�O�3�FiC�Pw�x?�,Y"t�իWŐA�ĕ�Rt�����S9R�!555u�!2 i�ҥR�Ƅ�c�o��=ۖWT̻V^.����D}#ZA/�^2�����oRvfg��WTV.!�ٶ��v���O��W����9�F�Ja��{�M��F��B��N�&�?���;��$e���(�]?J�G�������$�1�!�`B�I�C+��s�Nu�oU�)�&�E�{�3����{γ�]���w�c�@J%|#n~�+;����KD�Laǽ��N�Ú���e˖59�T5��G�}^���@���R	���c�B�D����+���$��b���F�"'\�@Eg�i$�!�v��AHZ
ǈ|#�%�o��a��/���Ժ��j4`��F��(~��F�w�p�CSB���C�������-[�Q�00(�+6A39)�!� IE��E��� �`o�$C���� Ȩ$�(�t)�C���>G^Ĉ�A��<�f;)=�S������sQ�	�b\��Ã����E��+?�|'hM�aD]$LJ���:��)~{hA2!�LJ��̇q�w��(��P�!h
��ݩ�ZA��Yj3����0(�d��Q@
�%�0�Ȃ�Bq��H�R:�ĤiG��� �01�*1 ����⒒P?#]��=	a ��W���gb�F}p���j)�}���VAڀ*���T�S߇5/=]�Xl�	Q�={ �Ϥ�/�2<-��@WM" U��5LG"͆�P�8�Q�!�(h��5	�%�JN�h�PKs�|��&h�U��C�f0�hC�f0�h����7�r;���!�������慈A�{�ɉ�XM���4m�lć���`|�р�#b�6D3+K3B4�!D3B4�!D3B4�!D3B4�!D3B4�!D3X�f^^�`�=��VC�!����䜋�K�Ta>��!���!���!���!���!�A:�����q�鳺4�SX�յkW|"�aֹ�l�3!��H�`��`�I#$�D���#�\e�F�{�:A �g�\��C}�H�bb������̌��T2��/����bL���
�u���uR4��]�vrb|#�	�9]��0���g��y�\��sB��v��;w����K g
��@����J��>}�ܷa���YYYbΜ9r�&g&!���={�ŋ���o��vy�͛7�s�΅�Aw��YL�4I���O��3��抝;w���"����:44Y'�ܽ{7���u�yO�~���!��#F��/�o߾��c�W�l�X� �P�����r��I�2t����W�^�7ސ�rZ �O�>�iǱd��Y����ڵK\�tIt��ML�0A����oJ-��S�Lcƌ��$�;��ƍ�iegg�
��H
!�v� ���R�LPMl�g�۽��;d	e�Hh�ԩSŰa�ć~(��9�F�'N��9�*l2D���[f<V�F� ���L̞=[8P|�駢gϞb�ȑ�?�g<u��=z�8r��O�6�3`B���}��?�h��d"�vlef�?^���{��+W��{ѽp-�@5�Y�x�.ȩš}(8\����
�����v5B��j��b
�P�1�hO^�uq��	Y��u<�9t��ez��!�M�z�Ѩz1��k�IH�\2�=!<͟j���<y��`d>���_�����:���'���?~\����8�$u4lCp�Y4�^/�:�)�����'�HB�,u
�X Mýf̘!��M�6I�����rދ�L�SVkB��%%%�a璍�@�!��@��2�i0��u�V���5�L�6Ǔ��Ӛ�R,+��&T#�R�~
2x�ƍ҂RӀ鋪����z%��~�! 2U�W6?4���b�̙�۲e�@8�j�!�aA��o߾�l����:��d@{B�2�Ӵi�d�B3P��l�9sF��(�Gn;ЦA�p<+����h�fE��"�=N����ݱcG�6�{���ѿ�Y�<(��nI�N��ur�����S������Pr���X�M�~@�`o��U�p_n�a�Y��ܯ�o� _\?��G}$��d�o�tB�g��;��mgCȍ�m�B��(��֭��M-�8�������)�ek*��p>�6����@�����7�Y$n�]��zg��	�|6(@;A�QM��k9��h)w}<U`J'6'���2{�!���	���`5��'K�#�C�C~��Ư��:X�6켬:g��jު`"8r&5��Xn���52����\<�薟Q�u�4���7��
q�
vL�:;���f3��?��bY��V�0����ĸLy|f/�+h���@���G��q±R��Wm
�"u"/$l�$<�y��!��C�t|� ^<&�"d$k��f�F�
Ik�A��ƻz��������aM�͚��j��ZXA
��|�v7,!\�9�V�[��ѐ���c�7D^"�`��c��	/���@>��0mȈ���#��X�׃K�s`�7y��0	*�n�Dnp`�Z�31h�!삗��`���Xv�� C�7���;�\5��V������=m4#>�w#��IVY�gF�b���?����ɵQW�.��b�of���e�����B�-ev�:��0�\p��喳M0�ن�&���0qY���!���!���!���!���1��/c��Mp����N�)y��2���322Zu�ԩw��q���QȊ�������ܹs�4m�Veiiin��([�{�7�������:'����� ;]�e�b�������<���:��"qy��'dff�u�ر�����W/^�x�u�6[%���ѕ+W�-..����j�=G"�0m�� ����z�{Ǐ�u�V0���1��?���{����͚5���`.�tzU^�ծ]�*L*��U̟?�_Vy�_��矗cvS��,L�T`zVzh/��iw�y���hѢ0���i��8�6��o߾��iZ+V�@�W�}����7V�f0�hC�fH�Ե^��G���j��LL�9�R�VS/H��r�d��q1ƴ���� ӓG�;�/ ��EZ��Z�1!BN��"y��A�^q���WH����Ztǐ<�>q�u��U�-Q�l�'�K��w�GZ��im�FS����!gH�%y�d�c$â\��'y�4[�B"����W�^E�z)ɋ$�I~E2<JZ����E�3�@�LB���$+If���ddie��L�o5��x2�"��
dc�����!�E26�� p9����DH�
�Z"o-i��?)BZϓ�1�=cHߢ��DHk��LLi�CB��(�Q.+t�GS�����
M��x�'�J+�MWbMK�GS�ً�R�Y(|�I�1L?D3B4�!D3B4�!D3B4�!D3B4�!D3B4���A�{㮞�    IEND�B`�PK
     E"BY	��} } /   images/bbfae99c-8036-4c5e-89fd-a87441410720.png�PNG

   IHDR  �  �   ��ߊ   gAMA  ���a    cHRM  z&  ��  �   ��  u0  �`  :�  p��Q<   bKGD      �C�   	pHYs     ��   tIME�#Պ�  � IDATx���{�m[���Ƙs����8��GսU���袍�i�4��A�("�q�6'9�Dq��E�HEVd��HX�d���&�Н��g=��n�}����ךs��?Ɯs����{����f�J������k�5�x��p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8���p8��}�𵂪 ʳwQʄRZ����k��{�Lǁ�%O�h	*T�J�`011@��#�QD
*B)�@ FI�"4"L�Db4��L[�>T	
4AU0����11��*��J���N�L� ��m��l@�(`\m.@aW��7W�G�|������%���<�Ç?���p8��h��@K�J���s�H��K���EFi��_j��R�kh�,A	P@	`   �jQb���!f(PA�U{�B8��W? � �FE}E��z�T�0b��P�t�>��1�yPr�P)[��7���I�����>P�+��T�hT ��ۻL���J��ui� ��5%Nd?#��z�vH
U�w�[��}��rV)R�""�%' ��f�v�U!�bs�!lJ���x�/.��Σ�~�S�����G����7 xD������%b~�]  A�=��~l�,!	"bz���
�*�E �
$S�
t�Nb�Z�L�WaEM����DՀ�Ĭ
�h�AU���!7�(���?��˯���1(��a��%�۽�����]���$���}i8���U�5�ժ��T�[T�GE�C-�J��eC�����	d�VE�RM��F���dQ�liO~M�?'0�w^d^�b�Op�x<��L�$����3x� T"��q���/@%B���w���w��ڄ����k��3o������k�q����:Eӯӳ� e�n|�Z��	U�M"�7h�Yr��((W���� D��@U�����y��䟽��� �6� ���X��D%"H�T�(�R��0+���	|KLO�x��8L����m.��>��m.@aa�]�%����P��/  �Sm/�J��eM�7h.�SD��J�$_+t�RM��
 ن^X�f��@�aJ��QS�t��k��纽o>c8y�l�BqĻx<������{MH��sF����J�v�������U�v�+��K�������]^\��^��������ԟ��|�^�/�-�p����; t�0�>]=����_.���FD�[%���P�)	R
b�K)PUÀq� ̦���2���_�+t�;������2{��W�~N�D�DF���k��q( �fB8�g���90��2�d�����q��o}a�X	�@�>�G�ᗍ�VU����n�./��'�����/%�n���Z�K*%��Pɦ�T d�ά��H��Du�Z�9��yeӕ�����}N�]�v�W-�~��;?��c|���	s)(���QJA�fB�C`036�`6q��F��,��j�@�.�q�}�_o��v�y�~���g��W~Ƌ��Ǉ��q�`ڿ�_�o~��-������<�Β�o�o��V�|����D2��\!���!F\]_#�(Q�W�Y7ƽ˧3]oqǕ�\`S���"ZM"�� J�jTM1+���y����M`��P���ϙ�gƟ��~�Ke�q�1^\!��1��,���;�������/b�]�����U��HI�Z2 ��"	���`^yۨ�j���l&��mH:��@��l�
^P]���u�{	@��9��s��{<��s�7��.���L@��i��%c��؍6���1b�<b�#��E�0�+l����U�_�������b|�_n���7^^���, "���~����g~�G_�2��W����O�����%�v��7�i��|8n��[���R@*��PJC��`�!9���E��^z�U쮯�(��RU����� p� )�z�5���5ki_2����&�5���5�Ye.1WEO�����9
�'����e~������3������1ݾ��}�������o����!����?��9�.��T��9���I�"')�
�慢�B{�g�Z{�^IU��mt�Y�8��ieٮ����$��qԮ�0Q���.~a�9|*���ÌL���9�((#cF�P��BDĆFly����.�<`Ѐ�p��Kx��|}��[����/�~���T�O@)������W�������~�ǿ��y��/a�yʘ��b�]���o�Ͼ��2r�~��p��3,����4�P) ./v�$ bLsƓ�^z��x�ʫ��
� "���ӅA<�t����<���])U��kH��Wy��P��]��� �r��G��C�U�/J?�!�(��#���,o�M���#���#��p}�����u�П���|�G�|���������e��_�|+��*�Z��BHU��(t�ͧg}	yK���*3
�U](y%@hM߯��@���a�y��`��s����N_�8�@IAA���`F �!�b�
��1�6<"P t�J@���p�勏��W�`xTv���8?I<��ƿ�H���4��.��C   �7��+��4�i�p�x�xx<D
�:�ߖ�߭i��A��8o���� � �3��Md�H���#��9g�./����g�N	�^~��������Č@=Q�z�I��;:_���LV6�^�l��H���_׾6	�<vQ q�P��@���Y���q�� �o�D7x�c����@�P���/�*��A_�����폐����_�^�����Ayz�� � �J�h�V���c��S�w�Vν~I5!�)t�j�/%]š� 뤸��P���x=@B"��%Ct��@Q2��j�H1�Z��JI#2fd8!% `@�� 	!d��������F��:��?����R/�t�{C�o���6=~��v��o�~�qw����AU�RP��Bd�p�:s)�ó�?V4��9�ߍi���p��·m)�I��{H:@JB �%�'H�(iF>�Q�H4(�>�@cA�	�M7�i��;()D �%oz����q�9t�:W�dg�o�;��#����u��I�%�X�a���|����(�߮y�#!���@o}���8~vs���[_�N
��~$�}�y��޲,� �Q*��9�%��kXӀ2A҄��4�z�P���oYY����aJ�E�*��j_�*�cYXk�PN��l-(/4;��.�S*7����S�����	��IZ
� H�H�.� K-��"
5�d0�6؅+\�x�W.���xix	�0"`Ѡa��4���g���e��2���x��p����-!����n��K�u����9��3 �����͗���o�*2��O�\~_��o���O�i��N��y"�3Ho�Z 2!�#JN`"��9!��r�0�nn )!��8D��r��E@q���5~�۰���FFV3#R0Yc���Q�.DW��ޛĉ�~��P3	j��6��*s{ͪ���O�u�y�T�����UM�0(�X
�'a:��C�i�ݏ�{|����Ȓp������/	_W��/}�!l>���(�Z��-��D'@Dg�(D$��I�\��%�-h�Ӿ_|�U�v7Zy��1o��B������״}��;��"�ܴMȋ�iT�b B$�j�,�JBT�[J�A�X���B� �غ �H ��`@)B�6(��3o��4��4 �	�kL�c�O��g���8�0��s�Ͱ�~i������w1lw��t-����@��m�$�9���M<|囯5��۫W?6�~�j���K���U��n�O!�-�dYfhI�r��-E��	I,^.9!oq�y
��0n�u����3�4�c��ͣ�-bܘ�#��a�K�J��J�S���$�U�ng9��޳�R_T�9�h�EƂ�@�����OՒ�J�I9D����)㯕0��D�ߺ�<�����~������������O|�ʬ����O�ւ�Z��!�㿡e�(�)G�r�j2[���T�<s��qن�R�T;�Ψ*t���F��9��z�Z&'銢jT�4*���-���9��ւ�Y�]D@PD
�H%�&����Q�VC��H*�b�#Ka�]"�Lϰ��pF��~ʀ(
�y�&��M��7s���Y���t��1�� ~!����g_�t�3�C ¸�Ї��43�3���/�ٳ=��
WWeh���u0����#��̀�rP@b-}�j%A���BH�L@mX����D���Iָ���Z�X�K���jZ����1�}��p�b��`@IJ�A��AT0� Ί�2f�vD���q����Q��0E�t�c���
����v���}����;�y�%��j`���A����o��I_�"��>z=ݾ��*�E�'E��Z�5D8���h�C��	�@��|DIGS� H.ȹ@0�	ДQ�#�t � C���05���uw��"_? �&[T$K||�7�ӄ@������u�{��KoΏ9\����%/D��=����f_tN��;EJ�֛R7J_#�@uF)�e��{�O�����~����~�w~�w�����V���u��o��|���W�|��K�H���"G�L�2�lJ�%ͫn��1F��Ϊ
��w�yL��M����E)��z�ž6^O�:��׾�aU �Z"@�lB��;��,O�@����z!�$(J��ށ ���l���p0R�Ť���3bQ\L��-�����A� ��RB�v������5���������3S��8��"z�oso!�o�?�O?���q(1��%��f�tv"�w��T�Բk�a � J�s�a�q���	L#�iF�G�M3�:Z2r���<�������}��ʟ���G�q���D��2LE��FG�b�c`��B���L��	, )�M��`bb��Y��I ��H�tr��7�>½�
�����_R�U�Fji����P��
U"����V!�K��R]
E� n�b#��:�Ah�t�����p!P �����^������ 8>y��h
n�S� xh+�Q
�60C�~a�.�J�s�JB��g�o��}�f�g��]4b��� )�����/�9^
�Hy@�!��H�q���7��oW�߂r|]U^*%_�f�P�W�Vb�%��@�y�e>"�(ǣy���-e���'@b��%c:� D�4�e����!�@nn��gL9B9X)Z) ��oN��%�T��G�ÛR&��!��Xe�$��nғ�A+��.R�m�e���Ξ-�K��%�i3 c)lT�D@��H��)�''�o.����nz���O��#���a_+|���f-�a�0o����5_)�R�Ũ'�H-+SA˃T]�oQ�a���g�8M�X�jU�X�6ֹ-���s��2�kѩ
Z)�wR��G�؅["D�Ь(�0A� 6A�(g(B��g��#B�dU*`Q����)^C�
�hA��43��A�!��A�^�^"���{�BxF����D�%����ox� �q����ՌF��� r�0��N����N3�W��z���y `_��"����.
D>����d�"ø9��IidC�qP�AJ� �1�C��n�	1��R؍X�S�4A ��(TsE��*7�\5s���C��L꒮oZP�7�7T�/IAbJ]�i*UΩ�Y�(DETUE��Q��q��THJ	�E��,Y@9�EU���PJ�&*��"���T�\��-�˂�-Ƃq,�~�_�9�B�R����٫Z��*���l��r�^�3=��C�<�������`�hH�޽P�E�#��HyՇy��\i�;���9�ΐ־Y�'ת
J� �(%[-�<��#��M	�fS�R ()4%d�ӌ4O��0#猔R�P#�b�R��0����f�� sg8툩9�M�5[���Kύ& ���K�{}��$ԭ����ԍ�ƪ��ηváv�_=]��p�b� �d�I�oU%��w�VDE�n��2��ܼ�i\����zV��*�ӻ�'{�q�M���/i�sH�G(gh��V�V2���>���@��L�QSƴl�N�t^~��۷}JQ{]/1��Q�&�v���^N� ���M^[�f��FR�`l8��#v�E�2CHl�Q��I�d���I�zp�`��DDe	 &&��Tn��u�b@s���\KE2�L��  03�Ja$#��� V�P�C��8&���(4�(QS&��L���U���(I��+���� ����k����v
�<;��T�i�����a���2���(��r�BsR��H�L��HDL̡*_��i`Bd!��͆i�/]1^}i
�U�K��q�u�V�����û��|Խ�6L+MD$���Ｔ}L_՚����R/n�7o+%Y6qVe) e0���([�DDC9BDTPP�([P�P	[`���P���VG��"�%�HI��R��Ǵ���V�!T�T�c֜7�������Z�̌�{5Z�v<UHUI�����V��b��*K� RX�0����b^}�P�*��g��S�Ħ�i�q	e>�oQ��d�Ϥ-�Rl��������
���cJ8���%��ْ�b b4�:M{H� �S�-iM�@cS���YS���3=]<4e�L��&��7��D]Q�2<f-��w�n.�~��G5�,"�mb%S� ����Cx5���k���n��4r�x��O��Z����~��C\~��雟�m�������'PI֛Xg@��=��F"�j��V��w~" O��~M��S4����z�}�,���歯�f͆��ڇ�d��fc5/{TƆ��BϬPeX�2��Q�D��p���� +#h@�!����!?E. �ƂѕD���huRTC��� �"�z��`G�� ��o�����Z�&�Qz�w��y��CUf�<eL���O�xrTd,�X2B����$b�:
�xf�<�3{�D*}K1�ĀAB���0!h��̀a�������D!�����жt����M޻��o�[}����F�,��'����ͻć��ď*A���Rt�-^V��$��%b�p��[HA<a�`� ���tܢ�K��щ�P��-!l*1AF��lbM����l�=Y���
{?�x�=Y��k�
h1o��Ĭυ4�C(�"E���T{OT�ԩf])tj��u{#I���|����) �֬�~��j��|D"R��<�8���8D���M�l"B$��ʼ� ��7S�(�i>�϶լ^�n�ﲹ�l]���{��*���F��* �:�et�볰<+2O�b芚���ĕ(�Q	Py���P��}������ȳ�O��)<x�[�aǇV��~����@���4���n��*�
��5Ͻy�B���4��*���{����z73׍ghq������K������������E1[���
2�P��  ���
��b,�F:� E�Rz�A+0p(��\`��y
(]Yk5����C#��jV��!�׃V�q���#�g*w�ξ(�/pW�j���1�$I @�3n�7�`�@����D�;WDP�@T0�	%[�b)&l+8�b76RT�	��U�h�\�	~'��}����N�25�6��~��	Z�"�	"]��l�
�{��)T��!@��t��i��#Xf��`�
@cy��4@C��-hs�v�n�p�{_�U=4�¼(��8�2�M�[S�XN?�m�(s�5	x.�5>�3��j�I�z�K���O�,=f�{���'��=@5�\�]q�P�#����JNV]R�0��V�V�3BP�t�����^_B&3��R�t ������ߢ��h��t%��2�O����T��^/�k �Tma��0�����?{�J�KM�CϷ��r�若�E�� ������������'���{�	�|�Sx��oy�g���R��޾�gሇ�UM���K:��G�̖"�f�Ve^�~	��!7�l�n[��%�ӂ�-J����ן�)z�+��O7�J�wLZ{Rj���5�X���ʜ �2�H
��N
S�\@�M�Aњ�7Ȥ"(�}ge5�t�@��r�1�A��`�8T��湒V:��}�*�%j�ΐ�E���m�"H���:��`�ύjڽ���D[̀�� �#O�,RD�l1gV�@��5r.�sF))���!R�e�0�-."a`���UjhדX�3���=(*x>V���-LY��u�� ��=�u4� pT&�NвM7
SX��0���vL3(O�<�'j���J�TD  <��:o �%�`�ov ���^rZ�U��Ր�5-mMZ�ЪL�p��Mq��g�n��[Bz��֥��m�h͏��_H}F�Xy�-��׽�O�}��)��a��$	��L77fP��
�����mă�s��2w�v�n��Q&���	6�U�!��o�N�Jj�u5��]�r���5[��ht�ʘj\���AlD���^�Q�2�~�*��~`�L3�j�Q���`���69W`{��$
�����O�G�+����`��e|X�S�
���ޔ|�'$�T�<hIF�kF��PG��r�V�V�̓v.+ֶ�Im���'V���wS�k�ܳ[�u�z�<��/[�]ey�)��ԪI�l���w&�v�@m��d0g(�*��%����6�%P�Q����4`�r�$3����л���ٵ��^&*�W�*ШUi��P�,lM�����Oj��w��(W�kJc�͆ ���Cf�"(U�81B��� �\��{�V0P�Zl��-×a��|Ļ���u��
H��O��T�C��]�rQ�͋�=����v��(��b�.�`���.��9�ƺrD��L��Ϫ	(
� �	�� %�����T "0,��T�2�)��!� V�._�� ���M�	b��GX6�+��:ٻ��5m�*��Z7�6���S�|��β(������h�Z={ċqQ=z�RKK�2��,Dl}�I��,N���9�!0(0r��b��#f�-V"I���`I��7�f���ۍ�<�?`:$�3dN����z��
�:٫��{�����5��x�M�wơ1w"+�[��`�G�����\�3���}4̌��OU�#֌�z�a	J�������9=���G���'�����q��gq�!m@�S�7��T���%����%�XӒ�e��l-=�]����+���f�����j��$��Ic�٬R:�컀&+D�F�¼��,����*�C5Fd@i�DA����2�b�'�f5+�Փ-( R$�FիoP��(2�5��Q��/#c/��2n�G�A���vo����Rf�;2\@� ���l�r�@�Ӣś����O�\ʲ2wj���k=1�B�l@R0b�u��	9<�f(P�le�2Z�p$F(&���d����Lur�Ֆ�R��
�12�����x0(X'�&�-���.���[����J	P�o�Jm�tU�띪�ꋵQz��-g�R�N_Dd���	:�V#���Wg��
��`L�,IrU�TD���*
���n!�-�b��PF 5�����B���O#�-�e	^�@lFT���<'�6N�5׵Z�ֈ��贌����3�L�Z�ZmHͣ�&�+����o�
o��vT((�e!OG�)a�8B�`�7�W�����O�<��֔��|�s�LG��"6q�V�K����YyY�nJ����^��:��*p���T���85�~�4�3�<�ET_������J *5�*˥�v3���k�$9�/!��O����ç�K/�>T
}z�H��'�|�Ki>|���:!�)	��lJڒF�4�Tzh���Bk1�"[�R��tE�uO��V+�����oS�M6,}�[}d}��x��
��!PH=�k%�����(��`�)�X��>6�	!��MHP��D	3� �z�,G� ݮ����,c�f-�|q�5�u*���m�cB��5���+/H� �������Ѽ��x-$R�9�T���9�Br�� 8��ԗ	`A���
)3�
���2z��@�R���RlT-�R0� S��`?r��y�]>�k���ݵߴ=q�e6�Z���<�~��{j��mˡV���Ȧ�+���6*����D���̥� %�L�3�c�j�V��?GS�f`�	 {!*��C@k¤�A��^I2&��0)jߘ�%le�w2�K�C<�<볳ؿ���[;�K<[����V���.��*!��m+��Y0�*aD
D[WHE)���h��!"�3?~�9M�\I�a`!������./���/DH�1����iF�%3�焠-n^�U(��Da��O7_Ջ���׶6'������ڴ��pL��idJ��.o��oK�]�����M��`�Ř��>��9zB� ��o�7_��v����[��/�>����Q誊��/!�Ã��͟+����<�J2�\l�o+�`�D¢Z�E� 5~��$�d�F�-�k�}+v]�D7VX2�W^�J�T����i{�	�槣�!U2�bk��Z'��`�[v��kw�~�%2� n�>�{�8ҌIf$(PM�#�f0pD�4� &�����܎$t��Q^)iՓ�5������Z�t�i�a=�R�P.��	�2$)����<!���JѶ��1FcD@�hID)�T��"P��{�Rޥ*-�K�=�z������(�^�VN��BJ�F�<�u��'5�AD�O���[�q[y{FEP������PB������ws�fԁ��B$���0K56YH� P��8��1�8�ᵕAB�~i��s^���^'���w��DO�ZU��_�.��B^����!��?tf�����0*~=DJ%�>���Ŝ��[�yBN	77Oq�&�֫���k��/�q��BDPR��`���'����'8�(s��4M� ��j�����@M�yW������BS��o���3�(���Bn����\������nșaѪs �_Z��%�ތ\�1�������O��;�����]|v�o5�&|(����������9������<�ђ[R�1b��%�Y\1KY-~�g�7ũ?���@��y��Q�%�ף�(zvh���3!��n�;�@�����7b�線�F���J�Lv�"@z�0{�v@Ĕe��$�P�g5�V"w(3&9b�	%�`W�}��j�����#@JFN�QJ�`��P��r �լ����h�"�(�F�׷�>k��F��Z%�2 �)f��~5\��@�i&���y�R�#�1 F�u����"�!�keA�sQ�T�Ů?FFL� �ϧ�q'˵�H盡��]��8`�ce���4�e��1&K�9��
϶΀e��ʘ��a�:im�|ʼP�T��R7��{U�x ��h� T�ʆ�5T�/D@f�<IP	�o�������c)��%~�i�n�/K��C��nG�V`(j������k�gM�=�S���I�Z:o�v�TK�<"BQ��������equ��d�>}�y*H�#R�8�v�ǓgO��l0������)%��<�\
�	����Gf��%l���7u�,,�%�ô$�َ'9K�@�r����:�җ�3Q��6�h5Z�:;-����)z�LY�u�2]�r=� ��2�������Q��|y���ǃ�+>,����"����]|�o��S����<}ea6��՚��I
�-~���Xr1�doz~d�z���������j-a�3�W��X��L�L��1*#��e���5_]p��aM�5�A{G&�L`����Q2a�#2f�Z
 B�� ;$��5�02�x��F��x����0F�U����W��r�%	���,KZ�v���߮�sk�c	�F�.��j��S�-	�Z7S��pn}�T�JAI�s.AB�H� �(IPf+�4`�ڎA�%F����m��J�5o�HWR��{�'�����e�`�t��S^�g���JʟP��fL'��d��`��ք�Z��e��["�P5LXZ�F��s�X�n{E������9ke+��u�v�1��Q^+�sZ:A��.9�gJ�mW��E�����]��wj���/	5����p���J�Q����R�tx�iNl//��G^�~������ FJO�1��r��a�ʌ�xDJ	Zex�)�sO}���a]���㥯�k�;"��Ȩ��\^c��V��$����z�S�W����I�z�^#3$��6B���?���/������}��O��cߌ>p��������7�v�돤��?U���J:�%�D!ɐ�{2��R��s��r�~��K&o#�j�2 �z-6Ӕ���9x�ڼ�x�h���z�,����|�r-be(b����q,��2n�P��0}��S��j�6���%aFƬ3�L�2c���l�!�pG�C�ц�l ��xF�R���,�z!��OX])t�$����x�,�{_�V��1w�J�
��� �1a@ҌP
B�Z��X )c.Y3rJ��>�gD�F���E)+R*`hQ�ڞ�4�*������S_���5��[h�y��������0+����e"��Q�EiA��iz�7&2Mlg�$��0��T#+t���Ĭ-�ь 5�Ό.!K�5�l�n.�����ڪ�_)�x�ٛAsj ��v��
���F��I�7���W�S_��("]�o���9\Փ�����QE�d�C q@*�<g�R.8'l6#�FpQ�qy}��|�u���x�����}�� �i�8L38D[����	i^�,����3��s���Qp�F��$c���oxnI���J�\�{j5�:+��8n=1L�����\�e ��L	N��
I>�����0=}��}o���x�o��T���%���ax���(��G�|T&�Z��6�	4Z��K?�Lړ��k��S�Qd�� K���Xka���Xv�2?��Kq��/8��V�t��=ʿ%C�6��"F���������ѫޓ�:oAT�X�M��Fւ$3�L]�[�j��z�bε�e�vW���8>@���:C9#�Yp�����S6���εRWt��}�L��n��lb1�w `�)،f�
��֖��c{(KY�KR��X�%�eA��`�C�hQxUkKlԟ�n�?m��
��;Վr���G-�g�hԽ�h�*���! %,^��>FcQ�GҌ[��5-�7�޲��%���q�8�&�ڡ�@�Pڹm
�Ң���[(Gc+Dj��T���E�:/����K�����װ��Y{R�H���3��(��#pzx{�W���2o�C7ԛ���3*�[�@ss@�qq�4g\]]���#���8N3�d#T_{�%�~�d)x��cd���T0�qs{���{�a
��rFN�ĠYd��lRks��t���8Y�;����K���:�������H#���ۺ�I�Z���~���B[�f	�"��A(vn�:m?rI b��t�^��/��>���;�>��ۿ|`
]U������_���{~����h>��2A$�g#����	�j<]!@� �Z��&&�-�D;�5i:��d�V�D�P������e��k���y�H�b:������;�[Љ
;�Ӈ:�KA1��0b[�Q��)����ژT�@�2*�n�aP����lY�(�R$HP䈩�"˄P�B	�C�Ad��$A�%=����!�xe�j�!<d�Bt���&a�1)���u��{+���E��qq���ŦTJ�BEj��"�pE�����焒	4bX:X��Ա�@$BΊTj�
� I	b`��`?�΄cV0�d=�j��P�h�0�e:��I��v% +ͣ�̖��R
��.���?ۗllPh	�U�	`LK)(Z :!ȡ6	1!�4����$"����JMk_]�F&k-j]�
��l����������4�����	����E�֑ �)YIT��ֹ'���ւ����v�m[v�,�Ѣc"]�-L�:�gevF~�>5�n�Y��+;��i�����w�l/����ݣ+l6�4�����f��^������	�b��<���,'�x8����r�m�{5M���#'
�}y���vΔ�q����L���g'���t9 �o�u]����C뫯'��Z~�U�؜�j�$��I~�������������߂����|�o�-�������=���I���t� 5���,Ѥ��-q2B�Y�u�A��ن�W]j��.�`��O(������W5��w�Z���|�$윾�Y��\� ���7}A���[�U-.W։)�M�b���,����f9X'�b���-CY��?:���@��:C���L��E��������� $�Z�o����,ٺ
�nNUa��ߝ%�����D�c�E���m$"d�q��fQ2�T�p HY�&�D"D��`���5z*�\�X7-����o=S<>�K대dzZ�*ζ:XNH�ԖF��=��c��Z9���a��\�Jw�)Ag��^"E! J1_�,fK����rWB����Lw��(�Evk76Hm?��[	(��a����e�`�|v�������a�Ӄ�&�E�5�Q��f��J. �}�j� h�H�S�f8�Q��q����z�-sga�Z�jkKZR��i\ (6�t6`ETPJF�'����#����a�-B���RJ��v��	2�9c�#a�ݠd`;��n�SB��)8��)M�P%�J�!�,,sKe��{�x>I�<Y�;G�����z���c��3���Fw�c/_���>
����:�	l���a.�24-�D"�%A�d��_���y�}+�>�<.}>0�>=~��똏��W��GJ:��Ɇ���#���T�]J��Z��5�^��K�.ٱ���ߟv�[���`
y�1�f�)�=v}rg_��(],����p
�u� m�.�bD`
��jrגd�(�H�ſ�P���EfZj�U�u���Z�EY��U�	a�#�	*���H�,�ea������DKM�Z���0Е!Ж��0�H(�\=j�GV@R��j�s�&��J�zܘ�$"g˼�LP@����Aр���@V�����L���18��ߺ�qCN�����CS>��;���@Kz����q��ǵ�U ���mF�V�3C�2їw_�Gv^�a}�hM;��Ty���"���d"Y�Bɦ���-=y���=�P��� ��"+O�5�i}�W�\=c�)�O�w�V���*I֝�t�m?\��f1�g��i��[_��&@5A���^�j� ˄i>b�#�`�MeZ.���߁����A�f3"��'X�RPJ�dWǨRs�Ob�f��f��}u�V�ק�)�ޟ��q�峽�����Ým��xr�r"_t]]�Ƽ
 *���=.�2�1���O�g���?|�����	�������UzH4g�o�B��$�w�:9M{)Z������dP9��E���U��Xj?������[��7�*rfMU���ݤ����sZ�Z2%���0%�Ɇ���&�B7Nl���i$��5��דs��SR˜O��:#�D��#����<�;ͳ5��d�&�N�������`j�nBAd�z��^/�s�B*�lXw[k�o����[���L�o�m��a� �%�Υ�Bd����T���U��CR׮������x��w��?���Q�]� �����s��vJe�X������֙��������J�+b�!��i��[+�:e��#v-���K^Rm���/�ql�^�:U�
ъ�4/{CZ��v����7BNAulks�AK|v	�-�	�>9�X��*��_���-�R\
3n��|#����)��A�@ ������vLs�������^sr��@���%��n�#�<M�ӌ� ��<�w��u��{KM}ϟ�����-���'��:z�*���V�ja=TÔ5�Xȥ�L�Kӌ m��@Hy�.�����|��o���>�m��'�s5�Z��+���m��_o�������_]�[HI`d�f����j����ZG�5;�ex/����<I����4�y1)�S\��� X�t3=�=i^�T�S+���,�co* fD�  �)b��V��h�,nZM�B��Ų�u� ��h%p�Ե� �p�������.j��[^i��*Beu�u`E�ʢ�O̵%[M�6/}I$�,N�K���B�;��R{����-�c[d��[+������S"�4|���#�\[̮"��;�t��[������?������$��0��.m?�?R2�5F�0��ތ%$cЪ"E����wژ����v��[��Z��z��+��y5"[0j=^�ʹ��\vHK<����-4�ʭA�'�����{=�=w�2p���i���-	�˂f�BK��?`�����
�,(*8LGp B`\^^ ���W^�v�E%<~�m�\����`��y��B����0�RrgS�ڷ�Y�b��������c0���g�wΤ.N���Z�ʥ��yYRs:Bw3��X�s�:��BbslFg")��ռ��o��o���o������k?��k��U��x>���%M�?O7����3�N��*(���-RȐ�@��̵��	�^�J/�ܵ�[��?>�b����+�6}�y��^�:n�ĈȨ��C��3O3í�zS�l� ˀ��	܇*�c��=%Q�
q%q�����-��X&�e�D�D��Źև�d4X��Xe|��D ���1ĥ�nsS�G��.����C-�8�d,��;�a�z)W{L�Q�	c�"r1ee��Z��h�t�0* �Y�S2�z���kAk�[�"YF<�g��E"��J���&,���������/��+�۶��B'�*��w  c7
�MR�#@�+t4���|)�Z�6��3.�	]_Ok'[g�3B���@\�z[�$�W+O\rmM���8Y�t��Pܺ2R�`�$���s󱭳�X��'�:�V�^-�g�>���������c%�|�*/8\�v�~� ���<ς)%�ĸ���؁'�����g��O{1c�6O�@a{�E�)'�4W�_��C�Z5rNo����؋��9�876ϙ���`w����l�K 3�E�V����$����R��UWC� (׮}���Q�ux�J�v�q��l/���n_�D'���B�����7��ø���i>��r�}%�#4Y	���敷6��(T4O�� n
�y|� �y��Y�Ve�R�W`�Cz�����5�� ,�Ks����l�1�����W2���X�dS�T[��hͺm��)�*���R�[Y��,�)��/��QɹR��h��z��&|c뭬�<J[(,Bz�G6���F;wA�9�VZ��m;��aE�v؍�0�=�f^�Q�1Ty��̵N�j[��yW  �lSڄ�����Ҟ�W�z%(��g�M4N=��/ܞ�#�t��m��z3��Q��5��S�}��Gh��"���޻��u���mQ`�z�5'$�RCkW�/� i�EW��]�=��]W���q�qzv��\�h1&{:�?�x��P#��7��|�|��[v�H�3�[~Ƹ����
yP�h�x�q������~}�5��?���/ �#^}p���#��<��^��ZA�5\rz�~�Ej���ߝ������P����R.w���@��3�)úGl7q����rv��kc�'
f�5�3�}T� %!���a�o�0�Dz�~��e�5S臧ORP��g���%~MI�������l�W�7��׺W�H��@��Z��N�u�,�RA����thZl�5����l���n�s����A�6V�Z�VJ{%,�W)� L�1�ujS���K�w�w��ʭ�����ɖo�;��PK��("�4�Ig3@�Y8KD�h-t#��m=�ﴇ�1���N)���)���Ӻb4*�F��V��J��Xp9L8@��c�
e�D��@�mp,�[IlP2PR3�IUPuN5��L3�d�T��($`�`+�w�����0B5Ygi����fw��oE�'��(�n�Q��P��3�����H#Ѯ��	j#F{�{�F;��]��(� /���L��Uᮜ��̴�s7Lq�����3��{�~qB�.�C��������j��ɯs/�u��G�!+����f�� ���BHHl@#A�`�[�������px���$�ݸA�{��b�C�#J�� l��jr�����ս�By����֖na@�y�����V��v�Ӭ��X[1�?YJӈ��p�����}��Xߤ��æ��bU�(/}Z�	P������c�~7��I��;�<��0��(<��>���|��5Q���u°�����u)�H�H������*����Zfh>2[-�m�:�eQ*�x�zB��E�%l�\����B�8�N�z�Խ�J*�+�2j��Qq�Sl[��*��6��D�m0{O��^��%~�5	.��` #x�R���Q�����:g�!����@T�"KX�?��Go�-�K��R�Ӟ-k�z��ۮ�e>].��ϻNAl��Vf�c7������B�,(��deL9)��W<+��	`%���[��U�)[׳8 � �8��J�t�h����Fo�z摟����t�N֮�&
W	E�=����Pq[Z��,K�0X�����ӸI� k����:�KkV��C����b{4��L{H:�,���،anSW^]���Ӕ岎��:�O��w�W�N��W�ѕ�������w� �_�aդ��$3���1[\<��������C�Y�%!�'�4c�8N�l���W��%A4��f�1s�5gِ�ߵQW}~}�Y�����%�@ݘ��,]1w&�Wj7��g��T�ڛX�j�3����Y��^e;�A*����*� +7���v�B�)�؆�گ���|��)��@��^y�o�q��%��5��o��<6��o�<���飒k�m��j׷�k���R'��X�;��V��إkTU�k�z��O�6�Z#�v�Z���i��}��鲉��>��%�K�����]���,�@K2�G�&\5���}f2�N�Ϙ�-s�T�ր���5���T D�jMD�D!��p�~w
�a�?|qo��{�j��Y��H�Q?���Fp10v0�i2Y��P̛��i
���y��6 �8@UpLq����p�/8f9)�i���%�4å��N�d���{��('��>�xH��H�ɇ(D`܁�(���6aX>�=}�gs�tc5	�v��s�d �$�#���k%p7��ޡ������<�O��\��rg/6#K�u-�2Al��-$�%�k��� :b��@�C��ѣGH�Ʃn�4l��KW`:������n/A���� F#�	�!C�#(
R��l�6|�:7AOBF����������٭r�� �JݘlFX1,�\�����������e�q`�`��T��7VT���h����*P��º��dk�L o?��~����Z���/��e�_<��
������݃������2���{h�!�6��%n��NK��gh��в��j	�Mi��ePb��\��i�ƾ^�u�d���4[B�	��%|��՜�����z]����k�n�[fk��V�<@1#�����(�ڶj��f

F��P{OB*1E��K��`���TP`�Ig���JR��
}�ث�Lt�+N�c��8�/����}5�̓�{	�:����� l��e�P�eEfE��."@jMgH��z%���ƪ.���v�EF�r�1)��8j�mfP�j�m�.}��#��X�-�Uo��;���:�?�A�ڞj� l�@�:?��,�5Ԩ�F)������ޒ�t.X��G��ZjY��[��^��<מּ��x��~�2�p��Wn�]3��\x�;�|�pژeG<x� ���%n���"l������C�f����K��n�!�	"2vW��!�"H���'dN���?S�11���0��+-gq���e�/���sMm]U̵��-9	�6/�tG�ܕw�k�P�=��Q�8��hg;�:TZ"rc�V%���ԉ����\�N�8|'��C��m�����l�^�없��B�g�0I�0>�L���H�o���x�2ی�>AMڈ�6��&ĕ�g=)���5����qIu%�Esr��k�[8�5��m�C�(��,�f=��]b�+�e��fP�JԖ����J���&�{9ࠊLmrي�V�uB����{�p���
��5�A�x��*�gɘ5�:�f8����X�_U��_.�"er�'���5w
�<gZ�S_k���F&l�a�@
�-KKQ�e�}�51�~����$dp����VZmÀY��8�Šh~Z��}�g����*��S��5�{���ݤ��"��q�\B�K����[-�b�-����PY���áf���
S�\2�B�%������?�~nD�oX�W*u���~��>C����j>G�{�'L�z��\X��J������D�,(qD^~����n��G�o�b�靈2=����T���C#�w[d��Y�g���m��3k�b�D�]������O����,���o!�u.��"�sQ�зOO�[Bx����)�X���S\�?�(�t���"��4B�� ��5F�Ǘ���7��}�ZP�_5�>��BJ���K8<��o,i����$iߕ���iu�r���k/�}k����uV�=	�	��X��!%SoJ6p�=X۸U(�,�T�=x�K���o_�����}Z��OX+ۯڶ�)��H�FU�����7$��r���y�@���Ba ���Y�� k��V!K�5#iFAO��I�{�}z�=كϫ�~�8����s]�ks�{��%[3cc L�T�Ú�D���ux�kB�5����\p��E�ՆZЀ��'2���:L��Lh���{���#i,Meb�yu��)����yU�H�-�hIo��b��kyd7.�g ��n%�������8�`�a883D��?/��ד�֊�q��z�מ\_Wk���dS��l�nF��>�C��@`_\�2n1l6@P� ��S��)��裯���o�`�nno1nF���ţ�݀I "�AD"�.���ah�0->��$�{�_�7� ��쒯�N�a��5��h7TE\�n�hj]	V��8yԶ��O��%(������%�K�@��&�|/1m~p����p��?��oc�|���ܗ���B ��c�� ��b��$y��(�CoʼNX+���1��&��zPa�g}��[�����"��,曶f&]!0�r&S�= S�ש`X��d������s]����ZJ�h���*��Uk+1����
BU��YۖZ��x֚1\=�6���X�u�9���O��{�a���4�}_hd�F�5,z�d����)��\yX�@dB�̢�@�Z�E,�Z`��52�PJ�V�!�E0e ��1�Y��S�SO�z� ��;��4�b��e�W��,���홝@�?�ٸϓz/���{T ��/B����?�`=�{�����sK�wu�"	$O 1Y�hZ�]E{�}���Yb��Q0gk�x��_��c�gk���nh�`�M�ٰfCjb�x����5�,	�c�2� 
�0"�$�#nC5�6dG2 	��&"F�$[��Z����dDkBk{�������p����z�¼(L'��u�Z���O�A���`H}_����'_�F3��'Y����%((BMn��Xcm➅�*�,5\l�ܯ1��Ç��t����돽�0ח���BWU��\\}�r�n��L��'���a+���^k2�f�t'J�@$V:C���VZ���,�'��j։F � ���0�u%���RK�L�4�ܼ�:I�Jg�0[BA���xemC�pk����}!V�$d9�G0cF�Q3�9"R 	!"`����j��q�mR�5�4'c=����6�cD�@(A�����&ݽ0s�Ծ�OA�o`Z��+V5�R4����Z����i糖}]�{u�g�"JA$j�����Y�P�9 Z]�%"�ጉ9�D;a�`�)����% ��CY��`T�� A��#H��~�U�6�	�V�mF��%��y ���3�z���r��� #�*tp�B��z� �<�(�V�&��P&�Z��ԉc rM�C#* �� ]���s�#{ُm���yl���r֦���L��lu���̩:�C���+�w�-���ۀ"�kC)1bă��\\���"4���1�@1�Z����e����K��x�Ÿ�8Z`�a�NV����8��3�pY2қ��
;��3��c=F��e���;�����`�:dy��B��UUPX��"�Vm/"�*�ɺ8�8�"A+%���t!՜$�Z�.3�$3q��C������O���ӗ~�����*
���~W�����=�]%�L:<�(y��r�^ �6 D{��� Wk�Q�2WS���|AM�iZ���[�7�
��8��h�!��$'��ڗR��A�4�
z�u8���\���r�%�ED�D���w��/h�}{r���D ͘e��r�Q2
8�0�e����5bĀ�G�&h<b�J@Q!��Y����g^��	E%��xe��ŗ	R�ss��	oX��~��PX�˒���c�e\k˺�V�96�U�����z(�,� jT��J�c%��b@!b ⚓`�������u�<Z��XM�"��"��rPeD(�3D�?=�w_H�%*�)�a��Kg�Seֽ��Y���������z�L�X��ژH	��^�P�Ӥ I�f@�w&K�$������Z�bN��źr5���^���0�:H�e��/��JB�7w�m��%����q�PhZj�@5 lPK�^c��lm	ow�QA����T��@�݈a�S����4^��� �(GP�QR@�;�������؎#<��	�no���*y���"jȤU�gW׫�yzX��	�ȩˡ&W��'x[����T��4�~I��Ő��˸Vjlom���.h�5"V��fК|�0Y*
�ĕ2���s5H �BTg�#�y�
�����r�����_�;���W\�����{x��s�����XJGk	ZR��[�[�c�;G��z�z��S�;H14���_8�R ��;�0��и��j�se�`od��^3����B�fL�ק���>�s�qO~L���(�tƭp[�أ`��ܺYu@��D	�D4��:�qd2CI�oy��b��TD�K��^V	'[��B��E+[)��z�p���K_���Z.D����] �!�ZՆ�T&�ƃZwd�gE2@���])g 38k�ôE��|���bh�s6���j]�kr't�}�֛�t�\���3�Z�J�`�� ,OČ�Z�ީ*To�NU�������Z޵<1õ4�.�y����~��>��A{ц��W�%�� ^ga!��Ujg��h���w`����Tp�zߵ�'x܀���K�p	�> o^�#�� (yh���ƈ;��+\\^�ٓ'�}�� ��K����MYS6��K'>c�*=}O2kk-ߜx�]v/����J�tMO�֏^k9�Z澨"��Кoo�**�(R�b���~�"�4!�J"�+��_�������S�W���WT��G�X�����9O�ߓ��<�!+���;ݞk��ORU�u��������2��շ�w�P� o.�����6h�(J��4C�h�1�t�f}��)���iC��{a�k�
^_�П�Da����(Gܔ=����q`%�8D� REfhIȚ��l�ݣM��楪��4%�C;�;UL9Cj�j�*],]�5���-1���Ig����)�JǞ��1^��� _'0�L��4�U�}e-H%#e���U)G˒堰��R�X��@#�1I�X��Z��R�ʓu���eo�m_����^+��{>�*�v���'B�y��������u�_3��R�Pb�W>�>	�<�F����a�6��ySpP� +��0ԻE�9�痽z����w��R���=I���ܫ��*����,�oz�Gݓ��e�}ev5.�1��L�#����+���a�h���T	2�@܀��|IO1�Y0O���x)���4(h,z�S�����yt槷���|�3���n��$Z���uiy5�_���NX��<|[1���;_�c��٠�Y�͗0���7��O���>���q�_1����SF�8���������f�t i2��+�d��9�ǘ$ϐ2e�t�tK��BO�@�h�vYy�-M
��+��)��#��5#�($g��OG��4�=lИ.4N�bP�^�꽓Y�}zS������ϧzn%�I�*�t­�q�G H<`�������b;4��	�6 rDd�Ԋ�l�e�pT�̄X�F$��5 �U��V�є����Z��J��=����B����C������.���w���B.�Bj�C��:u�fl���DB� .@V "
d��ÚpX����ө�J�4s�=�(���N���k�^����-9HWR���s�k[Ә��\�V(��a؀���J�Mj�j���Lm�*z,ݘ35j3XܝZ<^�|tB)�� ���л��y��e]Ob_��M��g�<ɰ31g�l�K��^}�RW�R;.y �2��'T
�9ˠ��_�x�1��'`�,Pw����Y&��$=��^B9c�#�e�=�JB:�.�V�Z�~v�C��qT��z_6gf����	�� z��I��>��UC�-����K�Ӛ'�T�75���H�U;(J���}�*4e>��0����DM����-�_����W�C߿��=x���������%�oAe����$��s��o�&�U�O�&��*o֚�~7��lr٩��#�C�\!lV�����!
P)�$h��!�(M}-�q�����z=,�)��qy�����zs����Տ��3-(:c�#�2#�BÀ�6���l�Y��1R �`3�À!Z����AҌY�L(�P 
F�ȴ�J�QB˕^c��~n} �IF�fdQ�tv�������U�]Z�)���Ϭ����j�DȢcғ[k�{3��%bY|��]�	<%F��5k�����QVh�R�GPb;�3�=�q�J?�<���kUg	�M�4�5�EkExn?�ӪҀB	d�(�:�������KfhJ�N�#k�ޛB��5]f�E!�*�v�5E�l_��l�������-�sf��8��טr�js����]�������,4�;P+�ۂ�0����q}C�a7� UwU����C[ JI��.��2c���&Y&��ץ5��2��ē>�,T�hw?�51�^�W��./a�u�%��yF�������-��@��Z(Hebdɛ��[������ H�Q�ï`
�V�^�?�O�=��)�_�B����8N{\���w���������&+��Q�g˾�t�J�ݞ34�2]��iյ�Y�ź��5����r31B��a�!l.��%4n!a Q��>���9� T9+d>��	����#\����k3�վ��ž]Ss��5�B�����[րH��k0('CDd�h#�`cgE��9?E){�F����2�L���Y�g��%wn�<�~�p����ڳo������[T����]^�b���]�;Yͧn�{�� � �ܛk����GjR����5-��W�ք�TC>R�q��ޠR�M��I�{��ŕ[� ��b���:ɮӎ�ۭQ���]�֞�B������?��Ѫ�[��t�0��V+�D����JR�&{N�l��➽��*O�>�}}/jvr���E�S����k٥%��=.�8�J�a��3�1���6�1 V�j��"(lL�ǫ���3��"Z7B�2mP;�Ae���sv��D�%gD&%����F������,t9����(xj�?�:t��e��慷�������M�6My��n{��1�Y����s��4MD��)���n�W���_�2�_�BWUdI@�1���y:��<��|�A��%X��kY��i�h��"ٲ�A�M�W)>���8n+{Yh��z��F4��<���ф	�fٚ`�Ƹ;h������o�iM����~����Yg`V�������"�!�k؁,V��\l/�9���`���l��aB� � �
�"b�V�"������_�Ji�j�D��/�a���]K�[ؖ�O:/�Y�%؅:*%��߮��b���9UO* !�1�����b�T���꺔�\2rQ�"(mR��b� ��L�G�����Ę���ݧ��#��#�sݱ2 @�HW��"�7Cc���<�P_*j�[hآ�����j]>���d�G{MO�%@�헚cCdm��(4[��h���P����FX]�6ñ�Uܹ��ʭ�n�2wd���㉫�iL��]�ڶ�&��!�(�J���lz7��IA��C �<nA�N�Bk������9��:T2(^��^EH�1�e�˴ǜ�eo3!<`��,��S�ķ��K�9u%V��ͳ���sWKN����������約7��-��>�X����{c�qҦ��\��������;_5�znB��f����V�,����VAdά�iSb��4�G����o�q���)�W I��V��e�ovWy������曧Q�[��7ŝk�j����(e�JsՄD+eVyh�����e�}�Mp�	���r��X�h#)����-��@ PV�6\�BW"ê�4�C^�U��v��-T�]���x�)9ka��D3ـ�Y
�*�H�L) "��1�כ+��Z�Y�(�ՃHFQgt� �8��8\#�g9���r�� �.h,V��8�u���������i��M��s�r�u��)�u��B�s���ֽ9=m��H՛�'f��1D(e#��"�6�Yj�W��fBa+��`i�f$)Hj�4	V�:q�3!�ơw�Y0���,�}X��߹�3%�ZW����YR���^�Zk_�uS}J�]�/��ј��Lа��B�(ı
��.(����~�����`D�Y�+26�(�Y�Hd�"A	��4�D�n�P�0��)�n0��n�>��A"X���X�qbʀk���3w�n�E�6",|��MX�e�i�����j1j)ku��Y�#t��$_�>���J�0@e5݂�����e�x�3G��̆IB�	Dl��f�۾0z`�נG�`Kl�:WC!U�W�pe7�$T�~&]��Y([މ�0�DK����ʊ��� �XS�
@3��ٝ����@ �t�[q��O�`X���B��d����������)�L)a��t��������r� �Ǐ�}��|�
}~�E�+��G������?7n���g��%[bKk�
IPI�bY�Z2T��shy��q�U��r��P�%��	}��Y���� �n�2o�e�j��P��נkņ���Uٮ�
��̛'Z�O(�R��;��VoN#v���K�-��H�1�#]C�D��4�0!)��_���+�m_B
�y�})O�*�*��vTkg�zl������2��̚Ʊ�&���)��J̖g�;_�xO�[���iĉ{���m"]^�ȇ���rm�	�m�������)@(� ��qS!LaNQFD0���ϋ�G﹧��:���Ӽ�j������`�7���E!ZZU�R'd������F]��~�c���X7�hQ��/˯�gY�+z���;m��RkힻS���J�8�ľ�Y�<�U�~lʼ��6j9��Q��֫�]�(Ue(G�q x@� �@���!8�`b���Ⱥ@��ҥ僄Z�Z�PH�t�q���3Ó�ȼU����=+�?���KP���u=4���Ժ$�M̀�Ϲ(��%���Ͱ.�i�槳]R���s�:�ψ
Y��]�"�&�3*6���QUf,g��p������Ӛn~��/�J��
}�]��K���_�y�w���7��3Hڃ�T��%���uQS/K+y�d��*%���%��[u��q����H�$7��uh{��(Ѿ3M�1� �q���Jn���@WnX�]��Z���(,_?�C[2C�J�Tj�oD���n_��h�<*
���K&<����.no'���\?|�_}#.����� '��|��6�*���v���=��(��4;���"��k��=�y_g����w~�_Ӄ�R��֫-{?hM>
dT;,���0ԟ�q����T�dƜ2b�՟�Q�(mV dUL	��!�J��w/�ݽ,E݇�����z�!uo�����ĝf֚�@�lUzS�zl�җ��t�^K3i[\�ACj65$ؠU�J�����ݙ�:�]IS�R��T��\���� �'o��f�/k~���)@��~�ү�gu2{��ٶ\�
��A�`D�&0���İ}�x�b[{T��=�pUv� ����GFjܾ��}]��F-�Z+\��x9�kw�m�5]��J�z;d{�b8Y�~�Mw*�a����re�Ȫ$�WA��q����J���n�递 &0��������2t������N�� ^��U3@�f���F�=@��䧆���Fn�z��O���|����R���q�3v����p��N�gߕ�O��(�M��*	A������ټ�R�I���.�G/�g4V�T�@�p(�d.�����Z�0�!��oISJ�8�������3쯵�
zO��[6����rP�
2	�����#<ܼ��p�Q�\;d�FTk3aƭF 3T"Bq��^��F���8�|���̄��;�ᖷP�w����F0��֔�gZi��͗��ti�Y���^ѕ����E6N����D�Y��"�����ǫ�^��+��	�h�~�t��l��by����y�\����\`C5�ص[��%����	�j|ϻV�^[&/���U:aIN�����2j�T�r9@C=w
H�B[�)�ɮ �	a�h���@��|���ߡ�K�]IQ�aս�~�������wQ�m��{�-���yv��:�FS���/����:QD�׀�Ge�F�x����h�
;h�����zK�[�ZC)�0hI	AG`�BV�sҜ��,�\�z���sسW�궩
ͼ\BAf�h�R`/Iu}�I�f q �h�kA<Խc��@����e�䄒&n߂Nπ�4�b����W{�$ɲ5j3��,���Ԝ��᎚@K���%���Ų�e��
�2�Oo��_÷��4߼���_������� ����r���|�����c.�H2��V�-3��+b�:�w��@b��J�B����_� Ӿ��M�8ڃo��Ą1T���E,YAD�5�ɳ�ʣu���E��J��hu�����hy�f��UA�bY� L�_p5<�[����%!��X���v�c|�Ww����#\�+��I¨#F��[ڢ �uU�4���Վ%���{͞Nծb����ђ8W��~Ч8�{O`���g/	;m� �j���r�C@���`�b��U1P��f�_a�Y�<�T � ��c�8��V�����������|ߟ�ö�jm,.�=��ژ����<����51l9�`�6�7 �y#��U�������ː�u.�c--,�(o �ސ�V�s�2u�x��ܗ5X��֧1�u�.mq�uX��?S����o�K����q�����Vi�26P���%(l���=�$l��^�kv�ld�ʭM�D�\�`�ɘ��Ҫ�5����Z�l��ץ�b��Y����R��A��� Es]s{��֗�r`�#�"�:G����aD/�h��1g����h�Q(���q@>��!T���ٺ���:���ۜ�����v��ԫ�o!HR��9�����h�%���̓7�EP?�(�����蛦�����x�}6�t ��h�2�4�Ħ�I��<uz]d��X -����i�G�g���V�ڽ/��@Sb��K�U��%�X�\����6-�5���Ք�)NsG���P;�u��N��^p,��#(J�]�jз��x�6@���C��t�`�M�Q�q��f�!��������!���f��y�m� Q�Y�8n�[�[�6(�,m]e�����bG��:�tM��d �~��R{�B�?gs�ΠR��ɠ�E��Da�Ը_�m�U@����ݰ��fkS��(C�"� ��%P����F��_|��9��l�Q�N;�R���r�˄���ӳ|Oּ�Gܼ���^Ŧ�	��b��[� 6��8L�o�PZ-��&ݨ�S&���04^@ɼR�r3�J)h��E�V�v��N��Z�Į��t�f����l��R3�z�0��%?�Nd�赗,	�=L�.���aİ����#4�P
�!�#��5��Fѿ��u韮r��[P�@����� g�L�4��^r5hN��b�-�ag,t��Ka�g�*���#Bl7�@W��}1#�!� !4A�#�a�8n7W���:����� �`	�*�<bsU�RP@&�t��@Q��Ȼ����/���;ZbvԚ#im*ղ����9 
K�.f(���_�a���?���Gt�D��!~�x_
}��	Ⰳ����r��J�?������2=��E5j}�>EU���)�˽%�L�[)��˼���baXL�y�Mq.Y�V+�F1J�#Y	g(U��S�U�Cj̿��!e���ZXh=���R�²��O�V��)�ZA�����Z�
-�&�0���1Dly�_`�[l8b3�@6A��#X(%Ϙ��WyM2C��pa`/�ܦg�ϏqC��q�0\a`�:<Q� �ڍ* {BU�m�(P��yH��@�x)O��noc�f՛����/��Oz&�:F�|�r2u�,Gf��:8F
�d޷���B!P�ҡ�	�)��4� b����YB�Bkˤ�D�ʬeX��
�T&�d��=��߶>ն��WyZ�׽G���'Dj����� 3ۭ�0��]j�3�P)6@f�!\>��	�fH�}N��@���Qfh$�m���k�w'�)�0�(K�s����,��:�ê�
y5�r=��i�Z�/#E��K��&�j��=I �U��.  � IDAT`,�� l�4����/!k�����Xe׋CN�qX��j����,G�t��'h`Pe/�2��i�M,`)uݖ��+c��������^�ꥶ��v�\x9@����7����h?0���/@�7V��e��h��[�TD���9Ȅ0[h�ە�Z�v�?�q�on�<�,)��ͩN�@���Z���T��#���4��B���*�..�'e��R���/�S��|�"���'�V�?�e���� y�"	H��֞C���tD�G���$V�2�)9Z	�����ĨEi��]-�q�J��"�ʹ%d�B�tDψS��ob%��>���j�Y�f^oՅ�0gT�ԕ�m�R���=�6`D넮��{�'#CsDF� ���]���-�a��.0� bE��(e`vd�DŁn0KKƠ���%�7�P��K��n�4���F1�0"���W1n_�̚.jG+dj�H�VE_U�H�P��-�V��BJ�}�P���dZ��b����P�X�ݩ6����C�f �Q1cGT0�3�K���)�H��Tg~�	(e��q�3�9C4"�F�b����{X��b��rY!ZVa��K��y�E�/J̨��T@)ٌm4��~�51��lS5�T ���v��
� ��I�#�8_����j��@a��Q��Q��ٔ�0�6��G�}�1`��R�ڌ���՝���?�����@o�K溶��'�;�P��,��W�Yz�=�:>��$&؋f�����y@�=; lA�L���
 c��V��{Й�׺N\@�Vהn���5:���hA��4�\�"�%!���o��CK�DN��� ���PB�E�uJ�v�0�Ȕ7x��6�6���ot0�Zg��/�Za@V�Ҟuի!@�����yzѣ�Ij��Ѝ2"��n��2�L�T���\�Zե���J���FD���nC
�P �L�8�/y��u���cl���� ��e�|�. ���4>��k����_ȇ�����2�@��!%��y�טۺ,=zƘs����|��jwUu���v����F�b�8a"% K��A�� +	�eǎYF� �KE
v�H�\b.����۷v�ۮKWWWW����{�5���9���=_Uu���|�m_֚s�qy�ϰH+
�T�����v�Ik��#��#�8�O��9����|��yR�*脶^���?!��P�IoN$3��G�Y���Pܔ��ω�?���^�D�M���u������3���'*`%4]q�O��Nt��`)x��>��z��b�{]�����U}��5���N(���5N?�	w�.��_.攈Dy��oƙ�=ݢ>M�7��K�X����At1�~'��ȕy�g�>��
X��+�T���dI�*�ԂR
��
X���P債	.�a���Ѻ�cC��l�[�L5����d]�Fn�A����@�r��
=#x���y�Y�5�ܨI!0J9A��`x�@]l��W��c:{!-`-@i����<~��~���}�����*�\��r�K�<2�?䱯���'I����F����)�k?�����hj����R����N�M����S���9l+�F��H}��8�L�R�(�W�z�l�`Hc";�~ݔ7��'2�W��+�\�i�����@�D[�u3�dl{����3��1�z-V���p�YUp�%��@�dj�U^;����p~@_ΐ� }�н�]:&�n�Yٞ����$Qs�qꌲtD�l�ҧ���gk���Z^��S�7���o~�~���(o���zk����_���x�3��B�+>����{~�>{�������m}����cP��ڞ]_����h�
i�'Y�WF�(��U��m:��c�8L�o�`S�>~�YD�P���"�?S
�Ջ�ċ>�<8����sl&�Go�8�Ǣ/�]��W�F��v(���0��$0�**���k{�����-�3

�r� ��� R+XTi(� *�V�Vp���k����QO�Q�/��e$����y�e�3>[߀���v�"ɨ�� ��+Я��l���T��aN�l���X�`��T�v�'}:_9Yf}6�T�sQT%q+F�z��өb�\±#��B�k\y��Uj�o���1YM��d �z$�4�;53��7��ʹSߡ���y������@�,�k�xq�
�g�j���	�ɯ����b���f
��=��� �s�	�}?	@��@_����c+G��m�Q���ki3���=��$\~/	�AB(����]z��_�x�y��7e~b�J�Vh�B�3Y�l� �D�_��'�t7:d���gg��+P�\�(�-��R���y7�i8�#]�'9r����bD(*)tKgٮ����ݧ3R=jq:�����s.���R� �6ݭ��9�����b;����#o0Іw�x�@���^���{2��z.}���(��Q�|<��Vl D��E��(��S[�����_[�?����G������b{����_no?zC�\�oQޠ�G_����}����z���������mO_�L~�>�����iޮ&�="����}p�>�h�xi�B��!L�f��3Y%���!w؄��Yu�a�/�x�<��!FL5����C�������^�Ƶ�u
:�P����C٢h�q�
��q�.�l\�S�C%,�ONjF�����l VT�(�g��	��8-�V<���'c*�>�ؐ�uW�����]��q��mX����3����"���ZO7>o��G"���C��ۺ�p��,X¹*^UE��]�5�鼸1�>�a0�T��X�������D0�*�p�B�5�ucT�j���QDy�����1�a`���N�Rw9����G�M,�JJ���:Z[Bm��nV��c�:W@�@���i���>�y������ ���v���A�R��@�6ɻ����&�:N�i�t�T�s{���<����á��u!C�
iF&%,��|��j���޷�(�>��@���$K�V�/Nhå�������<�@#u���P	=���+4��ܩr�~G%	¸,8���(�.�֝K���
��d8�B���+�Ā�[�:�_|Ljj�<9}L�#�iԳ N'�,
�t �k���j��- 䱫���������|������!�з_���;_��7�x��[����vy�ej�_|x�/���?���/�?��U����7~���Y���j����vA߬��*�;�wHo�	X��f��.aT�O���?-��yzꇈ�5�no��:��C!,���\y��|��=<
��B���S�N�\8��D��1w�����oq�����N�)�.T˩����j���
����	[��, �"��(u�¦^��k*��,1��R\�:[r�PyK�U���T�T�6��9��P<mh��ޣ�RQEK!J�Z�-%�v���kx���qQp�h:�g�F.���лL����غ�IW1?bEaB!E�B���^�)�`���(�Ƙ�����ķ�U-�B��x��h~A�Y�$�{ 1��4蝬����
�#�9W�� �T��Q3��D+��"V�|��d�� �+*���;�A �C4$Ip3*�G���|��v"BQ��݃�ŏ����Ӓd��X�ݠ[o�BG+�Re����A����/<�L�"�"@{�^ߠ���-����O�iUE���	Z6_���0E�z=�s'�ȓ�2�"3%�rwh��Yg�^X}It�qW��f����NP�է̙~�I�	��5�P�N6�7"t���� .[�hD���}R�1נ��S�D���P�h���������S�.��?[ϯ�����,^zԧ��sr��W��-Z��]�ٷ�K�<�}{�E^���ڟ�m�+z_����B�jB�F�!�iJ� !�α0{���� �yM%yH�U �=?���f�J��U �H�����T6Po`�J��ny�~LQ@���ï���L�=�*V��	�����ͪɹ��&�����L(�����<��S�����v@q�o/Ox{���U.P^��g�͊�z�sa��/c�*�Q[K�p(��Z�	`:�+�@�9?�����쫥H��6��A�1���G��ɣ+���X
^?0F��3"h�
R��3�R��pm �Tl1�\ԩ_G4@Xj� �;ZS�n���HV���1�?8e�<R����L��t�FGEj��܀��+Sqv7�uq�n/1�>=؜t�|�B�����%�w3�_�hӣ)}=;������8}��|!�(�o�����rҕ�H)��ie��������̍NKz�N=�
��������uȋ-%{:
�A���3X�TـM@�t��i��>$�hϠ�-�]��[��d�-3�Pj�8�O�zE�f�E�����I��2yd�n_<���J9�Q�
݌��r�K��!o��y��p�v*d[	U̹��Es9�2���r�t�����
�N�0(�h@�����;h GsjFwN�X�H��a�=9�*5Eӭ@�?�^�~n�G����7r����|�>����ǅ�PW\���7��K���|zD)�ԧ? @�'H��Z��v���f�U��l�8����~3�Pv0W�~��K�1�/�̣K��M�y��H�)mt�x���SRoW#�F*�F6	���+��񏾧D#Ű_�P&,���wҨ�Y�DVi
Ewv�M�6<h��g������9�#l�.�1�D7@7+(%2��ޮ|�UW�z�U.h�rmD���R@'0�<�e�`DE���M>�P�L����f�5�
��٫��<x�Zn6h���5�@�&HY#lq��P��2�
����6�B���{�s+��������G���	��
ҫ� �^�'���$.w"�tTu؍d�:<>$��+�O�x��&GA�k6�tre�� ��٠`/�R��|Z ��O��y3��VK�vg�}{��Q��-���|h��R-�B>���G��#�6շx��<p(��&+���ɍ�ʒF4Y\L?���m�t�`�Qg$$�v�d�]BP��q*S��B$�в��o㍻��o��Z������V]�b+��+П����'k�9�B
�.�ֆ��f��r����q��M�hJIL�H��(ȓ��BE_�~Q�lЭ���ë�q�aNw��`��
ft�X�����LK�68!2� �X^}�V;	���(���Ay"�!I&��&� %S��(�Q�t���v��m=E��`��p}���T~b9���?/��~��X�y��ׯB�!�l��v��_�"��_Ƨ>�Y�+DXW`{F��]�_[6���@�8,���10o����(���BD���5u�a�H�d0vB�1hͪ�IɊ�8f�GH�j�$�Z	Ee��5i�4s!\��%��$�yq�,�6�,L�����U�ʨ^ ˂^*6U4o���x8-hz��
\����9ٮcE��\�[,�!6UlҰ����EE����S��&`w\�v��-9!r����Q8-ֶB��
�E �cU��j��@B ��H�;�Ժ�dC�M�8�ՙ�xR,��Ʋ��]	�z�e�@W�R�h��;���@A\�PϠEAm�\Vh/Xj�b�z��6ԥ�C7�W�mw�MC~4!�(�DH�8���0�h�8!y1�.(w��j7���xP�ttS�tk� CB�-�0PJ�/�yO�����#X���ryB�P��j�_���1��yd��G�R��ܣ�(f[2sVd�c�]l�FW��2&��\����ȟcgB�{���Hq�s
�21D����m�mC����z��S�p�J��[�R��j���ؖ��2������?X.֍kueU�����l��:W@����'$�d��,7Q�A)��(
u�\T)�5��2G�: �a|񔎢A���Д���Rn�F&�Q'� 1C��RP��&}�ٺ^A�
��J�K�b�������罭��e#`r�4�v�b����j��D=��T/�44R�Z�:$��u]��"��g�]��<���6-˟���oy֟��F����}�����2-ݮX�~��7~	�w��c}�Lܝ�]�p�{qlD_� %�KDgn�)����/�!�8 �)�����G�Kǟ�s�=a#F�nހ:j�4�����{�O�}mx�/�����~�4�{ ��;�'�|D]6���+���Sõ_qٞPE����	B�k��k���䊭=cӆ�b��.���(Y�Ђ�Ū޵����W��A��2��n4��>��0JF=r����rS�JT��`�TL4�,c@��٪@��P� ټ�ETr8�Q��t��(l~�L̌�i��E
����BN�NaWb,Ո~X?@W�ed�(���T�z9��D8ג
[I�����FT:�!�v(W,4C��9�62�:F-�XM�@���P~Ƅ2Ph�f
��9�>���w���ޕ� ��զ���d�(8^
z��`Q�|���o�.��g����@�[]���zG�BA�8��>�Z�k!���]�Y�i�&��w�B�1��9�cLg8���N�XJɌ��v(+:YMJ�s�^a��:�#VT�i�n��E;��aݮ�v�yfݩJ1���3�H�<���5VR�+0X!r�&��g�U:��#3=�f�
��kp��qj�@A 
�O��A���f��,�z��CF�;�����5�1r��Ό���M��7�<�v�_[١=Q�n<}��R~h�$��7o��@9�����{������������Q��c��
���;�	��y�m}�~y�����*�p�$._�9�0����c�`��1��&)�o��;fJ�#���o�;�J�Lč�i4�7Qls���~��{�AO�}��_�!� t]��36y�ϸ�g�L�=�\�X��*&�mõ]\�+D��M$5�q�V1��F��`�����
 �] �B��c��(�{����ChV8I^deժ>瘼5���[4t��i*`W+�"hm��r�N��
:Tx��Y��$��	�d[΋1�5�iw�
���h�lmk�O�����(^=���%ИXd�y Y����=�2��0�AK�����A��D ��o���Fa���EUS��C�+h��=��8�+�Π�ЭB�g��{-ZP��gm[�T�
�~t���)��5t)��������	{
&:J��$�P�Ls�3�>:�{W�Y8��]�r��(�E�C9�����a�^���wb*G�f��*�u5�V�|��i����jzK7k�m+�]���]ѯ�6U���M �{�'r=GzpvZf��ᨧ�:Q��2n)	�ӥI���j��r���C�B��zq�9�V?eN���+TZo�����~|�&��χb��lz0.z�?�պE͖{��4�ϵ�	�i����LIa����W���t��S���?-��O�����˫�!���J����:��a���O�_�~|0:�S��F�2�˳:�M���ѻ��m�nu����bFr��LO�/Y��x��$#7!<�8\�Ccj��o9�o���q�Ј�.h�T�;y�&,M*"<`�} �L]]����z��p�J�x�x�+<���k������s��+.�	�>� v�%��Q����̆"+dSl]P��6���	Qṩ�f=: �L�:ds�85� ��ә�@6w#_��y�v�P\Q�l�l�n%JP�jGS��Bj6�����X7l�Fѝ��7lm6`[����	}[�[�R��x�N,`uR*�x�1s���(�J%��K��a*<e��.���9蚽�(@�y
n��[9|��5���<X�Y�n ��H zs�+tmЧ��7_G9 �؀B�ӌ���pxzKT�"�Ha�g�{^�o�L'�����_��g��)E5���Nۥ����hZuؙ=%Aݘ���/��>F�rF^,��`��͸B�o�����zIG!+�%7L����BXN�4(�]8a�w�<Ń&���"�>	���5�T���0j�/�U��08�UBV2tթ�3C�*��qdH���/�kV����ޝ%��9����H$�`����slZ�q�X?��~𖾜�� J>k��������g��������K9����0�z�[o(�	��4.X��'�	''��= ��:q?K�aO���4�&�Q�	H�`(���w�����v�~Sseo�	� ��Ͳg}xD#J�8����c��=]0AX#Hl�`�c��Z���D��bECG�R���i�z�0:z���]m6��1�i�ł��7���+?㹿�S{�k�"׬���x6�f���\��).�D�Oq��ϱ���A6#5'�����`|�$��B�G��m-#2�Rs�T*�&u�֛o�=���E���s!�����K�"��o���n#�\)غ`�����x,��FDUlr�S ��ȳ����i0�|�ff<�N�5�E3�1�<��|5�{BdU�������.gT4`�B�	R��d��-��7C\�+��
m@��Q��).!�e��}��:�T(N���Q(����h\T!2ڙ�ԁ@Gwzt�|�	�TU7��|r��L�թ���q���<�Q9�Ե+:72�aB�\�׷~@��TG>��P_�=���\?�^>�\?���z[����[G[;.��u����� UΕ��n��w��@V����Jwƴ�#�G��m��)o�\!A"dd. G��@�D� yoŃ�pܠ��!����T�����]�@��K>�������Ǫؚ�{��i�z�g��m$��sFJe]�lo��#��Ղӫ�^y!ccr�׷X����V��C���'��:�sB��Ob�(���&k!��6�`�Ɓ�ӚE?쯔�@��m�C�ǔl�X.�`F��C�Q_��wK1��;d�a�v�т��;�Q�:ǻ.غ�/��s����PX��$�njк�k�nxӁ�����{���y�e|Ծ��훸�7`�Xѣv���UZSM ꄾF�����e��  Q�ut�D="Wl~��Q������]�`���r�a��8�0gP�	��h�hM��P���L�BY*�+���P+�'��J�V'S�1ùsAg���a� 8��&̚�YD�ٌ�$0dDd|<���ߴB�:IED�H�n��vf�b�+��YA�`���J�@؜�� /�,'��ڊ�r�"�b�B�3z�,��~��P�+t}��BsZO7WN��<z4Ek�K�Ѡ!O�8���3��[�w�	��
a�ς��fj#��x����"�D���Z����)E�t��z�^���,��xOm�6���<}������_�-�!��IQln�ۺ���:G�r���N�"�R&F����i2��Uy�
{����@�ϵ�N�S�$*T���^(�f�l((��s�[Nei��{J/�3e]F��82qWLޝ.�Ƕ���j����]�\̝p�%�^�J����P�9�n[��ޒl���rap%+n���_���_C��W���HcC���s+��ibˑ�����tSp��{ĳ70����vp���O�Zk��l�2���ߘ74�'2��]�t�˛K)�%�h�t#!���G�	]�C��JX�к�����&�d���
��N6�h�hҽ�Ԕ��/��|z���o�'\�W�b��sW5�Vچ���u�t%)N��iЅ�OQ�2r���s|�Y��#�ɠ�n����hE�J�qL!	��g����~�i������o���� ����4T&�P��X!�n��X�^�:���NU�rfs��N�P������9��t2m@hL�r�����y-�M�M�)��Z*�m�oP�L����ؼj�O2ť�����[����� 0Y�NZ��>~�I��q%���������\&%�8􈤁�Y�&u��mhP�E94�w�z�� �H3z=G��D�Ll�g��'X�@�؞P�[$7A������,*m}���u�� �o�/^Z��ۊ�:�)����s��������m�>H�kBZ�e=�Oq�?W������R�ѻo^�G��!�NX�OT�g)x�_�-��� �ڞз7��Ջ��ta��7��4���#f�T����3n���1��/%QT��@���[��|Ӂ���1C{��.�UI_y�	� �گ��~EU��kk��2�c/R ��z���%�8����ɥ��*9�u���P(1���!sZ@T�Z�����
�9L�^Sю7��P_�(�	SN1�����7����>
�f5ցgB�|y�5���A�����'W���0o���Tl�*�����}�t�mo�XW,� �pU�"�UmD��Y���*!�F �^�D�Ԋᰏ��� �%�h_/0j[��"Y�N�DE��`9��;z߻������=�5��FWkœmZg��j~�J��ֳ���U�z�支��V�b��k3(z��J~�ݨ5� ,rX0z�:H0%�Fp��N+F�="�ؽfa��C�ʚ�*�6(��cR��R���Ũ �~�� �0Zˏ��@V��M�������
*����庁zGc�d�AB'��ijhHk@5+jjT�Ng�9�t�����N9,��u@b�"�������u��8KF�dϑn�!���sC�J	w���q�C��P�Ů ���Ӗ���U6P{���/�П��X�'�j��-����7X�>�N��>w�U�}�X���s�7�8I��S�}��U=�:8�^�z��)W���J
)�*�6%徏��{K�=�ih��M�x�{��R"ڡ�f�t�v�����}��}�� �W��͂T8\ng�F��u� (ڡZA�H�ϐ��6���^W2�,�hc�à�)-ÎhJ3�e���eQk{]��3��a����+�Ӓ�i�S?���RR;F|9�p��0��*��d�`�:`���FN�y��Ë�@�x���y���B�+��]�e�d���!�}NP ���8��"=[��u���u�<9{qQa�@дa���@���5zF��du�Hq��¯p�U��t��64����gT� �8c���[{��dR�vs�:�)>*��d��! ��׾yk�5&�����+�y�F/���+�(�q:�3"�����7��+x�,�o�n[S���������Z��)s'�7)ˬ��H�$��A��ۉ?�<�M%��pBU��]��
Ō��W�h�
�iA� zD�oW�l�A��A�|�z��N�/b�$ h[Q�'�u����xOV��a���1Q����`T#i���B=��G��@%��d��Tq$-ȵ8�S��*2OӨ��GQ��k�:UD�ӹ6��~��QHgU�$�������|hV�.�<?���[�4h��}���� ]��+�nX#�g;����0��'3�9)Q�"f�b�5��&d�Eq�z����<󁎆�R2�F��t�F[.�"
�F
wju���(*���L�"`�&�;i�8u6G$�Ug���$	�:��P�z*Ղ�dnd��Qε��Y06ul�	�	�{�C�Gk�oF�As�-��ذ<DԜ#j��1�~�PD�/�تs��Ugn������B9j��&��Nަ|Qn�M���ܞ����G�x�y�Y/p�u�I����l`ݬ �/\5�s1c���a��醆��l�����*���1D����_��'����Mqך���}'��!M���(Y�����c�J�a,���	��K���}�q������9.�(\mNr��`9�ZNX;akFw{]-�ۚ�DֻN����hǶ�/��*��a)���Q�zm�y�Ԝg�� ��y�C�����n�(�w�k��f�5uj�h���~
*?���`~��^�^4�D;�X�?������������T|>�N' ''�q�i(��#Z�hr[�h���2��a��#�����O�����L�����8�}΅3?&IM1��3�=�0�S�m���ѥoB���6��,` M6���>���3��'�������z�v����
��u�X�ڝ��c���ѻ];��T�	����ޏ��1e�L�F���ӳ�7������0����rA�ϐ~�����{���D�͎��o��C���g1t��ɓ�E�fsS�&Թ/L(]�xGd�Z�;S��������w}��V�6k��+�snL^�{6���8%3�0G iؼ�8�)�d�I�eZ��x�	�U�b����v��`x�Hd|޻���:���	��:�`*"h[б��B��rE��[6UP!H�·&V���4}���7/�s��Y.�1H.f�u��/h�-:@�-@)SMA��!�1̀!�]s8'�Gv:s���ڬMN�ރt�27:��9R=��N�D'��(f�A [�>E�r�u�!�-�
�W��ݎ:�4��2�X��"(�)0���:������:bJ9�#��r*�O�<�.�.ש@P)�#��^��#(��VeDE ��N�
���lx�:]7�ј:�I�@{�<9gy-��P�����#�@����rD��9���z�	��=Χ�L�:�8� b�̓ZtD�B��y�kn���]P�"�����u,����B�+��g��P\�|�7��5\޼�	���u5c.��ʨ�V��m�d�,�Ϝ�~@���O?�g�>nJ=�F�g~]�hO�HI��N[Ic���s�(`����	爴}y_������'

>�ƽD���`�<��ݬݬæ��$#r��Vp��H�H�1���^�nW�^��}�1ZW�ϯ�u�z}��x_3cky#P2�!A2���7�p����ޞjrI�@��Q=ڧj�[Þ0a���g���h� �N؆�}��o��8��M��}�5`{�5,�� �`�c�>uUl�{�T�T*V�% `��M-m{i���
�킫nX��r�"2���M*��:)r^6� �g��U�=� [���yn*H��vW`l�"Q<4+��%ۍ��ݻNQ(Ie���ܶ��nx^��J%�Z,��<GF���ɸ�;YL��'V�^��`�
wDME�:'�9"�@��~xr����RG����[�E�K��k�Hv����h4�1P���h5�U���7��3J=y{����(%&�m��HV@����@����Aj`��	���c��ڤsxR���_��b�U3 ���������pB��޵�Я.S�^�����B����ր�!W`�z��]�,`|��_�}�7�^���m}ݬ�:�IfN�"W��Ϻ N�q�F1�Q�{�)0��h2�����fyJ�>��αWL����������~��m�4�TZ����#-u��)�V�i��i�#�3��_RH�l&�`���'���F�:ə�\�pFb �TjoA|E[?��7�D����M+.�'+��x��� �?�� L8N�&�g�^,v4��q�q���!�ʱ��ا�}���d�!�&
�s�C��?�!�?kD=\K�	`�Ć��+V��j��

0�d)C� 6�.T�Dq��U�EM��8B׎���'yT�o>K�ɀx����'�ݱ��_1��Y[�qs�\�@_�_zL�S�ۖF{���@9G���{������%��;����
<oƿ0Ё���u4� *�xA�hG�M�w��x���<�@���C��H�lǡqE����c�K��u��J��i������70X7�� Z���؜IU�bI�{��=���b3�9W9&C���Mz4c*�P��T��EU�,��ͨ�H�"=셭����%�猼Y� �*'�,6.v��pwN'dk�q�H$�LA�ۆ���7�V
J�3���z��u�mE׎u-�����5�����3Dt�>%Z���
T3���=���θ�;������]|B����D7�zE4������D�ܝ(����@��9.�y���<��`���H�Y�:��p�	lY�E��*�+�������A�#F��l++�ШCP���7�U�/op}���4J)�}�z�ڻ���؛��hIF �t&�6+r�ۚ���ꕂN�p��gwrǫU�w�gm��� � �8�gH��y�q�$��#��-����ݣ����l�\��3?�ay�C=�B�mOX7E�ŋt4�@��)p�+6l�����.];�V�����#�oO�dÎ����S�n9s�d^˺�"*�*�h"ن��E�|$/�MhR�;�fhZ��6��H��+	�>{��u�xz^q��{�a8k��$w<Q	v`�Z���:Z��fc�;���E�P�Aey��`߶&�A�C�����2����@:���
J$����8���(�kcE���
���m.�g����[t<i���h��Qt�̷H���{���֢(����E/i��J�',>hMF)�N��X��Ƚ��^��>R'� ����ʶA��f�K�6(f#i�9SNy�`�^wk���36�Ƭp;c]:�n%W�z\>�׷oPT�ʸ�}�δ���zE�]P����x����l�뛊ys�b�&�#��؍v�Dt�i�<���>(�]F�7��ؾ�������\v��uk�N6�r�Ń���]2�+i�1��8����裳mS ��R�#�Ք3�;WOqG�^�{�u�&��U֯����h�ety���7���uE�T��]!X-R��#��BHN�*�#��'CRޛ�Xe�Y�>)���-�O��� #��I��)"�ؙy�G����"�_'/|�@i��*B���T�E��}�*V]�;p�
����>j}g��~�ju�l��:�l&4:_��8$�s�+mt�.�O����kG�l@�/�w�Q�TGof^�P��;�v�<gJ��D��M�% ��OnZ*�)eC4�e�_�+bk�ѵ���-�0�#�q����V�aU��wl]�MQH��F>�+��3�מ7��o�%���8�*��N���\���Ly�"�X�#�:.�h(�����U�éKm��ϥ����hs��.`}kH�����X	��RFR/�2��ΣݿW��l�3�_@��ܖOT��O=��ߕ�6��|��F���,b�C�1(V��%�hf�\���(��Jg�#G�ԞQ���Ԋ�H+����ס�(���b�aU�`������ \Q�(/V��l���>�m+��NX��uC��|��i��m��z���2��=�O:9�:4�>���{Ę&��Y���9}f��iD iT���II����<�	V�GD�q?�:�~5٭�ŋ;&A�Rk�C1<�L�&���M�� ����H���P��}�m���ذ�5��-�&Q#q2N@� U����'@�"���=�}
Yӎ��Vo0#M����3�-����VF3}h-SԚ �k4�S�<���.��qB��=p�9t��Y�����Q��ݼ&Q5K���tM�v���.����*'\�׾Z�I ؊����s�J2�G�~h�Cx3"��Z�t�[.��V�:%�,(�9 ����ek��̧����I�����z���S��lQ���o�B6`@Ĥ�����ņ�(l�r���&�歞�h��Ώ'ŧ�~�x��R�)��]͔�a�������ԛ��E��^�s�$��k�p��@:�љhR����Q1������֙�0C�N�h�ܽ�ɹ�<r����[�����7ٶ�M�3�����cT�?�+a~f�i�B�ר�>�ң������3��gyu�C�uK�j�q�VX)I�R������m]Q�G����Ӳ`SB_W����Y}r�)z�O���h���'�v5^�-�F v��q���*�}�7�8��p�"�KcJ�HŎ��k�G����9�p�kc��n�|x"f!�|��a�H���Qw(F�v �R�)����
�gڜ���W3��l�z1�<F�`��R���;c�>cY�Z	��h���W�2��kBS=�|�g�VD$��צ��N(��0Uj���X�r�w^����E���Ǩ��T����j�Y���ȧ0k�hF����������g(VcC"��D��'�4���sdv��S�s�s7v|�~�6�<�c�6��k<�Sz8���-��y�zBG���G^��*��=2:Ӂ�ZA\�1z�dd0��p%�R�z\� ���r���,
?����W�K)�L֢e���;���"�ދڝ����;_e�g�]�{A�C�U�ZpN[*-�Gz�X��
b�͘aC{'�Ԣ�;���[ݜJ3�An���UB��;e����3��Y~v�iʢ�렰3���>A`d-���\��o�yK��p�l����k����{�ضRB��\�u3Z���#h[�Z|1*Z,Z�1�Y�n�j�i}���
)ya��S� �w�9�k�N�~"��Y��I�K��#9�=�B$I��Yu{�y�+�=A�ã������������d��5;!��U;��\u",KM�4����fr�ά�Pg5k�J�?�瓳c]��Q�!R�)��p��
$$!v2>r�79����:�C4���}�i�U3B
\w����������;zX''H��/�߾��v��p����qe�צ�X�_�L�TP���{�p��**�ӹ��0 ε,݇�(;ч��|��!w���G/	�⛟��܃�b�9��/��(k��&�s�8�k=}�D;ۻ:{t��Ϭ6uM"kI�����b�GN���Ƕ�'�w>|�x���0:���_; ��}�2`$�y�宋���<�
�\�8�X��[��~��	�V��*����f�[uv�T�����yad�R]�K�S!�1`�qpn4��=�[9�c=0����i�1��4����hO����[t1΅������K�?�
S�_��]��?��f�Sx1jYe����p]ַ�D!q�Z_S%�T�3 "ض��̸-N���N�N�;�`�O�3�e�kh�42L����b���,��`��{�.�����Df�O�32}��A���N{!�h(��:�r ��XĈn���B��ƀ����<��T1)1�?k����	�Bu9��/+�u�i�ц}k���xof#�E	�����+�ً,���X�#{so׀\^vv�abЍ��%όm���ΌzF�:��X���=�2�+`��eF�kְ�O�C�@��\*�r�Xk[�xLAZ5'#�a����v/�2��{kY7��G7y�I�������	FSĉ�[履#��)꜍ݽ��D���q��b֐���F���}�ӁOc���fk y!f�X�U�{Yp����
�טߧ1�B�X�;�z���5�!�8�G�E ��=�EyF��9��8+(
ubN7�bx������$E[aF�q�������^g�]'���ܸ?�=����@9��@�lW���͉.���@��}dlpB�MJd��J��qǪw���io�ڶB�b�v�@a9p�h�:��y �l�[C��Ō�f���d�-z� h��H�Gn�����0�٠��u���b�N�����G�QgS���=�b}8	�:�;�p$�H#-�4;���kĲ�R���:�|P��Y�\^`�Ҁ�#����cumDT��tA�6<>��ȓ�FX�{#�����ʾ��!a�>�������(v�zG�-�_��j�9?O��!�����[>�/�������ތ��E�6 %zh}�l��*��x�+
*��Q�@u�G\�)����$6��]'�A��E~S~Ky�)����3;6-�{R��Os?#�Q������#);X���'urVH���'u熺�ִS��=|�58ѣ�"�N�X���(Ҩd����DбΑ7��Ý�6S%��6�ܽ��2�mj(Σj���g��(�	��`D��v��ՋWI�n�'NŐU[s�h3�mFZ������cu���e3Z���T���^"��D����
*>���0T�����������2�)qA�շT6�ZAUP���X퇰b�}�ذGY,�V@A��Y�7hW_J��	G-��YާDtzɹ��M(�I��Q��lu,}$Ӛ�2 ��0hZ�]�?���o�srgh��=��!SZ0{j����7���m��Y��EE]1~��ʗ�)GG�Fu�v<=]QJ���ds���� l�7-%6�V1R}G��(���	�|˹�������$�6e��gR��ְ�`����c��_�pA ym�*��*gŎ�!���J�y��3��jᵙ,�
1�\7�J�/<���39��􊮴�jB��HD��J.����D��,���dq�=�0�\ϑ�9@d�P��K�s���ư�]p��>W�(�n
��e�2J�2j{ѓ���� a��h"�?�΍kC��3�y����G���(�ʳ�^1������;3���-T:���q�~�Dge~{`�-���ɻ2B��P/Њ����w:oq�ُ��U��S��+8̤KȽu�������z��5��ȿ6T���@�̤#�.θ#���jS��DֱAu׺X�T�S*
��}}F#�e��tr�Y�h]aL�+̰Oŀ;�gBG�3!�߫��Y�7�ى�����|��%�c��ĵ�:M������H�#��\vNǄ��^�uN�Kbסǥ�3��O�km�b���r��G%�R�4��,"��Ya��] �?� �����+D�?�QСX�8�"Yճ{��:Ȟ�E �9���z���v�غqZ'x&�!��"�}� ��Ө�r�3������Ɏ����ع|c|��F��+ht��)��	%��lchO�~FEEe���!��Y�����k�h�{�U��&���� ��z�#Y�]*pf|��l�=�x�2c���Y��ӛ�T_�ݑ�Q�������0�>�n�.X������]RaĴݮPqs�/.��Po��?Ԭ6z���E��U�y�DôKP�F�-��BvSu�vKE8�5�2u����2W�n�GXgB�Y����V��A�)}<��P� v�(i�BV��yĮ��J�w�qԭj^��f_6� �v���3�T$��!9�0�V=��x~N�aLR�a�_����߈ '��ƹ���O���q��{��3�����ڬW���=�b��\�@�X:��Sk���mPK�:�1����h�!CβX��4E@���n�/v'Ҁ��p*Tu�%l7�io��N0tM��Ri���H��e�_�S<�p����b*7'?^�;eb����n\c�.{7�@���`tP�:6����g��W(*�U ��j]Ћm:�a�>�&�	~��kh-K�ة��ܴ;?�S�ŰG� ���Jӽ$CɌ/V��[�/"=���O�"q{C�peJ�_�v�L@!Q�9�A�����C�c�|m!�D�aRm$l��EpXA���&��`��?ZG(ׁ\i�lnuN�b�2�!�k�@�:�BW�4�W"�}�����`����9E�~��制��{䮆Θ�7x�a�a�VKZ�L) -��&����M]��3�A��[��-�����)�0.
�&�������)[���&��P9�sm4*��4����zEi��0���r' �G�""{��
vN=D0��l}���zH���J�]j+(u]2l�Y�=el�����7�k"���K��h)����o��?�t֦6�� əR�eM�3Yx'�B���A!��TA��T�x~�n7���ޡ�c���{1�5K�$��@E���S���6�x>��G���Sƽ������B���tDZ�%a|�������3*�U�r(��@M��r��4x9Bv��m������Q,2L͵��X}�|N�ޣL�Z���* �i཈a�&R��Z���64�C=�������lR��hq����?`���iᮩ�~��_�]��ʬ�&���Q�p�sgOt��p�\� ��s7ex��������|��&��T� =���hS�1�1h��n�]����!�a�"s��ØZQF\�-��7Fc���K:���h}/��������ޙ���"����H�
Y��"Fܐ��a�S,���tϣ��xTw��<B )��q88&�p�������:9eq=Z��¥���vSR�	�*��C��b�������xE8WO�	��N��$����V�fb�؏{����{�{��`_=�	�� L4�ҚFoO���X�]��+Ԩ�/%X��!rsV�~E�(���\,�'>a]7\�+��+��y�fuA=��HpI�2�=�w�3{#{�u����3�����QX���榰�et0P�|KhE�+TW(�DHc����8[�P�M��Z楓]z�a&�1�׾��kN����G�z��� fF)D
Q��EP�BE����EQ£p�c�t��_A���L6�!��@z�T*v�uN��d�(�+�	�@�pw��+���犃�4��0N�!�`�CT4)�]!��w������ �� �v���
�QyA�j�l*F��FF~�̷�X��Ƹ�y�݉Rd�X��(�����J06Xq���;�k�W�ɎG��?���;����r2g\'{Q\x�ܒb�b�����"KR����h��w��|�|�At$#��;kp[��1����y�4�/�-_K@2��2�|��u�.(W0�u����]1:�U�A���P�ކ!>Th_e@���oPF�f�T��5[D�\ݓK+���1G8`���N@ɴc�Ƿ���Nn�C��e�{&��Z|���IϿwtti>�h�TF�6�vу��oX�뺡7A�n��'���3`-�u'g�\$<��u_���$������ڞ3P�q68�3�~dN��
�>��
hAg^��\���q���F9�����A�~t+�w��?��khl�KJ)#�6uT�ʐ&�m�E�bJ���9]bV=¢�d�i	;�S����kG���qgto����B
M|/�!*�'c��^�/>'���� #r����Q>u��x��
i�\v������XE*/(��|oX�������N�9X>(S@��Hr�A@����ɻ�K���e�s�	��N�P�ݪ��G ��d�B�H�P�
��s�5P%�t/C�ja,�`�֝����ZfJw�f�Q<�ֺ��I������{��#�?�H�?�C1xǮ�ńL�=��p��ו�TPJ�p����@���(�6��t2(u]�PS����}TFߒ��DL���-`w�>٨cB�w����f��q�;��RHS �ņ{*�Y�����H����+3����j�~{� 5����k�P���i98��;��z6G�Q {���O�����}���2�hu�4���B��,td�y-Q��f$_�, ��lG�H9	��,�cچ�ܑ��G{��i��U�V�~ھ,��$0�� �]�ć�
zj~���0�à"�ao��W�3G�s��8�)�;d�n����ў$q8�u�q���u�T=R@��F��J$�(�	�q�&%cn"N�C��Rt��(�o!���m�S�*�����C�Js ug|n���z���u�#�#�L� �~Un�B�WE�������	(�r������O��.}��U�/�ϐ�ŉ���w(�c�=Z�cY<;�q=�Fw=S�����Q�P.P&h'��oA�Q��yޝ���D㔎�gx2Q�<;�v�]jfT ��dw�S>:�G9����2��'>#qCF Q��^�}ެ%R`P�.o�v����ӂ�*����e�[Jźٽ�N�Ey�u��zu��,��6�o�Tx��60���uO����������x~��u��۞t�di�m�l6Q��+d[� 3Z*��ܖ�� <R�ש��&\LoG������G�z��t��!�rZY�f=�vY�=�E�Iޭ�,������	�U���b�����|DV�zz��Et��U	���-E�˃9wpq�ˉY�B��5TI��Ü�F���hB5�3&���K����p��{ւ�DN��G$` [�� A��٪�_É�������E�E]�U�yY2��8x��=x��_�ϛ�d�o�ҳ"�?ؽ	f�
�ޞgU� ���e�1p����o��WhF7�KG*�����j��{�D��޼b��(�ؙ���J��k���#6��)�d w��ą�6�e=�b�0N0��c{�c5�,i��a/}�j�=M��ٺ[� `F�D��m�Y�����=�!���"�����@ղN&
��ȏ�����cT8;s���o1��U�^��gU�R*��Y�0���+r��Sj��5��s?#�i�H��T�Щ\���f��
B�>\��1DH-c<�X0N>�mr��Y����i	��S�O)��gبy�>y���)���HTP���X!��l���B��:W/:у�<9�f^����(��)�>G� ,�t��ѓ�us�2Ⱦ�S��+TGaBx��U`�(�@in'�{׻�Ez�b��A�#�M�%��/ZMjDV���ǁ*T�Z� BJ�9%�ݞ'�G�ad ���}N~�j�,?_I��T!�h�u��'��5�e�>�2֏�{����#��$J���B�=9�uc<�y?23V��Qٔ�Am�y J���,ŤS'����B�.`�!�׽IG㫡l�����ȇ��hɋ�#��L���¨ѐ�{/�Q��U�S�j;�����
'��R���������vM�ɗe����^�U��b��"Ppj)4"	�yB�����!�G�yr��3?���n�i�\�$U������;���8�w��v�?�T��r�'�}�ea��6z����b�z������r�(����Ʊƴ�ӂ���j�]�E�ur('����K�ND�z1���q�P]��snU�c���~�D���c�p�%[��
��sC{#��%�.��>Z���A��Tv����fX}��d�-�r�H�t�*JN�BǞ����Z�n�n����-��0"�o��E�PVtCl �A�������!����E9���-��ux6����aΛ��="˱�aPF+�0�(�4�Q3�H)�`��R��=�l��E���sX��m#J4"t,b� �	_ǭ�G3X���
 �V��)�H�1b���g(G��u`bp3U���É��}��C�9����Y'��>ϕU���^�;�؞[w¤M=��M�2�zw���\�@�l��ȹCt�`OV�(6u"���5O)��8ס�2*�<z�;^z�3�)&�]c��@�o��o��b��ENЙ3j'�j_{]��
�5��q�
�A��@ݠ�`Tu��1�;��L��g��C���D�GO$��Q>��vK��/^4G^�a�3-t����{�]K�� ���u�tA���O�6��Y�2>C(}Ak�m 7P'ȲX�{]@T��.'�[4�����̎�]��U=�GE�X3�[c8� �w���	�sK��s�P�^�F���;lV	�i{F.�K�[Ѹ3I���vvhx���l�ehiP�Zlt���G�o�X�d3����6P���A�ѣh�l�������`��//�P��D/Wb��I#7��m��u�Q�8A#��|�c�L���1����;��/j�0o�+���)�����|�AP�$ƿ.`e'�]d��`��E����N�)0�N����G�kc���-f�V���6g�� ��!
�j��co�:2_�Q�'.�|b�!"#:�mI�%�(�Q�}�o[�'ӹ<[L��jI��B���2��?;-\VurJs���;O�B����U����fY��{ħ�t
��3�#S3nh�t�|h�
q?r:_�~F����Zv��LU����Bϼn���C�=���ƝR���#�����+My��5>'΁�)�#R��3��k�^��'kY3���u�)/��
�܉(�X��;{�ɶ��m��(˂�,�Z!��bw��/W��e"��3�c�ݎ��r�����@���;>lZm��A��� �~�T�?$��Fٜs�w�v�ns�{:f�'�GF���(�E��1�9���>����I���f�IFU�$���((*�WP����w4(��0���l��B���8�܉Bo����q̥�Wl����yq�n,]~s;�sˌ��l��f�΃L��;���3��g�1D�CW8gT��I�/�F_R�?�<��~E���m\��UD�/%��&f�:�o�q'�6�� b>#�*_w���vg&���?"��7Г(���)���ǣ
9qdn�P��w_��0��ş�N٫�Έ���s�&�q��`�8:���f���s�i�i� S[������m�D#}ـ���,�P7�T��
��E딒s} L���N�QR���q���4��=������	����I�f�!�w���*��ED�t�S>Q��Wmv���b/�c\�6�3:Qje�n ���jƜKF}��=��0������C��:�[Co��a�#H��]_���h������%6�A��@��E٬�,��k�A�T7��6� F��İ@���X8�%��sDO�l@�73@PU�kSH3X���ZE�K��s�5;�S�� �VvBI��`���ts3-/D>�����=��X6�r����i1E�C%��G��qwo�;D�=��M���Ӑ�@�B
���������ܔ����W�����r�a\�uν�;����Տ\�-���9�KQ���D����`D��}�T�NF�&�r���$'��dF�a�ZԸ�}78X�BG�HU��'&��P\'��䓓EJ��b������5���e�>�|�`�06�p�,R��8c�t���H�&yn5�J(���A�6�Ċ��8��ts��,R�W�i�t�*�3Й�}�p��3�p��#�r�NU�;���p����E �,���	�V�ɀ ��-��Գ�������[[Q��. .���[��s�I}�'��!����㬏����ry)B���y�7��7F=́�Pv���o�Na��N���B⻗c)8k����S��-κ}5���oH9r��$pn�-�6eY��u��2 l#�I�,����Ñ�(9U�*�����T�8ˊ��[,8�dy��c�n�+G�oB��K� {��dnQv�����^���^�;���ѣ�?N��".ಀ�Z^�#D"��U1D�C����_�������չ¥wE����K�Y�g�F�7(�z�9��T���ڑp��A4���ܻE:ꟛ�9*���^�Y�Q�@:�&��(�Č�uW['����bѢ�D٤����-RB�P�ec�"��F���D�;	Ԯ<��n��o�q�xN��i�?/]�H�JG�x�^�JΏ�GG��g�5!�ѻ�#���.�@�4%Y��ᡝ.�qYܙ�;ڎP�q���]Nh��Gbb�7ϛ���X�1)%D�����F�{�A�B��
mV�ޛ)�bP?�x�y��z~�r:;����ఇ�����9��o9��CP��Š�NjU����zءk5ϔN�N������I��91��@�w�=96�ԣF��,d��+H�,pc�ͳ4t���es hx�tA�v~H���}��o� %�o+D#/hp/���?�}E�y2%��8dcJ�p`�;A��j��~3f������;����#�sO0~��t@�G������g��Xȶ�)߷��]����+�bdEkB�F#p`E��H\	�s��P�����fnQh<z�؀��)�,�=p HrwMn+����,�A����Y�!
�s��(<)#�d\�00�R�� "r���	1j@��;�NםĂhǴ��B��Vɬ(k�#�n؉��0�@CXZ �6���)w�X�w!K�.����_4N�8����
��p������P�kz"�	_
6����3Nft�HGۤ��^��c��^� ��ޯ��yt8G��v��$g�N{�*�%��2�)Nxޛ�ZP�*��NtO��^�Q��ԡ��y���D6b�{�Fyx@=�@�SI�=�_jd���F������@t�z��)l9���'Ο��EpH��n:=f��3�-4��M�T� ������"=;������d�o�Da��'FA�CdF!��:`k6�k X����_�I��Q��n,�ЮoѯO 4s��xn���r.��Y+h�x5B����&�s�5ȸ7�v٪cy��͜=�/#����z� W����|�^��	���<A��b0C���h����1=�\ׄ�y5�� ���`t�:5�O b{�D�&G-
)B'G;a!q4!T���
h�iX��k{���tV��{��$��\�xF�7va��+t��Z�ڤQ}�8U�IG*-S�j���y=��-b�id��%�b}s��XW.2�E�3W��s���$�PBF�U��SC��}�0���	�-FD1$qj+T�)9�=
�
A+��*tWh�>������
����VW��N�fA�z�C9O���]p���e���|�fԧ����tgT���9���;M���<(N�G�55	��
��]-�Ĉ^�&1�)EL�Dњڷ�l�Wo��HS*(KO�yt��ڝ��wH���<�Q��&'�z+�&>)�ߟ�#���ǽϛ���(�w#M�@.s4Gؓ������py|��z���l� RP������k!
8�rPq����RS�s �U�
��hJ����j}��?���*Z�W�.�O��o�.O߷>}�(׏�킢�	d]���@OڄP����s�ݠ�r���<G�V������g��2�q B)%����{>�q|�[ͯL8s��Ul�<�4�À���yiFO��D�q�}��Du��f���"A����r�n��H�[���fs��@!Ik� 44t]mp�Ѣ��u�]�MȨ����!�<&e*�z>��i����P�4"р�vxʹ�,���I�aMF[K��;���P��E���W�w�����,��<#R�VPF$������1ʾ�
�T���ۄP�t��07���DԻ�2M��=e��]��5A�������C�"
[ZD<�o�_Nk:��z
�^�ItP�N�a�lvH�>뽓5�Z�t��K��:�x��p�:�Ml�촻(Ӳ����cG:�lq����>)T���Z�M/��8h2��b]4�^g=��2�~[4O�+|Џ�1N:���m��D�����P�޻��/j]tvcT]+���9I"���VR����Q��y��'�����z���F���9�j�5��DG���r~�������J�������
п�v������/���|���#Oo>�O��{��\��1]ߞt{���!?o��ʽ����	e����JC;A}��d3��l���1'�߇[����`H�,o{�Ȁ��������.7��mD�?MCvR9|�Ip#�D�uD
t!�"4)7$��B�S,Άf=�Pꝵx��3��#?���ל��.�:��P.<��g����x�#SᏑM�$@��F�*c����pnsf"6�X�P(����!.{��e�t�7�XC~f��x)Z�����M��Em�n�X�9E=��n[��@��&���J�����1ǟ��,Pm&�����
*}@���-p����9��v�������[���_FE�+�À�]����g�d3�:)�"���y��^#����0�Z�Z3���\R1��d.�j�E߼�4�ra)�����o��^b����9���wA�|����Y�3}<��=s�ߥ�i��DRc�)z�U�I����M
�U(���RO�`׷����_h���'P�`��?�����^���?�]�K�~��#���~Z#|�aŶ��?�_�[��7��������^�>���?��$_���p��(g[t�JW-:dT�igz�j��P-?`�K\s:D:%J�~�� @s�Y�=	�,x���=��.%��Z|!��Z:@شwʪ��4os��qx}	��!�b9�%��Ӂ����pbn!�o�5kj��2�PU�����\�^kb�1$����J�2?���
w��� e����	�D�����JQPͰ����/��>9�QB��?�������qRV��m�''���K�3�{_��!w1��>vM,:�8:	��w.�`f�zZ���(�1'�@��߼����%|���i7�V
��l�:�/�>^3��<H���w�}����uaAAcڳdb0N��HT!N�j�����y���T�r��ۿD������3R]����P��	�vW�����t�}��x��HV��4�-��<G���B�dQ<��� C�T�ڌ���O�zF==��G�ԟ�֪��
c9�!T�i������_�����<~�Ͼz�����?����+��?���կ�4������K?�7��ͯ}ܶ�����ۼ<�~��ў>�q}��UY���+�zV=�v���#y��R۫�{%uFRb�.S|qPǩ���L�(���R�7x'EGo\�3��Ľ',)^��A�4������?��0#����'�><ę�j {��k�ZYJ�yTmK8G����#��_R�dO�s.ܓ��>v�vݝyE�&A�؝�a�͞�DCJ9�9� !B�ځցnSkuR�N�6�e�������g4�w*�1��:���s��FP�mP0��1B�?o��I�I_P�Ӗ�$t/�p���<�����;��);�r�ɀ�:	���>rYC��wN�S�0���d@���,C/��;�=䥵8f���N���������X*�3��QWq*b���hR"����r� U(�	�t�����g�j��7r��h3l�Nr�c�rf�ˆt�uLR�i�{�R��a�u�_��O2���	�d�p�5���Ƙ���h=2L����IQ���R�����$�QR
e��c��T�����>���_����/�?�����?���|�+);7����#� �ſ�����_�����O��/����^�w[9���>����+X	�W���b5̉5����������z#�7��~􂻇˪�GE��D�����1��~��vH�ה����<�^��=�r�w�E�!��$�
t��	K��N4"t�KAQ/|ӽl�!Mo_=R�� ��qs:�PC�h�fg�%�~�8���N��1H��r�y	3�-�ށ�['�ݢJ�A�*�l�h�!@CF��Sňt�q�7�g��
���& ��4�����������'�3�^����2��=�]�m�IRd�S�V<\|N�`ϑa�aIMݟ3��mSq�F���#��_��:ݿ�[߿�������Y�����[f���t��QjEe���8�1��
F����vl���z:�>,(�RC�qJ�L9��{�1�#苑
Ǻ1����9�#�	�߳=G�!��|G��K{�x���Π���.RǄPN�G����z6�}yQM?��68��I��� ?���ß{x��\�����?����s?�����!P|� _/��z�����	|�w��_���+�o�r+��=���w^��+t�@H�	mӺ!*��<mB��#��iCW5�[tp/��ţUo���A2��������U�����=?z�zI�T����9�Y�~�D=BG@�{2�8����k��c�D1��#:�< 7��6�x��X;}�1�P���L�]Q�x����`lL������v�ݻX5/x�hV��a�l��vJD��T� >�G�cIk�h��O�R <ߋ��d/Ϸr��}q�������^2F�Z�k�6�m��H�v>���=�4VJ���HE���b�tPPa��7�oQCA��Hόvɻ�à�\D�<>�Z��c�{����0��ϰ����;�\����E��pH���-�T|0P�`��������"��(��z�R�sJ��C���Ngи�X��71��ɩ��O�+��h�=Y���Vd�&��S����X��;��Y��H�I�(�lQ���=����јhSV���a=?��W����?��_����ӫ������F|�t�t�h�?�=?Uŵ5|���6�����>���~G�X�w���կĶ�d�C�LΛ�����:S٪� ����*�A׌����#�q[ݗr�A�q��T�z�."�D��������g{љ�`%77�! ��g*��@M�N1a2V.2o�ݴ��ˉD��p�V�V�A�d;A�nS�`����!��Z�_O{�y��c^j^�DFQ�H���2W7\�w�</����I����&m]�6��AA�^͂�;�TLn5�$�S! ��1�jjSqGGG�����ar�g��m�F%���D�><7+�w$��#���9
��@�wV�6�]@�ԛU�������耘�,�ؔ@�Iǉlx�*l���a�����(��{���ؚ4���iy)ʞ��^>���P�{	���QkHf�[�>.ڊt��Jݜ���Ή����h� ��S=���H�`3$���J�6�E ���U!?,#�iݰ�!ϒN�4��f�?κ�^ڎ���{~�^�A����(�?�t<�!r�g��R� m�Z�^�zBYΞ)٩Hb�D�E��@B����������|��_�G��~�7�r}�^��}�/��~���M|��}<��gN�����imu�=�#��U�\�a0*l�}�T���!��G�0Ըɡ���xV����S�%����g�i���}�����͓��&6���!�=�Y�� ���FPAǆ�q(��S4�����+� mP���Qu���tX�H@���M�S��^�/�qWF�T��k�6ѯ�.F��;;6���#�04��fp)˾�ɨ���)�|��� ]��"�ֽ`�L
铧̓gޢ?tLY$Uk%��*@&�R����U3P��$^�T¡�z�D�w��"	�EgErV��x��;�{oc�-��c�Pp_�r�A@��>nq�� �'C�O�r��6�3�f �d["I�:l����P���m��MD7G��r�sQ�X�{2zgÑ�P��Nʔ�E���\_�\o�z�A2�"h�H�1�Z@�T���t����`ش̲�.g+]�j�iT�q�Q �BNe�����6��Q?�U�F6�w�o6&�����nF/&�7������I��j2":�Bs$��#C�d���*�:�Ƞ��drp�����M�^���(�>�X��>>sy�3�S���4z�S��s?��O�N���������x��=��c�W��~����O���\��W���r�����y�j������
�
mH�ԃ3zuJ��F���3���guzg ��}��~^͕�Tޥ�0�;>Q�z"��X���z�ҧL�� ��3΂,��{��� ��I��	�n�P��5�<N�r��i�������Jґ[rJ�=Vrxw��dx.{�~�y?y��c�^��έ_�R�������hTk'gDa\!��;=�˳�Agi�K^�;d�Nt��h�`��뽧LmNw+�����)g��Ϯ�5 Z��Q��S�;�4�F���Ƶ���]^�������V�Qйo���:�����c�%Ekf8���:0�Z��UQj�
�@�@��6���v���zGa��m��X+T�M^�3;�KIG���ڼ��b�^Xs�ĬD�ǹدW~���@��ⵌ=$/��;!�x�ՑU��F�b]I��Ǜ�Z�r��j���>l�-2G�������3��������}"����o�������2�-�x|ϯ�!|��� ������WUdٸ�����#6Q��bסh}��	�ä\@� j4��͌�X�{0����ctH�����f�Q����i�C�@�(�N0��_��"t=ٷ�����;�����KE�� uQi,P#��37��(��n�tB(�Nc�q����a�윪���)O���Sۣ����@X�U������
��XUU��)�9�V�*���v ���1a�����r��1R���	��c6�#�^4�p}�Kk�N�Df���zWE��[��JD`�AHs�QM|�ji�@��@�����%'�@�cO4O�y�x��������I��M��ұ��]4�b�,�H>\J�_b�;--'�DQ����k  {�IDAT8�)�R�S#��Cl�+��ST���/��h�q�bOj����9ǥ�Ss�z"�'�4ޕϹ���7` �w4���8G�8�� �re;W�bRr&f�*��F/vV����N��<6������?�����k������mt�r�_��?@߮_xx�ST7��V�'��p䛍9Ǽ��R�%�bԆ��)⽩]�Ź�i_��z��W\�{���qϻ���a=K��6����@�"7:���1�wy�c�v�#���&�3��Wv�u/�Q�wQt	%�)���ب�B�J��ή}�qǺL`��JhΔv�&ϯ��cjRBw��U�*��x
%j(L2ܥ�<�Maμ_���@Wc ��0h2�S"�I�Q�%t/זb�t�EI�@��|qW��䱘c��ˆ9�mޓ����	�4t�
��$�ĊW���%�G�~��ü�H�O���/�GBn0^�,��|�
H��L�R��^�� r��·w=���_��@�	����G'��='�G.(������|P�U�;�S��hC���lNz��/�����ebv2�{Mg����%�ِ�8�i����^�(�=ݞ�@����J�U��4lV\H�-�DF�����j������������|u�����
������xz|�p��t�~͏�ķ$����6��/���/�g?�����&��j�簾)��,���
���c���b��4�0�+ȩ?4�Jx`��|w���<F�d���� �[{4u��߇�C�d;4q��q7帱�*Niy�yVA����ޕlֽ ],Ci̠3�AL���o����ۜԢ:_����d�W��*�{51[E�k���H�n%�J8~�
��ٽ�euF-���;<�SC�<�C���f7�6'R%�,|�k0.�r�i����������;<�q���A��=��\H�U���p��D���I��=:'���b��Ɂ����V�E��`C����隍�|��*����,�Ѱ�2F��ɽ����l��B�ڣE�@(5�A�Xo�9U�K1�7��Ҭ�X��f�
pq�ݲ��s�{Z{t���<�[��T~+Ծ���:�*��)z��0�]��<�G0���L����cׇ��	�щD�R*J9���@��zYD9�����[ey���������g������5����: h|ק��?�������"�A~�n0���
1:��; �������ӌ��Zl�o摂�{��+na������`�o�1U;�Ӝ���=e/Գj���A7�(#�.^d����o��
�(^�G> ]�Ό�f�}b�QL#��.0x�&�tvL�6�ca�U��W������{J�4��R�U":1�k�쎟&��8�e�͊����[�N�] ���3i9���F�` ;�y�q�#"�=�̕D��f85��ǘ�(���Qr�q�*J%&�IՊ�^|L��=�3�אq�7�ywgX�����p�a�c�8���E�����7f����,�WW����[9�/�ɼ{Q�;�;cp���D�y{�:�f����ާ*��]�Jo��r#V�JN�$-)[}��5а���IF�]�e܋��2q�8GGv��;�:˰��n�MQ����$"�`�0�׎.�;��ہDEJT��#���c�ƭOlF��+�<������?����/������2���;6���_���ÿ��g�y����/����/��� ��[���n���;�
)S���O�WOաMσ���S�ӵ$�o�ncX|
>�[�v����4���k�홆3��}�0�&�ɫ���A��D�M�)G�&��� � �^R6#���͍	[4�<r�0c� ���R�ESTu@�3����r[�*�m�@̎��E�J����/� ���{��S5�
�ym��z�X7�eSl�8�Elڔ�s�>�`�t�P��Lh
d�vvx��1�]~g������(��HQ�v'�H��{zN�Z3�9���c'�N�t+�$o�;����[b��YC�l
]!w|�o���Ao����Qp_OS�_P9�5's������*�'�5
̣�h�+�!�8�����hZ�:����#��Uw`C�H����츼q)�,�H�:���,�Z�@�	���������"ք�����HA�� ��i��ApG6��ɩO1p���/a�o���>��|�����F�μ�=:�����~�ٿF�0� �G�LՌy�Pf(��� �������x9�������������oů��t ���u��O�5�3�������|��������i�=]�������w�^�X+B����"om3�늫#��ywod��n����6�n>襛�`�1db��,U�}��w;�<[#x(�P�0�,������Z�`!RXn��qH|`��7��1����y�~������aW�E*��
M�k��(����S�,��o
��U} ��}�<�x�PW������]Ѥ�ڀ��X�b�ag��9ڔ����V�nF*����g%�:9�Fu,�L�0�2�~�4)�5�Cs��(��i�]i�<b�| ��UG@ҽ���p����;��m��~~U�����BLA�������X��n������	Zރ�����,}�M9|�������򏜴)�a��m���Q�����WdUQ/3�C��ԋ��za����R@��h�B)F�-�љ|��*qw��9��V]L�ȟ���%Qk�"�E�a��aTp�!}N� L;YO��|sDC�C2h��ٹGd��=��I�x"�ʌk��Ȁ�i�*o���T�����&tdgj������\�d�I�sDK�
*g���W����㯽y�������S?��ߚ޻��t ����I���/��_��^_}��U�~�_�����~-�3( @�%��P�[�3d�=g�\��3
�o�������s��O,��zs�[O	��{��0�?
����P��#<� 3�1(��p�`���I��X�&O���,D6Ioҝ��P�}�G��1m�]�
fk$�N��v��0��\��
q�|#�V��Q���5!Wx2�k��L9l,YQk���l�"�BCfW���5vG-��l�Ս(ᥢ���A��Ĩ@]�rXP0s�W������Bچ�6������98�Ű��M��DS�v��d|���U¹p4ϨO]n��6G/<SzG�4��	�6n�!��3��.X��9�r��y��9�Jٙ���s�����_�d�����LPf�m�n��$�N�n=r'���L�i�;�2�,�����PD�/�^�og������g}.�-��D�3u/�6 ��\�_�������8p��r�B8��s
4	�KB�\�����@��BkW|�=~%�_�A�����i�>>�z�~���ڷ�E*�hW�r|�C�p�[�l-]�S�4ra�M��%�� �����_��ѻ�'ŋJ��1G���hg2��pX�]�4a�-:+����d�[S���ם��G.6�;����fo�b��x�*�l4�4w|F N���1Q�qM#g�{Cv�i�9uq#u�a���Ju���s� �֦�4�&�8-+[�%MF�����9�4���`�{�d3���c�(����>�W�v��9��c��hh�d&��7��"5!IC��K&�Q�x��{�����WH_}���]�Ќ�(y$b͐g���
��Օ|����2Ҍv� ��?���O�i���|)Ĳs��u����ñ�~alw�{�|^8uq��z�y�u�̗��N4e�32(�w�sv]Y��������dp{q��T�Ӻ�3�)����n�C١g��s}  L�䨲�C���c��=��j=�=����3W���r�����hCگ��5i%O��,B�ji�@/�<UPY@��%�ğ�������?��}������Wl�����	�����u�ׇ?V��GD�?�}��RVXn�X����
g�S��@�����2�\a�1HV�1�b2�����f8e�!_��'/�F��3�/�r�����0�{��q�C:���+��tj�ϝ�$�1�{��V|r�PA��K�{���s-w��M��)��v(T��鵻H��7 �{�A\3���W1�T<�#�hB�n��*X{8#�7�7 p�0R�ժ��͝5F���Z��6�@La�$����|�Sq20z�w
K��x��/&��[B��Q0����:����E�w���A�
��q��������<:K�;hθ �������':���n�#�Y��Ζ�I����$RK������
=����qxtȧ�o���N�6!u4Г�+�>�<.x_�0���*�Y�>S�:�SD�:r� �3��u\�/F��pz�d�k\�����B �(�0���V�N㭺S�g��wQ񌀌b9�qu�`���X*��<��l�K)V��S(_jI>:/A�GC}SH���L�1�l��r�3���d�{��4q=e1����zz�7���w���*n+���ǯ�A����o�~��տ���U�?ޅ~-�P"��&�/hޝ�r������&43V4��!�՝�=�$�6yn���/F(�{��7��S�������!�IHTSk4�;���t}@v�?�Z`2�Sn��L���W�P��8Eͨ����ɘ'�8�k0I������&�0b����o����Ús�1�Ȯ�5+��lk�h�6�"�+�� K:�F���x�G�~�UCl;u&I����k�0)���0\�p ����0���㛭P����E�� +{��ۮ^���.9=�&�m6��2-|߅r9L$��fA��ơP T�T����؛���4�Y�u�L�q*�B8��i�fu����M L�_�C���ʜk�`,3���X��k���
P27-6��{����H^�y�F�Z�bC����v���G,���+1���{6DT\�u��=C[�st8���r�3Z
	�N.���ʭ�����M������K�D;��{/��C>]�a�r�	J6�	��i�+�h9	��_ZN��'*�&賟ů��Wՠ�����.�-��C�����(~����R�ђ��&��w̥���/���z�ɽ�c$"�㩴�@2�x���杇IJ<.9`�Y�)'�vR��0��#
�C$ޮ�0r�$�D-��3�N,b�U�H{4~�O�"�%�n4��Eq�\�q��~U��ppr�o}��aBe��?����؋+����(������ڰ�-&V��r1Gd)x��qk�W�ϝ���$�]��m�������}d��es}����!�{e�;9
���'��f�U���]G���b�c*�$=2��>�H��n�
�hv5ǈ�#^r�tΜ�J6�$`q�������~��ŴV��LeZ*����ϔ��\��>g�u������~�F��n��A� ˺T:zQHS�1�ǝʜe��<U`yx���3tk�ۆm���,��U]�D�&�B$�Hh�Y6�Ο�p�����0���a����i'>:㳃�x_d�_�{�{�a�{��Q}��x�?�ʲ���.��A/���߹���?\N�oן����oů��Wݠ���������Y��]P�$��D�?g�1M�a���8հ�.��{���J�lƬǴ��]KD�M�"��#e�	��1M�{����&%�Gh��w���(�1}���# .3�6��&s)Ōs�9݅&�k�H����gT�֬&DV.��.�E:-hq�B��P����Ǵ�4��k2T����fx=����鸏��4gu�$��m?} �	P�S�^g���	�W@�2�
+����=#�
����yDP�R
ά`w�p�3�	�GdtB��l�D���\���A���1�>R���ϕ:�jr��̋&�к4wX:������tt:�8���D�u��FDsxJ���ȏ��N�i`ҹ���D3�����!ս1pٍ�m��@���J�o �N1j-�`k���H=΃�cbdt�E�O7d=}L�����e2�2�"JE}�^�`���a]W�m��A���;�j�iL�.���6��C��G�2��LE�CC����ռM�t�3ՙ�{s�s����`�p̵N�3~T4�h����X��\+J=��
.%i����s� ��-���x�������~ ��R~��_u� �����������k��_����?�x�qR��k��Gi�*�2/�Dl�='�f��ȹ�\9kU
���{��vo66/<�1�2({
i��̚q�S&��( �)�3 ��Ǜ��W4 �h��52R��iE*��V�,��x�|����v�*CdC#�(^�U�bɫ�TT<�{��%��3m|��Ӄ|�Bw�aIX."]�[��k��R�F�!9U��*[YA��nX�׉!ڰu`�*��@��nO�������(�8~�Lv����פ�8-��2�Hh�ް@_�p�$��#X���L���hҊ���{��:��3�RW�:�^=K �v�`m�.��P�(*0s� 2N�
��6�� ���ZI ���/ � ��3P�"͇	�!DP-���Kq�:E��@]�~�#�:���Oy�TA8{���ADܐ�jB�����������9l�AM����m-�샙l��2N,�4�|ƹT@�*ضo`�Zh�X�:d�D���r��a���t��1|�����";*?f�a���49y�m��&v�Y&�<��0�k�0�i\��/o5 ��h�>Ӝ�*g�ogCP�,8�k���Љ�"P��]���������~��X: ����C���_�y�c�友�E;��唹F��� e��q1���DKC� �Vc�#~�a���|���O_E�FD��VJ�N��d�%Z��]W)�B?�4X�|��G�Qe�H����[F^Z::8�EYD�u�C�ڰ�����xd1R9�a�#q��Zs싺�{Qّ��P
7�.p�3�#k���X�>9zc���`��Fh�]���J�B|r.uW�$t�*������XQ����<H~Vb���
�m���;B�{��X����n�ۺO����A����ށ��n��)v w�B�
�qD���O��2�)1�����y�d�����`�(��4u��[.�-{�����{��i���	Q��A΢���>�&�;�x]�� -Y ��y�Ul��9�x
ʉp~�@ߜ �P"�z�Њ�4gtv�ޱ^�^ϗd�d,�ps�����)9����mi6DՈ�DB�vw�x�:`�ӵ���A��NS*��I��T��՟g����W��|�������[}�c3���G�o~[oW>=�;��O�<��.`�@ڲb��\\�,�I1
T
bXTl^���{�I��}�}�j�W<\�	uŉ>4+M��<�'�NcL�����[�����Üǁ	UESͶg��t�ϡ֘�dF����}F�k۰��E,LL���$�{��"��%z�^���zג�R��,��w���7�7F�7Ի#(��fQP�CiT��]
Val=R4
5u�ϙ��nl>%pF\c�S�hI�����A,5��&Y�:�w����g4�_rA���&��)c#
(j���~B�BnU �'}��+h�5�ϛ�C�=�h����8�2v[62a��됋H��C7�dv��|�;������t��}D�"á�b7�m�cFa�h�ʔ
`z����j�2��V=�T���S��a���l&K1��A�ay� }�F�$�e���
�*�&��l�~�!/K��3�я"w��J�o��_H@�df�AȊ8M'�H�x��dDȔ����`^��Xu;U�؋s>?QY��e9��'�y=��[�����͠������[���|��_��?����h򛣚�,�H&�y|�8�������mT9{!���a�^z����5�>
M�OR��ÃӃڑ0�4$� ��wJ�	���!��5����hD��������n�& !�ްiCG�
�P��h�
P�y@����[z쭝+@�e������N���~��P*�A�ɫ�cm�`E�5�����4��	:�D4��{�<�%���C�����m��@��;>���V|(�a����A{eA�3�'�'�L�b"r���ioZ�����!�{�F��i��qo�-}���_/����� l�p�>.�f�,mAP$q܍�X@.�RЉ�!�)b��О}��m���8lf%��sFn+F@�H��j{8ڨy�(�L1����pPF��B�` zoh���0�8���[CW-'�v�b��+zP��|^�u��8[qQ{�>,�;�������!�����R#����SR:Dn�sd�dx�z'ӝ�|9� "�2p��?�/��G�\O����p�ys��'����[�/�D���_y̻���x>�}�����|�+�+Z���B L�ژUt��L�����OPr�.�|�DD��c6�s�����D��y�!�Js.*%���V�^\6yʉ���3v/Sqe�0Y�Td-�/����sLe�v�N6{%:�����������=��ð�2��:�Oާ�̊0�b2�|�~?����1c�P��l]�|��(����1��i��S��O5;��Q��t��r�n8#��2��fx��9����-u/Y�]�����Um���~ؕ|�l�$1��C�Y	��nn��}�jv��\/���6��G�
ι�|���v�����ɨz?�,v5���-�߀9'>x�<�Ǿ�\�Y>��ǽ����f��^������3Mn8#_?��TQ,@�(ݣ\G���G!͌��	��n��;�Q����'uQl��m�W�$�(��Tf��<NAԋ��^�i �K^i����`6��{�(�& ��YS̓O�@*���{�x
�E&Ƽ, -P��ǝ��ᖿS��������o������oK���?v�N����i\���v~x�����.��$Ҡ�-g�N!�YU��b�ȹ�(�k�����!�����t��A�ȫ��j��T1���A�|`:�r����3^E�k���.����95#�(��n����Ѐ�=�ǀ��4/�i@o�l��t3Ӥ��+��PeT����Z���En�q�V��,�^5�mJW��������v9�a�
��veFA�O�o/�u[ �ص��W�(�Xv�R���N]�n��V�DL(T�(J`�1��=m�\X�S�^x����*���eT��
j�6�C�(h���u�O���Y�w���Wˡ���[)!��A��¹�1�ƴ���>�=�Z�M�M�֗)!�8;S�|�U�Wh�o9$�gG���丅�G^����"룎�}2��@+�,�
��7HkPQp	G�u�s�
��q�ܮ!	�X*N$t*���7x{�#u����N!�����{<��#'՘6�h@�����h�c��	.��֙�uǣŞK��}ܷ�Ǎ����l޹}���R߂�O=��}��	[�~[r��<�����#?U�?�����l�[A�G՛��Y��A@L��,֩Vй@�8k
AVC�Lw�N�&{�b��ｲ���D���}z���y��!ǎ�v�lv �Хa��U�F��Ū��U���A#���A��|bu~o"g5�@EA�>w36_}@��f4��K
��`�e84�:�Z_��G��'PTG@��%VQ`mT�O�v�(�4��U�u�7��u$7h0.t�&7���\��O�/���o���{��l��B�ʊ�4ǅ�>X��^N�I�$"��HC$R/�SD�ٹl��G����������k��bmˮ��9��{�s�[-�"�H�D�UC�ɆaAz�yȋ���!yH� ���(q�8�b;Aذ��U9��P��I�H�b'���朽ךs�<�1�Z��[
`K��<>�X��=g��ךk���#yj��$�$�@�:���z�A�·�ȑ�B�y�E{�k�ܷ%OpB�m@�w�.��F�o���p�V���3���	�պ��F�ͯO��٢k���S��v5f򜮨~>$g[#0����� $���D�}A���A���A>g�{���1VD�{~�x͊=�{�����܈b�8h=B����o�C�U`۬o_�~-����jΞ[�]o��X�y+����ސR�hO^���������`\���ɔ�8�Q�)�;��	H�o����{�ӧ�o��]���|St ��7����3 �oӜ�
R��H�(�S��Y�蕚�b� � ��T�+G�d�z�����=���V��z������jk�ppxԶ�0�ȫo��G��Ͻ������w@e�,3N����$�W�A�c��X���z��+��
ؼy�H��!�[En;&ɦ@��gߝ׼��X���#$�֚���RoTo# �@�R����t�����r���㄄Rp�ͨ�!�����w}u�n��:+�C9`H��f�k3C ��isŔ*v%!�l&��6�m���ka;4®`�yd]�����i��{����f5�lMW�Yĵ��lb�$�*6^9ۺ;)�xBZ���Pb2�%���#]��=���"���z�a�x{ UF��q��+t}���ovK���%qփ��f�0��QN�V���f*�O��x�{m���	�#�� ���
���~�����Gћ��=�f�(�h��RF��(�6^C�" mH�.*eE��K�ǹ�:^�E�y�<�=�/�ނ�̣R^�У�ϟE*]gk��)�g��j��P�:�ڈ�wAu���̄�9�~�j��kZ�,h�lmg�3BU�{��Ϙ=gkQD�He�i�\~���'�����w>�g�}��i���>�/��G@��w���P����.���z�S��Y����u=�H6�ΊX�0�vV\u�}����<?�e�w6^� �J�uz�6�z3\�Tp�`�����-3
���e[DK���n،��o0�/t��c,vX�C-؜-����0�����*�9��}ޣ!�P�t���(��F8�-�ko_�ń#���s]�k(UsS����r�ن��D��K]���_��[r�(9��q���ѥD�P����F�i�;z���|�*X[nVw{=�5Jg�~nܗǴP����9��nc+.,#>$��Q��d�&���0[�^��0�.����Z���z{�z$B7+���{?��}��v�z�o<�}�=FNx�����e�_���>�U�~v=��Y�Y��X��u��ݼ����
²4�f������V�Zdu�d�9��mޢ��kŸ*ԣ}ԍ醡O��̍��j��k@�w�U���ԪEs�߭׼?����w��FPO�l?��_�fx�{�������Y��\���v?��5���r�4��i`�sB�T���rE\����3��^A�w�,�i: ��=«_�,T��'�?)ҾhO[Q�چ,��7��g�<E�Y��U��C]�4vcn���l-��}}�R������(W�X�]��������;�y�ɍ|��y�U�4,*�;���O[�<���������V=��&���Ekn^-���H�ҲjcCoN���_,��ݾ0ڒ t�|D4ܪ�n�9v/�z���Y%�����Bk����o���I�T��T��^������HDP&h�=8B�q���=�%+JR��:�=i�д�Z�u}���Sg:c���\�՛ܬS=�����ޓ�C��{Y��Mz���6�³]裙�7_�����ڸXxT�,"▛�3?�ܘ	�@��Wj���q����^�g�7���5�H��;7��Y��lk_n@m�W�V�st���[��lv�8X�c�B�E� eF{M�JFJӴ�߿��m��*���<f,}~b�״{���o����.(�'���c�����v�G~�����V#���Z+�#\]5o�Lv�����o�O�<����Fa�����ϕ�U������a�y�C�'��G��l��c���x�\�8.)��!�ݟ���r�Dx����7�o� ��Kb�)�ť��B�M���KJ��b�m]25 ���=n��ᦛ<2%h�X;7�{����z�ga��p�ж2`�������g���o'M�}�\a���ϓV}O�uS%W�S�!�	��u�3?[�*
ۃ��{*`�OC4�_y����Ln�Kkr��Mα�m�Ms	SHm��,Xj���ൄ&��ӱ��0"��X�p=/ :��t�ߡ�5�	#wj��ke�v}�C���A���{c} �����%�b��}z�iW]\0����#x>���8YΝ�W����_�
uc̨�H��R�Y��RJ�G�W�
�q���n��|^-���5���Y-C_���nK����@��F�˳N�B�aw��~�i9a96��K���r��M�K��!�P�I̦��Ƙ"/2�բ-�V��Ix����MM�#������~zc♉��h��������g��r�#�����CΞ�.=@�3M����<LV߰F����)�a�t�"m�P.P.@��\�Ly��D�"��/~�L���s�~/���W..���|/(�����]��f�Y=���*��@#�8���	�=�)��B}�w���r�k�n|��}@ȣ}���gS�zhY�Ko66�����7ӋlN�{�je���N�Q��g>ސ/d5˔i��>�9<��_�{M�����u���h���m��!H���������W&_)J���$����1�<mk�r�f�������6,�۠ɼI"/ SZ7]d��Z?pv��3	_�{V7#���k��L]o�Y��_�.Ȅ��EX7G����K��u-'P��z�^�LxUIܖH�z�����t���=�n����m�����=�k����'^�@���0�G��|�v����������	*e�[�����E���H���њ��\��׼������X�_	�d��"�Z+겠-ER����,�ݣtM\�P��2_��l"�g_�\�>��Pd�c"q끎��nu���o���)o�k�M�M��`�������|�l�7j�!YtJ�s�f|vA�Jy�4�/���SϽ�C�����|�t ���_��G�A�����(�zഘ"\J�Ruo|-8�n3�(���77����c�<��^�&\���<~jͷ��Ϛ
�)������f�=yȳ���U]�%lg�w���ga%�l�=mb���j���3dcWW/�7勈��9��=���������3��[�g5:��7�����&�������P\����4����I�&�j��
[�Xl΃E:�0ڼ�-9@M#���X`sK*�0�i�R�z��PzT�_��d�w��7�n
v#�~�V�C���M�ϥ�V�<���C�쇆w$���<c�W[�q}:6�v/"�?�̣m
C��("hU�se���M�E�?���r�����A|�N��ͪ�a\oWjԺ
ed����3d�|6�EE��N�,f�]a������۸
_��kDz����D梣���@��'BK�^�]W�j�ٵy$}#�ؿ��n�i���3}ܬm���&�cݳ���g`Ѝ��Jgn�*�k����f�|m�I/R4�=G�NR��5ev�JY���1󟑺,x�xCt x��n�W��֝�_l�?B���Ԓ}�J�jT=d�'J�����x3e�B��V��|�&��_��^
�}H������i� ������"7s�����p-�9�|{��Z��Y%_J#�:z@�?$��0�����f����>�	�L��>Jz>���B���M��>�_�q�}
��ʞ�2�M��[n�}F^�?��@�!>DVA���6<8Uk�iu��矂{�m��Ms�uH�Zn�y�O�d1O!%7~�`Y��%�A�庯Q� ������#}6A/�qf��C��=��HX�Fī(�y�D���tow�3t���&lFC����Ev4fh���u��ߪ�m�3�?0�זM��Q=��~hml��8������0Z6ѡGX��7���)�G�k��v��+֐��>� N
i3>|t�̋�f9����Sf{����Jƴ+���n�c�įA����z�R��lv'���t8E��&����$o����u��{��u����M�v�e�Wt�@m��9�F��>vw�l����ꐽ#�[��7�Mjek��1�}
�$�dav�l9���ze.����OL��J}C�s�<��r�í8��+m��?���-�Ia���B6�O���ΐ�M��%��@h��5�|�w[�لf�-����X�HCLHc���o������r���s�Y��7� �'����������SF/��;��=�N}������-z��ՠ;*��%��9�6 ����6*N������~h�5���	��W�ԧV��GkU�a�+k�lc��#2� -�tif��x����z���!%F&��8�A03�ZaS�D�B�s6A��@MAd��T�\UܛOk��<�m�t�����J�m*s����2dh��h��6�:�B%{'�goS�T�*ZO>1-C�$s���5�	=F�%������6
�Z�Z)�SF˄�Pջ�� q�skuYX�ad���=q�#�	
~P�z��3b���:[���{;�y2��+Z�F��$���X�Ao��{]�� �vrJ�=�������z�5���x��x<b>�����+�8y�G��� �12��`=�b����5�2j~d�Dg��x��Nz���gz�C�i�fk���b�]������������筱�N������d�̉2ɟ儔
R�����"����o<��|����;Пx����_���~A��~��OQ*,O��U�BR>�F�@�!vb��	D �E���܆47��o���t�����ۙg?5o�0��C�����zcaZ�N�j_��H`ZC�}ZQ����=�&�<f}k���N���ڇ���TLrec���C��/����ԕ˺��zЯy��
^�`���x�����͙�ޅ��U@X@X�z�-�i��it�{���[x��'p���W_�7�/��M%7�T�z��4�HlmhW��hk����GPl�L;��k�m�%�s����d\�����c�;7s�7�)�����:"c=}3fx{=��;�{h*eU�+�k�0u��`�(�'CϿ7bHJ.����5��Eic8Co�Y���q���7��*{��z�;{�d��ߌv��H�l-z��GkЍo�����l3�N�������e�jg.�i���=/��`'3��b��p%QL%Ck#ےim���0��n�9=���y�wQ���=�M%r��O?����
���f��MQܸ�����{���#l���*Z���\0�(����iw�}Ⱦ�O+�ߎ/߿8<����F�� ���| ����g�_TF�K��!�4MUN@+X{
=t�d��zA�`���3o��{�#F�����d=T=�=���F�{l� l�@x�E�CD^#�	麐��&^�m����(���7���rֽ��N�,n��fL(�bX���ׁ�z��9�ǉv�m���u�m;�u��%ll���5������긯��Ud�[�j����iͼ�:�q-�)����	/��9|�ޅ{��z>���0��t̨}^u��~��nMVcbՕ�Ȕ�{�
u�YU���VX�f�?K�=�F�_�q��_������D��&xr�zJ^p�Ѵ9���u���:�!xb�iy���:&�	u�u��:�_�M���2���o���#i��g���腐�P��AX�[���	�m�7֪���0�Q�&��Q��8��pA�i��eF[��lW��g��(��
"Eʄ��F�21���*r����tkA�mRghc �_�GS�ۃp���p�t6��fG����it���/n`f�Ƽi�>nO��ɏ���ޒ�t�b�����wNy���@y��g��O���'��[߃E+�}���z���_~
ZT��A������x�Q�
4�9n��U�wk�&����dV*�-����8��G���x�`�/��w?�W\�eUA�}74ȨF�����t�Y�~5r� �������2�V�V���V5 �
�K��bu�B7�9�<w�#�:��6E�g`h�����	����^=�ؔ����j��^��@85�q!4u�X��	kH�H*�:���{����k���]3ж�-5`C�Z7�2�*�&x���\CQ۬��IHv=�m��-kps�b�_3�'�z�lDf��������g���}s뽒�>�+e�J��{�����R�{�j��ŕ��3*%T�ژ��کG䚎��z|�.����c����a,���9��YMVCDקWim�R��@a�x�W|[��M��B� ��6S�Li1�ͷhc��GJDP]��9L���vhˌ��R�s���Aٞ�B7X����u�G���q�Ekg��fxG��yx�-ճ��f����\����T<t�7�~D�3%8�l�R��3(O�����4���|�o_?�C==���{�F��o�Ї��_�9d0���禩�WJ���w/����n%r�m��H�~���J�����5�C��|�M��������}��S{�����џ_�L=L?���44,RQ��I3Fz�ݦ�<�m���S�=D�����2��k��l������::
6�a��<���ڶ��P�m�Mׇy��4�+�[*���Hl.UQxQW}ځnm�T�cePb$m�m�	��V=|�T|�׿���������H���	=�C˶^z��I��g-X�"&��k�u��]|�&1r1��Z+j]�JM���ȑ�����vM�������=rn���u	S�"B3��o5e7%���H+���U��q'+2��`�O�j�N�	���M]�Jb�)eԥA�j�^ϱ���<Ғt���t����p����X��mn��Fȹ�i��=� �E�"k1dJ�a?d^A ������󔐧r�[ſ�Y�����q�����P1����� #��#����������Cfd<N�K72S�Tv`&����/x��|�bv�5��^�{nz�ݠ����"M0�`�j�����c���34����Tn�O�<�-���?�7�7�@�����  ����駾������C�s���N)x���e�2R��̩�=�ښ4p^���V[���<M�[�*�y�f�g?��2��0V��x�iC�f:���E�s�.�L����)������@��w��{n�<��D�^K6�md�c�pcs��yN���I]�$�����i�!�����9�x��=���b��ko@�[��E�S��y�a1�F�bf���W|��	�64졻V�#���޵_���d���є\[���0�h��9N�	���N�!�2�}���2c��?�ߝ��
���{��HI��z$��W}����7S��o=�|ֶ�����]b4�3R. f$ʠ̠\@egJ��%�Ȼ=�T�4�h��]�8T7�1�j�{ȷ#�i���f^���=�d�w=ܲ
	�1Hg�|_��O�Zb#��cE-cm����>AXj��T M�Z�iF��3ي{o�GE�z�E�8c�v�7�n�6��e��I-����#qs��F{J��w`f,�y+ �׽S��=Ӵ���Í�����WV��H7h�!�kO��6վT�#��N�l�N�E��O�2��e9~-�����!�xS�U�׾�19��?W��NH�w�ȥ�"��x{a�p����Zĺn���|r�j������!,}��}cu��o�2�T�6�;�n���1tKY�&�!{��1��]�}zߺ�F��t�*���ER;�H�t����ǯ����z��d�a��x��iW��Hcx��-`�*c�&�b�ns�z$�o�g�{/E$\#>����ЅQ��HIM����+$'�4AZ2O~� ��yM]#�ߌxn���%���L�ځ��ہ�̣��c @�b^�l��1.��cch��}=��&4��ƒD+oB�#��G=t�b��O�Jid�m������>uʫ��C��i�&�T+n%+n圁��){4���g�$��J��kB����ͥ��V�ƃ;�:�J]]w��{�X�?�:�&���=��������O�m�j���*V�����*C�=,�!���*č{��UD��������ݣ��q�=M�\���58.ɚw�iY{���tG����U�-��~���7�O�o~�e���� �il0�C��Ъ��m-r�� {�sB*;P�~�S���� ����x��:П}�{���9 ���r~+��H�X��ԭ4���}�o�@j�#]�^�*$ [KR+�#��W���s�Ƭqtݱ��m�|�6�]�ݲ$�|zYh[=�=��{zQ���f`�{CX��]cX=
�եz�e��i* 5�¾Ag"$����LDA}L����vA��!�Vo��t�2vۤ�o����j���ĭ>�s�����Jk��\,fqO:5+�Y@�����`�083L��&1���e0+r��guU(ߚ=�/��N(d1���WG�1!� �wX��̽���z�ͷ�kߓ�XQ�d�:x����I�H#W޽Y#)���:M̢���t�܈+�$K�d�f�]��D&I^�h9��� M٢>�w-���ugQ��������[�˼`�ŵ��ͫ��}{{���F?n����%��m�4����>��	�s귕��WHպt K���S����TPe��Ċ�#�ہ�Z3!g��tlW}k�Մ,�c��xh^Dp��Hy�Ϙ�)\ER-Z'	@�>Q�ڣ5↳�BU��?��7�������a����^{3D��m#�2ڂ\�������$"�w��;��9�8A�
��r��\ (�N`ڻQ[@y��Ȼ?��?�7�����?�7Ձ �����_�9,K��n�JOr��ip��0���P��NԚ�x!ء�:*K{���G�������c����_���pc����YĲ	k�Yi�L��M�0i�>�O7�77������ɼ,�l{H�7�Q�L�F&��5ܷ�R��0�> �c}����5�%��� 6���m8�/�Nv�j�$~	��A]<a�:s#\WEU=������hJ��-R��y�x>�Ɋ���p�4N���*�f�kǆ��q�'�:G˩E⑏��5�QJ��E��k;������0<�/tv�ֲ�"�PuHޓ��i�l�����'���f�71�:�^��)!!�Y�F�i��^��̮�X.���R�.��*VX^�6�Zl�^X��t�Ϭ�$C}r�n�I-��g�����]��^�W����X�����ӫ\k`�f
p̌R\��>�4�h�v�UR��5ۏjkX*0�Z{V6�͕dG� �_�{���P�u9�I��E���5r3��#�Q���-b7�"]���=j�Q�d��^6��SF*djp�<d�X�4y�������t����w�Agq�����~��K���7~���NzE~�HY���h2�7���rZ=��a�]�o�2�����,k���m�cV9�߬�'76Y�hm.pϫ��Pݶ*�o`�y>���r��e%�y�͐t%� �V�:B�6�I|��9#�y���@N	3^T}x��i; ų�ÓD����5�{�!�l��彘,�^$�)2Ī�uV�M�M� r[<�A�J��`��ŕK������J������@�N	�^��
4��Sww��3�^[/���ӄ=�8��I���Z�:�����������>+�X�����:�^�u[���՝t�+�48�b�/��	>�N���SO�)�&9�5�~h+e0'��m��R�C1��ٌͨ0���z��A��g�y��������@"t��q���z�7�\\��Ū��Vḧ́�ך�_l{�=�$�ު���j\�J���r7������f`8@�V�	)OÐ�V��d3�ن�����u]�P<m)^i,zlp]��v��{Iלޮ�n�l��gA�m+���Kߺt��"������ϻ<��2��	x% R�(�<�ly#�I=�)!BJ�א��s����2�^���A��xS� P���o{���?��~�����|K%��M~W�̓���0��F�Эƞ�j��e{�����@�l��l����]e<�}'H.[�19{xh�gW�z_���
�0�y1��؄�Z�W�ZG����f.���X7��X3#b҂ H�$s�x�i&{���3k��!^?K�ٔi��@���u���:�6a��#^6�x[�sU y�V`n ��y�P������h��=�f���\�b���m��	˲@!�rBNdS����̣*��|�K��]$�W�����f׍y�z�c�S&�������خ_���[���ӱ��f=�����}� aW��e1/�<$��{�잒��!�Ecm�׾�\���@+�2��<	��$���,�v_�쨧��K�6�MX�/����ֵ�][�_;����@�/k�}���~��x�ǟ��vcٌ�_����o�=K e��6�~Y��� MpCI��n͢�Sbp���^Y,(@"F���ڈ��LP�H �)��M�3�،G�{(6?\1�q[�G�H��U�p��9ҿ�h�����8�8��=j�w����!�c��E� W��8O�#�8'(gP��T�<�R�0=��~2��+ǫ{�=���Q�y����~��﨟�9�����Ͽ��?�����"G4,X����C���IA ��۵J�ԇ���R�^/���O�6w��鮘�mB�:�D-�	�.�V>�sQ�Jzh+���R�2]�!�ILloߋglZP?_��IU��b��EO*�����t �4r��mU�g�{}�ȉ�h۞���?��26�5f�!Cү
�MR�Q�Rd�3��n��{���K2V�,��V\^6<)�L��Vۨ�ruh�S �U�d�3 ���խg�!e3D̨i,:��յ���޻�cܧ�g���ՙ��z�F�9��SztC��9z����~���M�A ͞̳�1r�������WkU�|4e@���zw�}-[�;�-���}
��]�2�Ț 9����ģX�0���y�\�|���q�����#i��n?-g��=6�k=��n�z��X��kU���4��"�%'L�	9%;�`�L
挤�T9	@�l�Fk�4r��CY��
z���M�B܈�\�H٣~�������zQ�p��������7�����zU�Yn����n���zU���{�*m�ל���@��(Д�����7�\��mJ{ ����ɟh��}���aqޤ�it"�~����Ư��q�����OO	��1�H��֦�^A����e�B�aH����#T�k�]M���C�7��ƚ�G��.[WF�yzŪ=�ݳ{�_�(Z��Z�V��Y�_���'Q�VJ�D��Z����3�0��t�6v�����"����)ﯕ֜��ٕ�n�9n����X�g�W�ۡ�s�.w+�:Q�M��s���e��+\���-S�n�qy!x��@� R=�n��j/SL)#1#�Aa�2RS�g��L4[;���抔3���L�\@<�6����h��q2���zR�b���M�j�7����Gd���{�CZe�EٚK6.b�֘�(2sF��BW[ߍ�
2�L�T��y���!����sF+tqt�.��y��@/�Z��wz�Q<�]O���zM����Y@���U6��d�{�Q�p��l�x3 s:o�!o����{�Z��li��~�4M`2�k��b�dbO�JV1�'�ͧ�l�*���*cؑ�v9EWEi���O���Q5�e��`|@�����ݯ�*�D7��X�vO��,cF�f�z=Ł�ߏܻ/w.�^�z:]�L}w6c���{p��yO{����0s��e������ `�(~���ެ�it CB�s�(�|]./~��<x����0��ݽ�q�k7�M!��湨����z��u������X���æ�lv�&44���%��t�9��#��4<�ѿO�屛��L�������y�Խi �40��v��`$O(��K��;�m�%v��IM>��=3*(�9�++	�������ٟ{� �:Q�W�JU���QEէn	�������Z�
hJ�1-G\��oy�Ɗ��ZQ[C�L���PB.�zf��y����&X��V@����ē`i���PJ��eƝ�~���W��&�9�f�mk�p�)*�zlN{t	MҪ7��w�Ev������aHٌoej���v;�a�r�l:�P�6��&���N;H���A@*;�i�@��'s�tq	=��.�8����Ji�n��a3�'7�ӣo�`$�\9��#���l���#2�kH�+���p�ѝ��Þ+��I�^���}�Wd��[=���m���b��n����N>��B�x��-��V/n�����G�9m���\�\zAl�
jd����å�>i�H�!��G��,����U~�������H�)Rqs�~�	�ŏk�EG�f��;@��kDJ��C��Ɣ����2퐦�T&�r���i�������S�����7���M�M}�w����s�(>����������K*�	Q����˧���9���e�ՕP��=r`�ʔ,TBCAZ�^�Yվ S?�W�����z�h-�R�ԳC
O���Gچ�\�]�F�����Ⱦ �(�a��B��@�)���j���[�	9�0Q�!gܚv��.pQ�8�=&-��9!��vJ�>'�Z��ۃ��d�ѣ��MW�z���am�{# *r�P�̌&�|D�'���l��{��	g���A����V.�Z��ǓU�i��3�
�Q���a���	mO(��e^���b��dnD*NMq���'2���t+cAc=�t1��}3|��^�E���t�Ve�*���E�x��;��}^wJ}F��NH��9���=\��&{b��кN�y<�i�`KM`�ВВ��!*�߃�'!w��g0JbdΞN�ϚR�y�<��7d��(�ի����U�&��[����Nڣ?�Ag uY0��=?SA��K��郡l*[�N�
�� M7��6�<��#�,H�L�`ڡ���&�,�V�'IR�tEj{��p<][$*O�i�z��CS,�tid�r;��?�z�9���"M�������[Ov�)�S�Z��E�v��6y�.��3aҸX#�}��+Fl_�}��
'���#�����-��:X��D�+�?��2A��\,���`���:�>ޖk��G����S�7�o��C�3�0n������^~��9ܯi��+𣤺K������|�%՞�@nM{ۅ􇗺����V����V�@�W��X���K��m����xo9a��Dmآ�E���ƿ�W;���	9��5�o]�@2#%�BJ�����[�`���T�����3i�e������%v(v%SvO P����=����U��>%�BA���H�_o�̬Tv�DBDJ�oӴS����'䴳��4�ݑ[���Z��¢�V�dJzJl=����`�k(�C��&�s<����&03��Ќ�)�J.���-|�Kh�Q���D6��� �	�+�d��'2�'�����б�������Ƴ�j����ѾǤ;����/xލa߽)����?�+T��n#]6�\lP���*H:���(B"�5���R&P�x�M�4�����m*����S�˧�r@&'�V��o&���5ZU��`���Ƭ AM�A�H9�%e&eb]�E[�*M�*n����������N|�����M�D���'�UIDIUHd�Jċܴ��}��.��0�X�R�)_�̱��� ��?y;��3)Ӕ��_@�p�X�()�	cވ�Z_����dެx�@�!���RaKM�}��M$��IU��u5�!d�(�5�;F��(���F��7������7�S'=`�=#��h��SA�%���r�;�:��ns�3���j�������\��|Ͽ�����?1�2: ����_�ٟ��˸������{�=��$���酪���k��+���q�����f�KI���ja\/"���zC8b�=4z��r{@������G����xiKtE'�zPTm85A�#�d�c����>)I�"��gMH�(^�iyfFJJ9`��\pk���t�|�|@!k� '$0)Zv�>�����������S#JU�-��DG"����> ½�t���!�'�{<pՓ�^K[qF������
9��*�*�T�lҞiwU���v��}-�:�'ngpR�Xt�@p�GiIN��2��e�t\x8N[D��v�D�����E#B*��pk���-­���.����yL��X r��k�ivD�2���MWA���vf����^�E���Y�U@�!��. d*����
��Ҿ��4%�\4��!�"������3v���O@�L��K��'�O�佧��̤��&�ĩ1s#BUEm�.�<SJs���r:��� >NJ�>щ���隠G �rﵓ��"h'-j�,`���W��(���p��C�])�n�����>�|	�U=�&��-mr)��փjۋ�I[+R[��L��$���"�T��HZPX�XG�\���).��)��@�KL��Φ�ժh�J��Ac�>TB����H��nl,��&P����=� �
�V�Aɮ��;�ױH����}���I5��u�g���)#�؝��*S�g���X�H��{��}�E)�K��7��v~��,�Q���w�9���G?���
~���=�f��˷ԁ ������+��q���_hy����m���<1��k�/Q�"%ki�&Hb�0i�N�:���*&X�ܛ��x=��hxI8������V7�U�C&`l �U`Q�PSA&��V�'�W ~�0)R�P�ȔL�L2�0�f1QA��r��i�;�ܙ�`���<!���VA[`�ښ��Y����T���<�Ӄ������5f�� }�2^d�<����h͉+���ݾ*s��n���ҔX.�����2��r��Sʍ�y.Rk���&�eB]
8=U�߯����wcW���������T�E�ITx�j���P�'n)�4/x���Ǚ�JΦ���	9eH3)K&����S�>+n���pkG�mFW"D���+����}��6̨��m�.o�J]ꛣ�^�lm�Ex���~��Z�.���. �Z�����	uf�(�H�V��݄S�q:	��)���gԚ���%��ٕJ�n/|�����S��#_3�Cb<,�����_�į xE��,*ߨN/��[.��[ޕ�)7�,�rc��D¹4"m��kd�e�&Mx7)�De�k�,�jEz�Qr��m�@��r}dL�y*iJ�K�Xu�mn	@Zj˵�,�%�9Km���V淋���R���|�H}mym~B��Vkˡ-ׅuIB�mAʌ�����q��i�����B�N��]ɸ�`\��КE2
d)�vB����hb:]��HPP]Еۈ H��u�Ż+]�����dE�"����Q�;��'�#u�BDS�;oM�{爌Z�q&�a>�@0{�>���>xe�R�#O{�2]q�-�������������R�9�-x�v���Ox���_�{��Oѯ�ҿ���A^�E�� -&�)&<Cb櫶il��R����D��dZ��\���lz�{��f����!���&N��@2AQA3�넂v���z�����+de
��M�1MH�=�N9{�3�JW�c���].pw�w����z*C9!��Ҥ�,Dt��&ί���Μ��S�\N�O	��*��9O'N��ʇ%]ޞ?�3?]�|��r��R3���֟Ih�J���n(������-���Vlr�js�L��'���������9\\�5��Y�q}��YQ�KD�[k���i>��c��[A*Y/��P8=��J��e��yλ]�23@���5��ä�ĉh_wD�/3������?����²]KοNە�9���D�`P���F�1Е�[�pV(�GE�B��:V��� �MՆt:i�_B�	����Δ���K�Zv;�ۇ��R�I��x�s�j��P%���y��SO�r��xI�o�i�Uʻ_W�/���
PK�%���VJie�qj<q�����7e��[,�"��y+��v��	�fc�T2���tЗ#�X��'kgj3P��5�S�L�z���Pv�L��Ί4�EZ�5H���P����"�a������u��Xj�3Z�2�_��m^^���h�۲�g��nk�����T��z(:CeA[ԥ�-���e9��#)���.�*{Bk��:5��m� ���־�D6��SS��' $Ӽ��l�J�#��vng�k)��0A��}��1 h����n<EYi7587"<%��Z,�;��R��xJ;K#��W����^*��J���.>��[�����-w��K���>���4�˸n����?$*���/u~{�si���fH�!��0���n۵b-�=�
�<�����L7��^ �ʱb���߱�l	�W�pya��������+�
����`E6jU��.�֐S�R2�2!sƄl����1+ Ta�
�|�C����%����gO�6����v�2	8w�_Ki����/�gSΟL)����IR�s޵��V=<�T��'>����z[3CiBK�' �g�y�o�z��W�
 �ZѤbYf���=�����^�ƽ|��5?|�Wi̜H[�Z+��L�-;�tGTo�����E�u߄wJ�������rI�3Cs��I�LXTY]S��'��Ki��T�%����z,,`�jR�["�*-��GA��L{�`�-�z/�C�T�R��fPv�RR�uG�}k=�ѓ�Px�&�U�[U�U����Y��ki���R[b�K[�R�)�:/u��~��ݾ�P3�ք_���|Yr������?�z�g����4?q[�p!�ť�|K ��}�SH�ۨ8y����l5����5���?���x~���  �IK���eF���!��m/����y��Nz���г�������;�����<�xWP��@��Y󤏧X�+d�RL�XeW��Rk*��tD=^��%��i����������R���f7�Y�t���A�0N��st���6C��P<r�3�X�\� `��X���/�6ʀ���ƞ���P&Fd��N6��],���H��i�������N����������Oķ� ���G��w��~	iaҧ����.˿�d����&�TZ;B<N*�y7��f�M���G�X��+?Yŧƞ]�.�^A�!�⣴�͏Tتe��ײ�ի������z}�Wu����
h"̲`>��Dؗɫ��r�dNإ	S*&/��g�j�(�w8L�qQ.q�p�������S�Ň��ʴ�r�ʧ	��=�_�����WN��i*{-��|���~���r�0��	���	w��^�w�RI8=8�x\p}\���}������Z�ڽ{�ݿ�w�S��,���=,�	��D��,hMH�uB�ɋM�D�o\1e��.�rb�2A�k�+Q����c�i��~�wW�ֻ���-�N��d�x޷$i�95��Ě�sK��wAV��&a�=0�o�{�M�7\!�*)TD�6�(�q�nr�n�r�ׯ<���8����^�_k�
�gk��.tw�6P��2��O��/t~�{��S�[O���3�[���ew@��HE��}�F��7z������~�+XN�X���f`>bz�I��5˼�\�$e��I�i�z�b�E}7P���4�ҔT�����j|k�C�j}�&�,G���ꅔq<U\_/&*����4pݴ��6�c�F}*�����T� �#&��Z�u��Zunqs[|C
ٍK�Q�H�����5�m��
ǽ��vS!T�^�m�ZJ�۾�T.>���.��?�����C�,���#o�R�'�[�@���/�P2�_��SU����j�ai�;[��&kaZ���R����pk5�9Ϗ�$x.�+m?��O���#޾����6�ի�{�+|���k�W���Ҁ�r�um�>�S�������*6PD�]���p�i��~qUP+ �q��;�{�$��}Wn_�zpk��������y7}\���~��_�}��اtwH�����l��t���^���Ջ#ꬸ���)�N`͠�P�x��5�EЈQ�RFk%��u�_b�9����6L��z���X��^~���p��C���ⷿ�{s�U��g>j��`��p�O?�=}j��km~?D_$�}����\?�;�F�|��x�,f8���"g�����Ԅ�i�i^��+�
���r��;>&�%&y\=�]�pm{��u-�+�P�yʜ���M�Ȥ/{�ڏ�o�~��P8%3+��J�B����bG)#s��8�\v���)���xˋ|���?5���Η>�1(	��5�O?��?�aY�����I����iE�I[��XߢV�0�}h�o�ӽ���X#U" �/���i�-��ke�"�
WU������#��W��'�bC)���QR���(�$L����!>�b`�&ȑӄ[��ؕ���jŔn#c�D	�/���~�ٯ=y��������n�����ҧ_���$4��sϾѷ4��B?�a���{
����an3Z[px�����{���%Ǉ/��J��K��Z�k���bAkC&��^�M	�
�B8͋�N'@��i3/W�Zsx�����F%\�I���+���'�9#%B���d����)���pLލB��Z�l#Y}��	 2��4ٰ�4������k9��J�WA����>���8��-��7�������@�/|�ؽ�i\��h�G�y�����^�N��wf�ߩ�h�����Ui{�Z �Td��^��G��7mܫ��#��f���a�
}������J׆������,*�#� jC|��I��WhRQ�u�K���%d6�f���i���U����\���w��;O�}�c��̻>��/}�ݓ�s����p���7�6A ��_�E �VA�3�y��镯���t�.>Ȍ�6ײ���{ҖI*�r�2� ���s�>m�P���ٔ7��@��xS����]�>�
U�b5�UKIu�����e�i�GǞ�2��qA�x��y+RE`���{ΩW��(/�r?O��r��/Q��H��r��;���/E����=�;��O���`y������SO�vz[m�gAx*ߣ��Է�ջ"� �C2IUXUX��h��d5�㒮��R���Ůq4%+a����{�}�EM`B\���� �����MLPb7MP.>�E-4�4�\�����������������O��,������e���[Z��?��O �^�����>�j~��[o� <xG=]�u��
�>��{���і;m^��T8^�Z5u����54��mmV5�&�'o
�v�k�z#�����3!�U���(q#2��ܵ!o(��p�˔�g��I�.�,̩��2_'N��k����?���?���^�� ��}��F���t~��[��?�ҳ��P��׸x�S}����[h�Ro�N"����P}Z���[*8a�������խ����c_q��
���7�.?IB�,�m��*����>�0��וf�����m���5-˂��Jɨb�1S.Z�W%O��������px�s���/�{�ٷ�-�<�����o�� �g�ԧ���x�|��� rxn�,�����6�<S8�J�U��o"z��o�N�Ts���(��yO
�jz6O���"������
�6C����ܭ-nk�$))aۤ>�i�2"��2%%NB����J�f%>�
����K�ӗ�����qY꧙���F�^|I_��R�L�Uo{���ѷﷄfw�/|�v�j5��@� /����#K]�&�h�Y[M�IRQ6�g"�邈n�-�iOL;UL
ͤH`Ndc���X��J�d�G�*T�`�FB��5���B}�+��De�8-3��#�*�2�~�'�V�J�����<����������O������/�u�4��|��ѷ"�JT�}�8�M����p��~�N��p:ͻZka���:�D�ۙ���������nI�Q�h�k�y^��T91133)"�b��f��@�Y�Z�\r΀���W��X))1	@ں�-�1QQc�
�
�3���9�gN���U��N���,���>+���S�S^��N������¯��'�
�����w?�Y�؏��}�� � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � � ��1�Ӓ������   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X    IEND�B`�PK
     E"BYd��   �   /   images/a262aa33-74c4-460b-b0ad-c746896f6744.png�PNG

   IHDR   d   d   p�T   gAMA  ���a   	pHYs     ��   %tEXtdate:create 2019-08-11T01:25:28+00:00�d�B   %tEXtdate:modify 2019-07-26T05:04:57+00:00�_�X  �IDATx��{y���u׹���Z�j��ez�����L�b'������2�eH$BaJ�@�dC��`�@��![G6NlϒqO{2��=��RU]{��ۿ�����1�'��n�u�{�[�=�s~�w��ʥ��1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�lL �1d���1@�l�c@�a�z��Ti�R��)�|�H)����]ǧ0�Vg�¸K�F�Z���=:0��y��8L^a�&����4�"ϨH32ʐv4������>Y��6����=�n� ��w�H��)�~�����t�g��!�<T~V�Yz`�����j����ר�����Z�:@N�NF�ޢ���,S�ޠ��NY<�Zk��J��� m
& ̡T�nW���]����{}*f��>s���m�ݽ㯐[����u��)h~�����>�����R����h_�М�NݴC͠���ޘ�g>�?���g�~��P�R8葉ڤ+�T�O�8�,�`�UZ�	!�n�6�a���y6O"ǭVk��D o�D9~G��[�m���^�u�'^"�[^���O�N����+ DF�u
��v�����/M2�P���&���8\��
\��w�z��V�K3�K3���h㇟|������~ݟ����W���f�ȉCD�M"�!Y֕�.���n�Sf�	ch��G�&�q�H5���*o/��%�ݼIj��KI�Z����.J[�(�\ׇGk2�j�4���X:
A�tԿ�M?�Yg����K_����pkC通K�23�*0o�g3�$����0�v�g~�/+�W7��|��ּ�,un_����� I;���\��u��_},�~�n@"��-ob+b�v��X�I��f�L]�Һ^��U�8�E'?vV�x�C�k�;���M�}$�DLi�S����mQ�Ņ�:��(_Ug�����F�����	��ġ`VcrDqf*��q
4SU�NLm&U^�������G��i�8�3�.�۩.tؙ9|fp�[�D����W)�lSg}�����ѡ��0���%�]���pa�[���>PD���~󧢵�� �v���ԡ�����?�j�UZ��ε��@��_
��e���,�=McB�'�pt�&���.���
{^�K�zst���t��I��#���\N������r���4a�8&:��i�M����fS޻�0�*N�� ��%
V^��'B�%���w�1�@��Yuh$L�wQ&�0�3��	B8f��e�wA���Hi��%�?�p-,$|M^�0$ln���ÃN��'���S���;u���}���~g�| ��eP�>Gӧ>�����)3���I�+Q$d���򼴍�*ձ�aѣ�x�M�"D�ܤ,=E��Cdẝ��HKb�=~���kur��0!�-�)���!��D��)�px0D!�`����!��YҞ+sU9��x�T�J�,�OR@do6v�"�J��:������gB�K���E�����Ԡ?±��� ����s�Kh���+��7^mn����&]
wV�:{���i��u�Z�|�I��'��&��=�{��֠}m�r�<�r � ��c%ED��*�	���8k�0�Z��5�׃S�w����i@�g�ׅ�âz��w[�D'��I�Ar<��a�L*�އ\M����G�+�+��߰s[�����
��T�l1�z��=��.� �v+r�v��[�D�KO��c�	�K�N����[_|���S\�m#$ł��y��s��~)�oR�"�qm�ߵU�/�ԃpw��
"��U��2��Nڦ�<���w]B�^�X�U�F�ozZ�3d��(w�m����&�ҳɂ�d^J��)$��D� ]��X0�*\KIy,`Z�S�oا\G�څ��k�ԫ����G(4ED�+�i8���\r;Y_�Fa�bn���V�`���܉'�n��z �}G����#7��{�B���/ga�`:��v!{�%Z�A�q�P�w���~CYT�UM@u�C�D&�����m�O���KY`��Cs5�e@Q�f�\Z�m��-�%*$4�H`ٟ�i2WD�L]VCq�)�~�dQE�:�)IX˵喝
��O=E>U�)��:[[��Bβ�saȜF3�`H)E1��>>CN�?оs������=��;k�.�$�ҩ��x�~���p��_Α7�p�&q�@NTNu����	yф���ά�K���	]�WQ�6���p^S7����N�z��7e�WY��G�95�F��+�ÁBሚ�t�D�,UX�/��p $o�T(M{5�ր�2�gBrNa��r����
�7_׃s̟z���S��\!3X#߳�7��0��p�3��<��D4��Y���b4~�:��˝�7^�H,P��J�ܰ�K핛tv�y��'�w���y�����a2UNQ��8���/#z��!X�4Ee�w�.���9��� �ޙш���.U�5rI?��H�>��!���~�
S%6Y!
F��[ͪJ�亢�"PNтĚ�Ҿ��\�*Ȫ"�윬c�*#��%j��}���y�����﵌r+���Q����5��#w�<� o`Nٰ]M�꿞=��3������i#$�z,�Sm��}ݕ��}�{���ޑ(P���̄ZP^U<P��7�E�)s��p� �Jg�"L��s���8=�8�&Q&	�A@����d��U��Z%p@ e�w�C�� jT���xbn�[惟^��.�ӶxmhI�R�8��X[;��Dn�E~�^��WR# j.�5�RX�_�r�+��]�ʜ-��"���^�t늬դ^��G� x�s�⿸���ԉ?��Q���:�o��� j���g㝫���8��/�(���E�a���r��j�Tܻa/k8S�PY$����I:9s��;��1�M��0RE��<�Rھ��DR�y�2���D�*��$�ETdF�(�8*4�uD)1{6G�����@]-��=F���r��q����0��؜(y�s����@onm/;1�y�&�'����YH��.�KT]xP���SY2�A9qE���	r��������������έ����{>�����@S��/�c��eu��ʘ���	9%�Qڪ��x�"�4a�$ۡN�o��t���"��Z�m�O�ȉ�/SmΞ���%���b[�Ap�����29?gi�IH+�� p"��� xH_�\U�#�8 �=���� �Ʈ��Π�P|9�G�ex����)ݥT�$��5����)L��H��=�c-9Q��3�C���"��BS��4�=w9Z~j;�~����i�ě�}Ű"a��$�ڝ{<��X�1x;"g U.�*Y-���$�0��=��FG*��wi�f���zK�l^���~M��!t`����E�ޗ��5@���R�3�7(T�rl��<��T��;D5�PD��ѹ���d����\�p�!ё�I�#&��Hn=�Afa������[�M�����ox(�}��jߑ5*8�ҷ��D]�kduƵX���E��e��g���s5��w: +�KaS��q��0Y*rc�dZR��+J�*�G�Zc���"4A30��7���ޯ�Q�/�޸D���xs��D�p���.a����6�9%�3ա��XYn�"L[�˭"� �� 1��MR��(a�F��Pcs�6���w�UD#�ƴ�k�:&g�ɻ��P����]^[U��գ�W�s�%���@X���f�S�?��:	���.�B�r8�魐��57�ڛ'�G�͢�k�$�\.�Ӳ3�������|�R�|�|�܁�ڴ���P-���ץ�+Qhlo�)�^��˹!;�S��1C'�aT����Uz+�t�$½�;j�9�d(t��x����m�0H�Հ�"�Yi��BT������5���8R��/6�̽L�FKn�M_r;4��<�\�؊K�E~�%ut���ص;�2��e�@4�����*kY4S���X/���9������
�Y
p=���8�8,Xp��ͽʶ,�{F�>Q�H�Q�Ĩ�SCsnF���g���T���胁őX���}d�$PJR�_Ξ)�
���֠�hGh[���j����'M1��'�>�Hd�D5��8R��,
k"�Y!���C��\Ŕ�AqY�(7��=�b�H�Kr6���e�Nو+_2Kc�����]9ڪ�£���a�Y)@+[3N���?�u@Y�I��2�a^I
��a�|&R��e/Ki�Y����������<}8���$i��{{*2m��"��ZjF�R9\ c�YZ���V�#�j)y�*j�Pj�T))6�����Q�Ƥq��(؟���Z�K�כ�ό��bЃ�l%"w6�s9j�k^\	�m��J� ą�|�(�MҜ[_$9��.e�h5e��ؾ�eJ�F�M0>ߵ�����C���W��4n�&8A�{�^�U,|^x[]��~{�/ۓ��S���r�*��VM:�Ibh*,J2�{`PY��-s�&BU�S��!b%f6zx�"(���u��_NM��ϯ�]	p���[ِ�������C(A��ʚ�&V�%n��Ҳ��m��XZ)�77�lH>�~X���w>�ⴇ�P8Y��e�z��>�!,�S�}%�[��˕�P$+!g�0��Qd�F��-¬��X5�@�iPE�vٟa�T�r7����hޅme���-�a�����Ɣ��;GМ��`��?��{��~�ɿ��'�������C�r.r��Hf@�޾�ѹ���J�ƲЛ�J8����1��� B.N0���=6ۈ3ei��0����E+<÷�V�sI���ϋ{=)�[Q�����#�Ap$�r��q�a(�`�FQО�Y��jî1��X�~�ʍ����C��V!��e���z�3�r�[)W�`�'��?�%��_x���gg�~�Gk�7l>�UH��E�ǡ.J!�dv��:�Ք&�6N���&�1�Ri3צ��=#*�!>�
�mI��P�{�0$j����쵲�ABf�Y֒#����j�����K+GDA�iy_dv�Q��M��T�b���xm.��P�vű|����g�e�X:�JP�W�})B����qQ���H��=���t{��?;�U2�1�	���`���'�~?l.���!Q�w+gD��w��<F��8� ��#$�I�G^�Aa)�un��-O!
c�	����ԋ
�	i(6;��R��	�����|#M�RJd�sRa��
VO^'ANL��Y�k���PY��6��Z��<mMf7�4�t&{,E)�*v�t$F[��1!,�Y�y�s������}2;7YW�����c�q�u�x��T_,.y�}?}�y��,�Ӱc���Z��团�`����)&��|,Q�%�3�Z�T���OD�R����M�όy����|DJ�s�<���O(]��Yx�L�|��X�ǀ�ANY�ؘ 2��H0/n]��z�̍�s�B$+D���"Ys3�T�
Z9?�`NY�h$�(ͲQj�cIQe�_�)��T�~.�t�̳�z�U:�����!�����(��+/�����_s���n�E}��P�{o�����\P���r���J*@S)GG����Ae!ȋ�G\^���P4l�ݞO��+�;�,�}!<��F�R�L���=T`��v������[C�����8/QV�I��@�[�%���-s"� d����uH2��<�P1��:h��gI>�b��I�ѯ�Ch5�������7���st�]��\�v�~7-_x�K��c����YtH��O�-��:�F�"iK�\Ŀ�׏���4�ϐ�x��
�d���Y���Oi+���V���!���h�w�e
 Ң)�;�YِR;@nom��@O���#&���V��UBq���ͯE�.E��4�΂+�5YO�{�F��`d�mp_>��A�Q/���t���h�(��;�_�Ï�|���|����k����W�n�u�1��H꿡������H1��;�^�[��dQ!G��Ȇ2�@qN��A!)�k�ҶVE�V��u2��f�u�k$xn��(0p��]6�F�DSFF!^���+
��l��?W�yn��\Ԡ)v(�6�r�u$��k�
PEO!���$c��'�,]
�Q=�st�t�\���ׇ^�������yo����G����!�v@fg��k/����?���������S�ҡbЅ��e�~i+e%BVG��b�f�n��Cb,�N�w���Ƚ �T�k\�K��'���V��h���]�B�� ^�>]�����lM+�wJ�2u������5)Ly�2�MR�UI5�}��L��k1����k�	oN9Vy�߇�#Y1a;T�&�.����í�~��c������c��i���?0��e|�)�u�T���[itď��FC��'�Oūx��i�\�s����3Μ�-���'���*��jו�6$���-��4��"k����z��J�Z��sը�Pvo]B5��\Q�{߳5�[%g��ٽ)8�eC��0�,~F�_�J��@t�4U�*(�R��#��>�M-�hQ�3�܀�t�m�e�l�a=^s��������~�wx�̇�w�������K��|�vV.��}�?���?b��;����"�e��=�f/.��kT_���En��u:��!j֏H����V��|W;^�K���MD���*��4���AUy���Ss)�f������|��#;���.�u ɎHw���.!��#К��BZG�����8�%��N5O�zGSY�u'�}����O\B� ��Ȯ�H�N���a�'.j�.Ҝ�g)�#p+Ti-Qe��E����a{c��n.�������ճF��w6�S'�������:���H�}R�sn)���>���z�&�3�Uϣ�?M3�����Go�V�3����W_s+��&��N/�G�+���Q���Yz���k۝f�f�����@{��㙄�"����Ju��9�r�i�v������������X��� �:��LT��N{�/)<L����l߭;�f�y�5����ߗ{�<r����.��y/��^"�@�ZI=�F?s �<8^0��U�s���t�s;���H�}oJ��y�V_y�q�����d�����~�v>��n�%G GS+]A1��4��x*�������D�ۊW�=W��k�>��/]�򯷛G���	��P�_'�*�.kqgv{��RoQ7�d�*qR
}EQ��0�і���|�>9Bൕ�e2�-�i��,�bؕ=>'K�w6h8�KG��� `<PRvP<�)���y���?�ɠw��G%�:��=SSt�0Eu�婙�H�Z��S�z��M�yם��?[�N����s�<E5�X�����w3���}ȁG�CwΝ�J����is��*4������V��6}���ȼ���T+�����ڌ)	w�9�_����W~��W.�C��%ZlP-h������}/^�L?N/|�b`|P��֚l�nܜ��U�y�ؗ��ڇ2�[��}�[����<t9`@K���w:�W_���BՇ�{典H�o�4�f��2-��_���[�p�C��
��9.'u!\1���tz�5|�|��>t���W�9��D<����Auߙ'�~�s�"�?�7i��D�����G~��_{)�]D�D��.
ɵΦ��j[Mz��ץg�͆t����q����r�N<�m�W.~���CTi�݋�%�W�ƉluKu�P����FS��5����� ~i�~��wt�?�}�w�����O��O���wf��c�W�c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2fcȘ�	 c6&��٘ 2f�D�{��w��    IEND�B`�PK
     E"BY?S�2� 2� /   images/da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.png�PNG

   IHDR  �  %   ���   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���   �����
                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                              �ك     ��FPUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUUU&��M    IDATUUUUUUUUUUUUUUUUUUUUUUUUUUUa�ޟ<+;�?�9���/s��f a *�K e'�P��xvf m�T�w�����a��j�T*��$f�V�4j,%� 1\gg�/����y�/�*�9}y�~���~<���                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                         ��Ū    �jkw�yIou������h�g�R��e�qQ��c��,�RY�Y�"�zL�ʲ�~�u+!OE�N)e�,���w˲lǔ�B)�!�����t�
)���\J)Ʋl��/e�8Ƙ~��S�Ն?��$�X�B��̲l�S�;�1�1�eE�qc��,�Gy��2���eEȲ�"����s���hƸ�5���x�ޙ�Y�����k��      �>�   ؒ����p�g4���c�UŮ,�]�t����L*˙�,gBJ�4�v��e��R���l��hƲ�������B�y>IY6y>�Y6.c�dY6�Z?fY?��/c�Y֋Y�k��)��q���Z�|Q��Z�����?      ��;    �IǏg?x�ˋ�bJ�EqIao(��yY·��+�r.�L*�nV�4���tڊ�m�h)�k�Q��)��1�7R���Zm=ĸZd�jȲ�!��!��b|)��ԥ�_�B<~���     ���!     LZ\����WN���8�.Eqi-ƽ�(�Ĳ�U��{�-�b&N&�4��չ�R)��T���<�Zm-���S���<?7M�l��?H�کZQ�`_��|\Z*��     �)   ��]wu_8�@=�ק�|}*�KCY�e9'�=i:����0ͅ���{���Qj4zY�����)�{)���Z�T-�_HY�Bʲ����T�
     ���   �`iq1a0�:��`*�+�x��T���$M&{�d2����X���[a��y>I��Z���b�~����,;���,;���g�����     ���   lc'?��+C���,���drE^��䒬(v��xw�L:n\��'�X�z���e������<?���z���d�ԁ�z��N     ���   la�...��7���XN&cQ싓ɞ4�K��X����W&�X�fs=��gC�~>���P�=_k4�N��w�e�w��Ҹ�N     �ׂ�;   �&�{�߿&���N��_��q2�4����pxI*�ZՍ�ŕb,c�������8����z��㓡^lay�LՍ      ���;   @�N�v۵�,�K��~z�F�ݡ(�U�[L�6L�湬�x)��_L����,{���z�ɪ�      ~w   �����Ņ�`������`6_�����p�'�e��>`g�1��\���h<j��k��ө����O|��U�     �   \ �>���j]��F��S��r<����p��M��������f�ƩT�?�'S������?ZZT�     ��    �Щc����五��x|m����eq8�R��^b,C�������:j�'k���Ӣ�ځ�z��<     `{q�
   ��X\�,�ظ)��[�h�r4�<�F��dҩ�`3��F/6��S��B�����E������SU�     [��;   �����b�����drS����+�h���]U�lIy>
����n?j�'S��x��|����sU�     ���;   �c��﮿x��i:�1N&����W����l2�K)yO�J!��l�f����h<���;e�����f���I�}     ����   ؖ֎�۟L�^����h��0\�KSQԪn�'b�E�j�d���E��O�f�Q��wW,-�Xu     p��   [ީc��R�F7���8]�����h4�Vv��)Ƙ�Fc5�tN����E���q���+�����     �זC^   `K9q�o���o����a8|S��x}�N;Uwp��(��gB��Lh6�����{�;�Ǐ�U�     ��;   �i�c�~��0����`�y��F�kqi��:     x��  �M��m�][�͵���p����EѬ��-(�GY��´�z��h<2��o/�'��     ^��;   pѭ�y�%�kk��drc>����!��Uw������9Z���������XZz��,     �g�   ��G����77��w���-�`pU�v���� �2)�����v�ټ�z��j�Þ+���x�=���     `'s�   \P+G�^3�ߓ&���~�-�׻*��W� /'�X�v�L�v���oO���^y��OT�     ;��;   ���ƙ���b8�9�F�Q�`���. �`�����>S�Z��z���w:shiiPu     lW�   ���s��~is8|�n��ᵡ߿,E��. �XR�Mb��b�t�(k������,,/���     �w   �Z9z���dr8��
צ~�> ~V����'B�����������U'    �V�@   ���w���b0�a0�!��o���ު� `˩�7b��L�j=Zk4������/��    ����   v�t����'O�'���-��W��Uu l;�Z?t��+��oN��W��~%.-Ug    �fd�   ;DZ\�ό��*�Û�`pS���h� _ʲq��(��G�F�s���/�    ���  �6e� [��;     ���;   l#��94>�7�^��Pͪ� �W�V�n����~���?w��?�p�I     p��  �v��[�.Cx_����ׯK��l�M �V��c��tj�nt:˗,/�S�I     �Z1p  �-d�ر������~��ac�m��_��	 ��Z����>;��;��KK��N    ���   6�G�^�l�R���-76ޖ�����< �bL��9��GC���݇--��    �Wˁ8   l2���E�wkn*�ׯ�EѨ�	 �b�OC��|��>�7�[x��/T�     ���;   T��ѣ�&Eqx��0���#��U7 �D����'b���h|bay�L�I     ���  �E��66�c�N�7��n������ ��-�Xf���C����l~f�����TT�     ?��   .��n����ht4���kko�I��& `���qf�43���K��    ��  �k��w�u����ol*{���-� �fc
���0;�������n�b<~��:    ����   .�s������}�~��qu��4�V� �4kav����|��h|lny�l�I     ��   �+8u��u���C���C�׻*��W� p!�,�����N���n�c�[^~��&     �/w   x�N9r���7���+�SJ���#��g���7R����o| ?^V�    ���    ^F���K++�L������x<Su ��P�������y��t���}��U'    ���  ��q�����C�׻9�zoHEQ��	 `3KY6N������~��v��KK/V�    ��c�   ���#G~=��76�^�`H)��	 `K�1�n��43��N����[U'    �5�  ���>r��t08{�76.O)yV ��R�}6��}5k6?���_��    ��ˡ=   ;JZ\�O7���
kk���U7 �(��J���Vj�>y���Ǐ�U'    �y�  ����Ɖ��;j���am��a2�V� @��X����v�ӗ^~����N�n    �Z�   lK���'_|�q8�=���3L&���  �%j�a��{<t:.\s�G�=���N    ��3p  `���Q����өQ; �Vd�    �c�  ��� ls��     ;��;   [N��?n�y�M�׏d��ׅ�hV� �EP����7c��Ʌv{9.-U'    pa�  �%����d���� !��h����7R���7��@<~���	    �_��;   ���#G�އ���o��x��  6��j���ه'�ֽW>��#U�     ���  ��>r�P���nX]}OwW� �֑��a~��N���g��    ��1p  `S8}�o���X���'{�� `��1ř������v�-,/��:	    ��g�  @e�]\\hnl�^\]�%�zW��<� p���47�T���|������ݷRu     ?��    գ�w��j
�ޱ����R^u  ;H�����c��yp������4�:	    ��0p  �5����-q8�=�?S�N[U7 @�Նa~�S���x�����$    ����  ����#G�^�����o��x��  ��Z��a~�˵n���oU�    �S�  pA=����\[�HX_�@�����  ^�N�T97�7i~�O�XZz��    ����  �_Y����K?���bu�����SJy�M  �+������	33���_ť�q�I     ۝�;   ���#G�އ��ʻ�dҩ�  ^+�����o���??���~��    ����  �W��m���)VV���uU�  �Ŗ�����gF��zpi�T�=     ۉ�;   /+-.�/�w���_���%��U�  U�1a~�;���_����?�/�n    ���  ��N�v۵i4�H<w��a<���  6��h�����ess�,,/?^u    �Ve�  ��x����z�����^�ꔒgG  �7J!�lv�{a׮�?�������A�M     [��   !�N9r���>Ο��0���� �-/�Ga׮G�����O}��U�     l�   ;�ڱc{{��nK����{  `ۚ�9����?p�%�=��_lT�    �Y�  �@'n����`�ùs7��hV�  ;ƿ�����������U�     l6�   ;ģ�w���VV~'��_Su  �x33'���]���?���3�:    `30p  ���=����������ɤ]u  ����7®]_����YX^~��    �*�  lCiq1i8�c��򑸶�����?  ��R)���^ص���]����{'U7    \l   ���ѣ�l���5;�����;���.�|�<�h�,ɒ��q��)KK
��=m;Rb�
n�a�f�iKSZ�����2���4t:�-�;�q�b'Mo�mg���8޴[�%Y:�<�7��[ ;����~�o��_��}~
��{  �g��j&Y�����ʛ7��{(v    �R1p  X�>�=���.LM]�����  �i�fIS�w�MM���K.�J�kW9v    �b2p  X���oo/��^�NL��ͱ{  �EVS3����bC��o�����9     ���  `��<;��tb��\���  ,�4����Uhh����u�_��    8��  V��mۚ�O��>LN^��<�!v  �<���cIs��,���{�l�    �3e�  ��Mn�v���쇒�ǯHJ���=  �2UQ1��_�?��՟ٴw��s     �-w  �eh����03�3LL�,	!�  X�4͒������}��{b�     �.w  �e"\}�ГO�+LL�5��97v  ��54Iׯ�rg]�Ӿ�B�    �Sa�  ������������B��.v  ����L���{MM7���7;    ��1p  ���UW]R9?}:>��e�{  ��-�r�t��of���=�����    ���  ,��ۛ��Sir�]���ܗ  K*$IH���[����.��+�]��M     O3�   XGz{[������oJO�l��  �$I����l�    IDAT���;�r�ʻ�    `�  ���tw?7�������+�R�&v  �3���K֯�����lڻ���9    ��e�  ����/33;���˒r�{   NE��Y����|C����{O�    `�1p  8K���H��ޖ��u��  8#��L��������t׮r�    `m0p  8C����n��ݙ��]��Ϸ��  8�Bm�h��z[W}��}}��=    ��f�  �,Mo��:=;�������Ph��  ��Қ������uMM�n�뛊�    �N�   �i`���$����ؕI�U��  XR��'���{��}j����    Vw  �S4��7]�MNސ?��P.W��  �)�狡���Om����    X�  ~�����'33�$!��  �g�4͒�뿕54|f�]w��    X�3   ~�cW]uu:=��dj�y�[   ���$!mj�n���s�����    X��  ���ۛ����剉����c�   �HG���?�|�+�K�kW9v    �r�  $Ir_oo���ٝ���u��|K�  �� ��	--�����Ҿ�B�    `�3p  ִ���[�gg?�ߞ
�{   V���f*kn�j]Sӧ[���b�     ˗�;  �&l������G���7�YV�  `M���K[Z�ַ�}����b�     ˏ�;  ���������b�b�  G��
ik���kl�x���#�{    ����  Xzz�K��>���_��"v   �4t_hi������b�     ��  ���֭�I>j�  �|�    O3p  V��ۏ�,�ˆ�   +��C�BSӮͷ�>�    Xz�  ��2��s~yn�F�v  ��+�狡��k��    ���  ��@O����ڰ  `u�ǡ�����n���?�    X|�  ��6�}���ӿ����&	!�  ����    �w  `E2l  X{���kj~�cϞ'c�     g��;  ����T��|${M0l  X�B.WL[[�   `2p  V�v   �����u��}���;���    �9w  `Y��y^:3�+���"	!�  ��'�r�|k��曚vm�����=    ��g�  ,KGz{�ɏ��Zz��e�\���  �����������5�v�X�    ���  �ʑ�ޖ��ԍ���5I�U��  `��8���7vtܔ~�K��s    �Sg�  ,����n����dl캤X���  �ʗVU����u56~:��+��    ~4w   ��ۛ���Q~Z(4��  `��=��������q�kW9v    ���  Q�]�rC�������������=   �~��~��������=v    ��� �%7���������\g�   ֠��#���Ϝ��G�    �_2p  ��`Oϖ0>���ĉ�c�   @�n����}��{����-    �?0p  ��5�\Z���1LN^�   ���$!���H��������=    ���  ���5׼�rz�?&��JBp�  ��Ҵ���<�����{�<�    �*  ���9/���X:6��!�|�   8U!�+���_�56~�s���=    ���  g��������'��㗅r�"v   <k�������H�����9    �V�  g,\}����b2:z]R*���  ��%TUͤ��_�jl����/��    ���;  pFFzz�\�Hz�d[�   X,��n0ݰ�w6����    V3w  �Y�<>��dffs�   X2MM�+Z[ol�㎇b�    �jd�  ���[�^�;yrW8~�U�{
   ֠��崥偤��ƍ���c�    �jb�  ���mۚO��ޔ��^���=   ]E�|hk��X����{�    ���;  �C��������'���N����=   ����L�6|���/��t׮r�    X�� �h�������/�����-   �܅��c��哛����    V*w  ��8����tr�tj��c�   �J��iH��Iׯ�X�w>�    Vw  ���tw?7?;{S2>��$�   �,��\)���uC{��o�m,v    �+  @2���trj�c���4˪b�   ��QQq�����s��>���b�    �rg�  kX��������;�B�1v   �Z���Ӷ�[������)    ��� �5�ӳ-��07��   ֊���{Ys��7�u���[    `92p �5�Hw�s+ff~;���$���    �Z�������56~�s���9    ���  ������w��ӑ����rU�   X�*+g���?�jl����/��    ˁ�;  �G�n}sz����'O��n   ��PW7�۰�7�����    �� �*6�m�K�������n   ~��$!���ºu7l��?�    b1p �U�-[�+�>���t'!�c�    �(�_(o����ټ�7�/|�;    ���;  �2�[��3�p��o��   <;i]�p�����ٳ竱[    `)� �*q�������O���ύ�   ��4MC���Hhj�������{    `)� �
7�m[���ٛґ��B>v   pv�\��nذw4M?��{�    ���  V��kWn��_�p2<���X���   ,��������{�~)v
    ,w  X�uw_V9>�+��97v   �Ě���ZZ~���;��    g��;  � O]{mW���o'cc�KBp=   kT�˕{WT|��w�=�    ��  X�C�4�5ɲ��=   ��������[�ٳ狱[    �l0p �e���W��jj����sb�    �TS��bK�Ϲ��Gc�    ��0p �ej���i~|�w����IB���   ��4�/���=]�{�G��}n!v    <�  ��l������I���   XYҺ��dÆ]]��w�n   ��e�  �ȑ���V���v���-   ���$����7tv~����b�    ��2p �e �����%���#Ͳ��=   �*QY9�tt|q�޽7�N   �Sa�  �vw��|��'��ٍ�[   ��)45}����Ϲ��Gc�    �c�  �Ll��|�ĉ�I��.OBpm   ,�4�/���=O57�xi_���=    �L�h   ���[ߙ���BXXh��   �-i]�H�aïw����    �5w  XBG����NMݜ��zQ�   `�
I����:;?�x�mc�{    �i�  �Booձ����##oI���=    I�$Ie�l���ō{��;    ���  ��-[ޘNN�f:;�1v   �3	MM�ͷ��b���ߎ�   ��f�  �dh�������&cc�KBp�   ,ki>_
mm{�jn��Ҿ���{    X��l  `l���td�áPh��   p:Һ��a��7����   ����  ΢�����cc7'Ǐ_�   �YK�r���w���}x�wL��   `�0p ��d�v���%�bm�   ��!TWO���qϞ�c�    �6� ���9?LO�&&^�   �lK�4����������7�   ����  ���UW���JJ%��   �Z����ut�fמ=}�[    X�� �Y�ܶ킓�㷄���n   X*O�����|}����c�    ��� �i��S�>)�jb�    DQU5]jo�����-v
    ���;  ��C�\���o	���.v   �r�67�[hk{���o��   ��`�  ?Bص+7x��7���w��rU�   �e��r6tv�|Ξ=_��   ��g�  ?��5׼(����p�ď�n   X����}���������   ��e�  ���S�ӑ�w�,���   �"TVΕ;:nٴw��c�    �2� ��2�m�K���φ��ͱ[    V���y_hj�����ñ[    XY� ���ުcSSϏ��\Ȳ��=    +ZE�\��y�ƽ{o��   ��a�  I�_sͥ���O���c�    �&����������?�   ���� �5-�ڕ���ӑ�w9�   `�TV�̵���y��;   ���� �5kl���FF�09q���-    kA�ܼo��c��}}C�[    X�� X���jg�p�eձ[    ֔��餽���{��E�    �w  ֔���ۓ��ϗ��_�   `�J�4�������Ë�w6v    ˇ�;  k��֭oMGF>
���-  ��U\pAe~Ӧ���p)��SS�$��Y ,C��v,��|d��w-v    ˃�;  ��[�4�W(ܒ���.��  Y��s*�~�g��ai(C���,����Yyx8ˎό�H�$	iZN�����?���/|��   ���{  X�F�n�2�d��o��  kE��'�@S����g�aa!�'&�?zώ-����K�	�2S_�����w��P�    �1p `U
��U�������\�8�  �\ݛ�ܐ��8������Ѭ4<��GF�lp�������|������ƿ��O�n    C  V���ݯʍ��~27��  ֪�W����Kj���'�lh(+f�GK���YRv�;�����x][���;�x"v
    K�� �U#�ڕ���ӑ�w�,;��" ������+j����l��P*���X�����,;v�����UT̅��Ϝ�g�c�    �t� Xƶo~ad��'Ώ�  $IRU��{���4]���!���d�<8X*d���,��w��Җ�o֯_���ݻ��n   `�� ��^u��00��$˪c�   �������Z[�K�{��\�<:��JٱcYyh�2�w��,���
�������-    ,.w  V����ۓ��ϗ��_�  ������ڪ�(����T
ah�T��ǎ��c��V��$!ݰ�o�ji�yi_���=    ,w  V���[ߚ,)�c�   Ϭ�yϫ����w�B(��e�#GJ��å��Q�w�$���6l����b�    p�� ����ު������W��g `YKr�~wc�)�Byp�Nx0xX�\����߶��{?�   ���  �ch����CC�Ofg7�n  NMû޵.]�.��t�R)���R��އ��$��Y <���o/tv�������)    ��  �[��?��$˪c�   ����+�*~�ǫbw��P,�0<l��L����iG��:ﺫ?v    g�� �e�-[�+nIFG_�  8}�/zQU��X��l
'O��c�J���*�*���r�&�5/M�I{{Ws�i__;   �g�� �e�Pw�eU##���[b�   �N��%W���5��XL�ĉ���S��'��ѣ���UD�n��l����uׁ�)    <;�  ,;a׮ܱ��)?<��B>v  p�4iر�1����NYYʃ���������W��NwXj��'�6|j�=����)    �>w  ����^�)7:zk25���-  ��Q{����_�#�p�D�9R*>\*<XJ
��	`-H�4����}��e�}}'c�    p�� X6��6�J
���-  ��Su�%�կ~um����P(�)e�����,v��WW7�l�������N   ��� ]������dd��$ר  ��Ttu�k���u�;������������ҡC��Tr�;�"�\!tv~~�=���   ��x ��ƶo~ax������b�   �$�Kv�lJ+*<��A�,�KŃK��/���r�$��&mnޗ����s���-    �`^&  �Ж-�-�R�eձ[  ��U��7��6m��ݱB���hV<x��<X̆���A �EZS3�tt����w�    ���;  K�-[�+nIFG_�  XU�zUM�+^Q�c%
'Ndŧ�*eO<Q,9RJ�w8!M�i{{Ws�i_���    �w  �����W�����'On��  ,���<��v۶��+��|�t�P�t�`�x�`))B�$��*]��\s�{;��y2v    ��� �%3x�CC�HB��n  �Xee����oLr9ϥϖr9�JŃK��/��G�����j&�踩kϞ��-    �/  Xtl��x�����Ǐ�d�   ������\{{E�U*�������W,8P���� �*MC���ծ��Ҿ�,v   �Zg� ��:���򊑑?LN���  ���u���z�K�cw�剉�x�@���c��䤱;�)�����߾���c�    �e�  ,��-[�[��$�X  ����+k�l��ݱ�������D��������c�    �U�  �u_~y��,�������n  ����&mx��Ϧ������G�)cw�g��i�ut|yӽ�~<v   �Z�%  g�@O��������sb�   �O��߾.�ܜ�݁�;���kiy��a�{�����   ��� p����-;v�cI�T�  X�j/�����ϯ����T-��/(�'���VS3:;�?�_���)    k��;  g,��Q9x�����թkL  ���|��j~���bw��lh(+}�������0?bĖ���RG��ν�[b�    ��G  ������҉�?���.v  ��嚚r��xGc�NA�|�X������ŤX4vֶ����jk{��}}'c�    �f�  <kǮ������'C���  X9��ƴ�>��SB��S������Ť\��G]�P��㽝w��H�   ���� ��v���ﾛ����3�(  8-u��u�.�����fg��'�,���B6<���Xr�Ig�omܻ�K�S    V#w  N����\��ѣ�975���-  ��T�җV׼����;8s剉������03�Xw`�H�4���{�.�����P��   ��� p���__�l����  X��6�����u�;8�B64��{�Pؿ��
!v��hhx*�~��:��y2v
   �ja� �)غ��tp�!�*b�   +\�&�{_SZ]��*J��=�d���c���å��`w`�����uv�j�]w��N   X�<  ��
o{[��c���]�  X=�o�ϟw^e�W��+��/y�P���tV�4-����l����]��   p� ������Eax��07��  X]�_��W��6vK�<:Z*~�ۅ£��R)��Xis�RG�;�����   �R� ��zz�%ǎ}2)��b�   �O~Ӧ��7��!vK/,,��'
�}�
��p��l����6���/�b_�   ���� �c��+>��ޓ����  �Ni>�4|�MI.�9�V��Ȋ��������S݁գ�b���y�y{��;   `���  ��{����7��99~��[  �կ�-oi�wvV��`(�Cv�`���#���å$غ�@�����wν�~$v
   �Jb� @�$Irt��Ӊ�?Kgg7�n  ֆ�׼���e/���������w�[,~�;�0=]��p����׶��������-    +��;  �PwwOyp�SI�X�  X;*~��*k{z܇��B�C�J�o�P:x���m݁�+��N���ݹ{��c�    ,w�  k��W|4zw!�  X[������oL<��Gss������C����TQq2�����={�b�    ,g^  �Q_~y}{�pkU�  `�����ZZ|p˩)�Cv�`���#���å$��E �'Mˡ��+��{�Gb�    ,W�  kБ������tv���-  ��V{�e�]T����<9�{�P|��BXX�tV�t���u�������-    ˍ�; �3��}Y������  ���ϯ�������\�Xف�·�Uț���    IDAT�Ʋ�= ���n����m�w?;   `91p XC�l�p:8��P.W�n  H�$I׭�5��]>��(���
?\(��_��;�TV�:;?�yϞ=�S    �w �5 ��V��.�"v  ��V��w5�֭���`�'O���=V(<�p!LO�c� �0i�fiWןt�sϧb�    ,�  ���k�ݔ�Rr����[   �I�-u^X��U(��>\*|�[�ÇKI�� ~�����jk{��}}'c�    �d� ��ݲ卹���&�Bc�  ���⋫�������n�����C�G-�,������ׯ{Ǟ=O�N   ��� `�:r���PȲ��-   ?L�ښo��u�;X��|��装�C��= �FU�L��M7��qǽ�S    b0p XeBoo~`|�������n  8%i�4��ј���b����ˡt�@���o.dcc�t��4�+�:;o9��{n��   ��� V��mۚ����<LN�0v  �騽�����ϯ���ڔ�
���B��'�I�s �$I�4MChk���5�ٙ���/N    k��; �*q�������/%ss��[   NW�O�Du�O�Tm�ֶ05���+��+$���;�,������_�ʻ�   �� V�����'CC��º�-   �F�ƍ���^�4,a~�\|��Bᡇ
��	�&х��c����:���n   Xl�  +�ѭ[ߟ���e�[   ��4�Ov�lJ�yϭY>��P:p�X��7���,v������\g����ob�    ,&/
  V���_��th��u  �
����6��9�ǻ,K�G��\(>�T)	!v�F��|1���[�{��Y�   ��b ����[�yt��&��/��  p�T_ziM��_^�~���xVx����c��r9v��iH:;���/���b�    ,w ��k���-����  �l�ؼ����kbw��(�8Q.>��Ba߾BR*9�Xz���u���#��+�N   8�� V�����%�÷&��-�[   κ��t�Ν�I�zv͊��˅}�
�\����J��n����ݻGb�    �-^  �#==o.=��$˪c�   ,�����!�aCE�8]�X�����}!�̔c� kHm�hn��wv�����)    g��; �
0t�7f��;�r�[   S��P[u��>�e�*�C�����̗''݁�QQq�t�9�z^��S    Δ�; �2v�|�?HFG���  �*/���f˖��p��q�>��o,��ǳ�9�ꗦi6n��ƻ��l�   �3a� �L��m��y25���-   K%��K������kV��:T*|���Cw`Q�iB[۽]�y��t�.E   X��   X��n�zan|��&ss��[   �Z�;ޱ.mj��-;v�T��7�K��b� �[�ܼ�P}�u������-    ��� `�ٺ�����g�b�>v  @5W\QW���U���R.-|��'�(�nV�P_,��v]g���-    ��� `9v��!7<��\���  K�EU�\vY]�Xl���bKkj�r]];;���-    ��� `�8z��H���K]�  k\��9W���7�R*-|�����\!ٸ���ٻ���-    �";  `��v�v��OFF�5n  H�0?�.��*��t�Ě�64�*/���r��0?���M�ꑆ�ϝ8�_�������{    ~/  "z�������NL�8v  �rR��]�������݁Ő�i��_��W��[    ~w �H��vV;���33ω�  ��T����5�}mm����X6�MWK˻Ӿ�,v
   �3��  X��tw?�jh�+���9�[   ��4��򢋪cw@LiCC����*7o���<1Q���ss�g�����[�����9    ��� �ر��������C��.v  ����%;v4��՞c�?ʆ�J'�gK}��rW�����ۏ�N   ��  XB�W]�~3�2�  �u�^[�?������d����ώ+�nV�P[{�z����v�~,v   ��� ���֭�O���$�|�  ����'���������U�����������p�X�*+g����o����N   H�$1� XG/������$��n  X)�\.�|��bw�r�66�+/���bÆ|62�����	X�������_|�ˎ���Gb�    8� `�;*��x��0:���-   +NEE�n���$��,~�r9���/���B��)��V�4M���s�S�޽��n   �6/  �×_^�6?��tr�ű[   V�����!��Y�V�P*��}��}!,,8�8-i�����Ս�W?�   X�� �S�^�U=<��ω�  ��U���5U/}iM�Xq�>�Px��BR*��%mm��ζ�w�}}Y�   `���  Xm��o�(70З��v�n  X�Ҋ�����bw��SQ�V�{ne�_X��J!͒`����'7�f�O���w����-��   �'� �E#۷��t���B�!v  �j��Ԥ�{_c�y6����dVx�����݁S�독���l�����[   ��� ��d����ţG3�2'  �E�o{ۺ\K��H
gAyd��p�}�C�J�[��!��=^��|�s����-   ��`� pl�zC8v�i��-   �M�e��V\tQu�XM�#G��w���X�X�Ҫ�������=�   X��x p�����ñc�K�ĸ  `�����.����I��)_y��U������P�
!v��eYU��ܖ.����|7v   ��� ��c�_�����u���  �h��|�z�K��g_�kk�W^|qUZS�f��YR.�n��*r��?�/{��g�;   X�� ���kWnG>k:2��  `�+B�EU�UU>.�E��ri�����/�JJ����d���e*�\z���>������'�;   X�� NSر�r�������&v  �ZQ�ٙϵ�z��(��J+�?����~�"LN���ӎs�I��w��u]灦��g�&� 1H��8�3�X�5q Ip��Dr�T�+�S݊ɝ�z�0�VwUuD٩NuW�R�Tű%C2)S�%��Xq�x��XII  A ĝ�9g��.ٚ8 �wx��Z������|�;2�����ͱS���6     ��n   n�O��-�d���L�    @%q���w_�tPI�˗�o}+LM1���-Z�R�_��o��      �w  �4��Uo���zf��-    Pi��+���T�� *Nh���|���.��im:@Z��[������I^�     ��w  �p���fgd�Y�J-1�    IJQ}�D�����"�rA�G?�~�Ü�}�5 �LP_�K-zDvw�M�     ��g�   (v���r�ge:�d�    *���j��:�l[�K�:Κ5��dt01��f ?'3����?��5k�����=     ����  �]�~������n��,2�    �Ώ�=�@����Vx��X�C��-� ?����/N��vu՛n     �M�   (V�zЉ��/�yQ�-     !��;��Ue���i�B�[���lV��Pt,Z[��vw�n     ���   o�Jg�Qgx��f�    �G0:�	�g�(�^�ƭ�g���ݺ5$�� !S�u����2�     J7�   �dh���p��2�    �o��t�7����B*t�=���W[--�� ��L�A%ώ=��t     (=�  ������+GF~_c   ��##�� o�jh��]]����Q�I�= ̒�|�78��cǎ�m�     ��t   @�ٷ�##�B�     -��p��5��I��`9�ׇD���Z�n`J���́'�o�?���g:     ��  ��{���"�xT
�v1    (bA:�C۷����߀"&m[��펳f�����`j*0��� �e2���[�^�Lo�k�s     @�c�  T4}�:aY*��:M�     n��{�JWE�|}(2VΝw�vs������X�T"�-53s�۶͜���G�9     ��1�  *���FΝ�y��L�     n�Z�Ȳm� n�����M�\aY2�f��@J�����֭����     ŋw  P�tW�5z������n�-    ���\W�+W��; �$���d���y�����`j*0�`�I�L����nu������     P�p  G�8�~A_���t    ���lV�[��Mw �52R��5��x�双�"�g�;PY�H&w<�ys����M�     ��À;  �(��	'q���brr��    �-*��n�#C!e:��SX�ƍ��R�##��̹D�Tj�[�ԝ��c�     �� @�Џ=y�/���ͦ[     ��jl�UCw�@��JI{�R�Y�����~�L2�T)��͟�뮆�����t     (\� ��𝮮��������`�    p�d$"�+� f��F��~�k��(oh��o:	���2���M�ZO]��u�1     �8��V  P�~�wolY"qZOM�7�    ���g������u�����jg�j^`*����޽�1�     ��  ��]��]�N?/���4�    �=��d����t��'�Q��E��ɚ�e�K$��|��5�     ��R  ��ɣG�r��i}��J�-    ��$lqʘ���T}����Ν!�x�T���}�     n @Y�<z�.36vF�̬0�    ���o���,ڽ;{�j���2�`���~���h:     �À;  (;�c��GG�"��e�[     sǏ���T�p�����"{�D��J�= ��3|����'O�<    �
�   (+�c�����J��n    �1�D��>V+��n���t:�}�;����M� �c~����Q���W[     � ��  ��@WW�?2�<��    P!�@�[܁
#�Q~�h��3*c1^p���į$��?���,�)     `�0�  �B���v�ʕ�2�n6�    �?^<�FW�BY+V��G�q7mrM� �;�ڵݣ��ݺ����     T� @�=xp���xNf2�L�     �W����`2����F��ɚ�{e*�vmk|l�!w     *}  ���;;���ǟ��L��    ����q_�6��,��͉���W��6�BJ�9 怜��+1:��~챐�     0�,�   ���#�D�"�]`�    `Hg�
GVU���pҲ��|�c���~<��l��_�r��6&�����]���o�     ��  �$�;�ڎ�?/��:�-     ��x�7� �xX��v�#�vw���(C�����v��    ��ŀ;  (9����^<���1�    ~<�W �Ȳdh��H���R��<ʌ��ڐx�guW�k�     �>.�  @I�8�=�3���[     ����t�⣚���#��t���PN������h�>q�1�     f7y  �d�;;���ĳ��v    ���lV���� E�M����� �GNM�5���y����m     ��  �$$�[,�ǿ(2�E�[     �'�L7 (n��Ѯz䑪�=����,,P6�]��z����I�}    P&8� ���8vl��H��t��    @q�}� J�R�ݺ5��_���rʄ��ؕx����!w     �w  ��]������J-1�    (^:���-!� J��F��a�+��Ȉ/�6��ve2�f��7>50��     p{x�  �ɣG�f._~��v    �{�ׯA2�� PB���ݻ#���*UW�33�ȫWH<��4�     n�u  �(]��͌����d��    @iFF<� J�jj���<R�n��np����=�={��t     �u� ���ݎ��\<~Z$��L�     J��3���HǑ���F��ɪ*���nt�H����2�     nt  ��|��+�4���33+L�     J�?4�n Pڬ�6'���T�+W:�[ ܦ���=�3     ��c�  ��tuE�%�����-    ���OL�"�Lw (m2V��c�C��2��{ �:kl�ktϞc�     �� @QЏ=Z>:������t    �Di-�D�-� f�u�n�#���.�M� �u��د����/Mw     �g�   �'N8�7��SSM�     J���Q�ҥ�� �A�B�Y�֑��
�\�֦� �<)S�͏o�R}���oL�     ��ƀ;  0J�8��/\xFNNn1� 7E)�l�RѨ
&'�9   �9�[皎 PV���h�+W:�訯S)�܁�#��̖Om�b=�����c     ��c�  ��������brr�� �Vc���9�օ�+`���4   � ����CBJi:@y���r֭s�eI?g�;Pb�R&�;?�m�~���{�{     �;c�  �O�T�s� �]�i� n��d���x "��,!���%�����(L'  @ka/[��je:@�R�K��βe�?8��\�)w��H=3���[��������     ��p  F��e���z�n� pC����n��ᘽd����@e($���;>�?   �Ԃ�ji�Mw (_��J9k׺:���W�= n����߶m�To�+�c     �[1�  �]|Ϟ?cc�Mw ��P��*z�@�ټ9,m[��?W]�dM����Y�  `��,a�Y�� PޤmK{�J�Z�@y�/{"`�(!J&��>�cǕS==�M�     �_Ā;  �W#����H$~�t �'ۖ�]����QY[{Cg'����\�'�\�  ���m���/� �\P��j���N���P*�V:�|��۷��ٞ��9     �a�  ̛xG�'t<�1) ���z�9|8�,_���P���f��LO��  ��ΪU��F�� �A���Y���'x�(Rk�J��~b۶|��g�t     �).� ��9p����2���ɪ*�쌆;:b�����KJ�ȁQUW�y  � /�L7 �0J��=�D�ǎ�d,�P*
���H���G��3�     ~��5  0�F����Bk��8I)܍]��#�qf�LM�駟N�\���  �Y��� P�t&d����w�/� �"�T��ǛΞ0�    @�c�  ̩xg�^=8��2\�- �v��+��C��h�����gΤD��  �� c1Y���y�� M�_}5����}�- n��FGessg���c�[     �d�t   (_��&��?�p;��d��ݽ;}�᪹nBk�R't�����  ��t*���� L��ƍ��?\���x&� �N7cc��G�+0     d�   �)��y�=:���P�2� ��^�Ԏ9s��R�闭��f[��A06�p  �<�/�UC�� ����r֯wu*���qΆ@���$���ܵ���x���     ��  0�❝mbt��:��1� o&�aٳ'9~<����m�)|�}����*  �y���� B�82�gO4�T8Μ�h`LO�M��}Awuq�    �� ��J;�X��~Id2�L� ��9�׻�Çc���B��0���^��)��D>����  P�<O�w�2� ?�,w�j��u:��(f�lKJ�ͧΘN    �Ұ�  ̚k]]�zl�[��M�[ �gdU��9?�PT����@2U�Çc¶��  0O���@g��� x3Y[kE~��ٸ�5������������     *� ��Џ=���=-ff�0� B!��Mn��3f-\XgU;v�    IDAT�*��Az{�[   *���b����  ��?}��Z�@y�.y"�]�h�Rw~z��EO���t
     ��K}  p�tW���x�Y1=��t !���U�C�bΦM!iYE�1]-X`	��?<�n  ���Z�mm�� x;���rV�r��!_d2�t�w�Jm���͡�����t
     ��w  p[�ɓj�ܹωk�v�n��mmwv�T]]ўw��VKOM��+�   �B8�ׇLw �;���r֮u��L\��9(NR�R�?�m[���0    @�+ځ  P~ǲ���z�~� ���T��ᘳqcH*UT[�߆��-s��O��l�  �CA:��m�J�7"�
&-K�+W�VM��/_���!)gfv?�m����s�c     (g�t   (]�={������ P��Ν�أ�V[�Ͷ�%m[���h�A+  ��B'�� ���u���j����P�����ȿ�z��C�S     (glp  �dh߾�Y�����������ъ=Z�^�
)K�G2�VK��?�g;  �ܑѨ���l�@	���r���׮���T`��/�Z[~*���۷�3==q�=     �#.� �Mڿ�7������$����}{(�kWX(U�����|楗Ҧ;   ʙ��QΝw:�u���e��R�󯾚Ͽ�rF��� �D�n�]����ӧ{L�     PnJ~  ̯xg�^=8��e8�[ T&�p�ݷ/�-�M�̦���M����Lw   T��ɲ׭s�U���6��揌x��~5��I��EFG"�VK���ӧ�L�     PNp  7l��������E�5��I)�-[B����,�����:{�l�00��N  �Ҳ��l��]�X˗;e�;@Y��l�}饴w�gF��TW\ji9�+���)     �.� �:~�����f�M� �<��V���Z��e���-r� ��3�`r��|   �L���^��u֭s���t ���:���fs?�ANhm������5�w߇�ɓ��     0��  ��ZWW����L�� FJ�n��;;c�����/�-��v�;� |�t  @e�<$~��W󅾾��<m-X��m�(@q�RZK�:Vc��_��qn���d�SW��qj`૦[     (\� �w�O�p��?���֙nPYdM����Q�������gΤD��/   ��e	{�J�ݰ�U����N@�����/���S�@�--���`�    �RW� �m�����,�]�n�@eq֬q���d}�m��U[k�PH��/{�[   *��"��
��
��t6��:K�B�0J���Y��&'���5ގ�E2���[��������     J��  ��<�п�cc�Mw �2���{�V{{�mm;ٿ��t���;   �&J	{�2�ݴɵ�����4����r��}/+�6�@!���%K>����|�t     ���w  �F::~O��� ��^�����Ѩ2�R4�@gΜIy��lr  (B��Z96��M�������B�k_K�\�)w��v�[��mg���t
     ��w  ������W���К�� �m�н��ݍ]�孲� ����`z�O�  )iY�^��q7lpUk+[������ٳi=1�n ���Tc㱦�gL�     Pj�d  ���#�\���;�[ �?���
�������bLL��g�I�B�M|   EN��+g�z�]���/��W�Pйo|#]��)�n ��FG��K.��f�    �R;  ���~p���ӢP��nP����Ю]a���]�Xȼ�BJhf�  J��Jg�z�ݴ�Uuu��	`>��������Yΐ�y����������Λn    �Tp�  �B?�*����|�� �M�֪ȑ#1g�ڐ�����,�����L�   ���	���+�`d�S��TuuJ�x�ܓ��%���ly��}�=@E���;N]����     J�  @|����mj�"�j5���9�׻���H��,rkt���҅����<  @	R(g˖��v��ob �A_��gΞM�W�2����x����O��     ��� �
�O�p쑑g���J�- ʗ�Fe�����ukX*� ϭ�ֲe�劧S)�3  Pbt6������+y��h�p�%]��� ����n�����`b"0�T2�N����͡�����t     Ŏw  *�����L_���t��e���ѣG��ŋm�-�@*%�+�BOOA���  �"��Ȉ��J.���UM����2��<I���j�#����g��`R�R۟ض�����4    @1c3  ,�g����#�; �)���kW8�cGHH��c����~�٤���<  @9��,�C;v���v[pw`������/f����4`��,O��>�|���L�     P��$ �B�vt<����֚� f���Q���������9�]��ϼ�b�t   f�Z�@9[�����]�gv �.����_�rJ_��n*��Tk�5=����S     (F\� P��<���>���L� (?���N��""R�[*A�o�6���s�;   0�d,&�M�B�]w�d(�]>�Y��� s�l�O$�,`��D&dKKG���c�[     (6\� PaG�l���(
��� eƶe��{��ƍ!�)FgΞM{/L�   `��t7lpݭ[C2�%R �'t��HΝ�<	"kj��������     �	[[ � �~�!;8����jM� (/VS�;~<f��9�[*��W�p��O���t   f��d�/��'9��j�B��� f��Ҿ�G!�x�3�T�\�>���S�.=g:    �b;  B?�Xh���3"�j5���H)ܭ[C����2a��!Ҳ��|�]8w� <f   ʒ��O$|�Wr��끪�W2�78��%��V�Z�Py��=@��d�>�eK���M�     P,p �B�N,�����f� ʇ�e��3�l�R�A�0
)���*\�P�E�   eKk����W^��㾪��T4ʠ;�ۢ��-����
�P0�T�dr��m�6�����h:    �b�
   �w��$��� P>��f+��S��������r��f�t   扔�^��	��R�ۦs �6�J�^H���o��4Z���|�o.>}�oM�     `�  ��������%���� n���ݲ%z���B)��R�r��V:����Mw   `I)��˝Ю]��-��t����^_�܁y&��i��x�����-     ��@
  el�ȑ_�\�s���� �O��2������-xA�3�?��\�L�   `����v����E�tp�t�������ﳦC�J�c�x������{�t     �0� @�=xpE0:����M� (}vs��舩�je�7(�R�<����)   0�no�ݻ�X�� �����g^z)#<O�n*���{���ʓ'��    T$.� (C��訩��|Nd��[ �8)��uk(�T����ۖv{�]8w� |�t   ����k���q�Z�В�(���U_o9mm�70P����rd���k��O]����     L`� �2�O�T���y��*�- J��e��3�l�R���$#e54X^OS   ,��
���ד���h��˫ n���RΪU�w����Y6��D��k߶M������     ��  ��a��^OL�c�@i�Z[����Uj�"�tn�Z����-�+W<�-   0+��򯼒��d�/����"+�"C!�^��$���C�����m������^�1     �'.� (#�>%��~�t���n��>���P��B��ٯ=]8w�M�   B!-K8�׻���a6��Q��t���^?�K`��v�Z��W�{��)     �V  (�VCC��Z� ��uet�ވu���́ Йg�Mz##��   Ǒ�-��}{X:� �7�u����~����R�Hd�ji�h:}z�t     ��j  �@�ȑ����3��[ �&U_�"��Ԃ�$S�t:��~:�gf�-   (.2����v7lp��<; �򯾚���_g�֦S���kjz[������     ��+  ���?ܐ��|�� ��Y�։>\�b1e�sK:��[[�¹s0�  �7)�?0�y����J��z%X��]X����h�*\��q�����H������M�     0�p ���.wrx��H���nP�������;*�bp�B�XLYuu���+�n  @�љ�.����AO��[���a�#�`�e/]j{���y�s��'���Ol�\s���e�-     �%� (a����_���f� J���V��Gc��U���?�p�%�@��o�   �)��х�_�W��vS�%C!��-U]��ի��eOg��tP�R��>�m��gz{_3�    �\aK#  %jd߾�GF~�t��c/]j�;:�2a@����/���~6�  �]I����nh���9G x{�l�~ᅴ?<�*w`�i����֏��=�]�-     �� (AC�����֚�� �qR�Ў!�}�)9@�BAg��Ť�*��  �d8,�;B���!�g
 o��:��250"�	����t����     f�  ���C�Vى�i��W�nPBGF��X+V��SP\��� ���3:��3�   �!j�~����wp� �VZ�췿�-���9�)@��uuo456v��n�     �
[_ (!��Gc���/�lv�� �C�թ�?Xe��8�[P|d($���;>/43�   xo:�Յ��B�Hx��Ŗ�D��& EDJi��;�u�?8���Z6�(i��.^|�t
     ��w  Jȉ�?'��ך� P:�����ѣ1Y]�o�#U]�dM���   ���tPx�ռ��	�K�6_��sVs�m��)���/TsG��k>�m[���0�    �la� ��ط�cc�; �)��sg(��CQa�lS�{�,��~"�'�  pS��q����y
Ik�bKHɠ; !�����-���A`:(WR$�;o׮>y� �     f��  ���>�����К!U ��qdt����b�k:%Fk�9s&�]��'�  pK��F+t�}���6��x�##^���S:�c�;0Gd8|M.Y�����1�-     �.� (r��Y�='
��� �O-X�"��T}=_k­����O'��)V�  ��H)�ի��#�����!��]��gΤ���M`�蚚ޖu��?����     nC/  ��vt��_������nP�����ȑ#U����:ۖ��e�w�|A���   ��`b"(��Z^h-��fKH�����HD9+W�ޥK��f�����-L�r+N|�t     ��w  ��>yRٽ�ψ����[ 9)������>����n����h�U�p�m_   �uA ��!���-�*YS�3	���PH9�W;�А�S)�܁9 3�U�ڼ�{����[     �U\& P�~�q�P\���� �MZ����u�+$�`��F��Y�q��g�   �Mg��p�|A��VK�ŋ�@e��#�;�t��q?��
L� eH�Lf�v���S.��    �V0� @>p�a�H<&V�.du��?����-(OVs��S� �M�   ����~����"�Vc�%�� *�TJ:�W;zj*&&rf�֖�f��]/<u��u�9     �,.� (2������2��x�--V�С��D���� Й�Kz�8C�   �5֒%v��"���E<@%�Z���L��W�S�r$kj��֭��'�-     �.� ("׏[荎>#���- ���v�9x0&]��v�=)��b�S��-�\N��  @y�33A���"��֒%�T��<@%�R�˗�B)�y�s�����'s�5�^0�    ��`� �"�O�TW_��L.7��HI)�ݻ��{�
�?0���Hk�R�p�\A|9   �DkᏌ��
V}�Ruu<� *���,�e8,�+Wrf��d�xb�V�T_��M�     p��, �H|̶�H^�v�� E�ue�����aC�t
*��F��Р
��|�   �+�Ӆ����u�Z�Ė���@���l��N����0��L�v~z��ן��0    ��`� �"0|���GF~K
�\ o���T���*���6݂ʦ,����f�   f]p�jPx����F�Z���P�TC�e56Z^o/C��l�Z�L��Ƿm�ʩ��i�9     ���  0l�С����_�g+3������ȁQ
)�-�?љ�|%�����   s�^��=�@TUWs*�?<쥟>%
�܁Y$��/6�����y�-     �6� `P�ر�2�xF
U�[ g�7�T8(&�^���<�N3h   �9LM�W_�K�VS�%�daPATM��[[�BooA����|��f�Z�����M�     �np �}�J�;��L��nPd������=�D�@1�JIk�rǻp!/
,r  �	�_��������b�H���
�����l�������ʆL�W<�m�>���=�-     �� 0���kq�ꃦ; iY"��u7n�nލ���d��?��E�   �;zf&�^{-/,KX��ls*��Ŕ�|����x��=2����;~�TOϐ�     ���  0���!�\�c�5/��9YU����Q�x�m��Q�����K/�Mw   �2X�Y�}��j�B�T�
LM��/})�gf�-@وD��mm�wwO�N    ��q �<�8�.FG�\�~�t��a54X��ǫT}=��QRTC���y$��   �?�Nk����¶����6w�B�pX�+W:�ŋ���1`6x^,�zד�.=c:    �_��  �HwuY���n�N7�nP<�e�����U*U�[�[a���zl���ؤ  �����\��A�Z�Ė�0g)��PH�+W:��K��2����4r���S���6�    ��1� �<:�����ڵ��� P<�M���}Qi�lD�R�˖�^?C   �7�̌�^{�m�@��+�ի��eO�Ӝ?�Y S�͟ޱ��'{zL�     �3\� 0OF;;�._�W���B�D��"�ƍ!�)�l	�����O'�\<   ���bG����Z� � �2�?��FF|�)@Yp�����K���M�      v  ̋�ǎ��_��%�y�- �������Q���1��6p��>s&%��t
   *�m�н��ݍ]�����\Ng����{�[��P[{���ȓ'��    �&  �~��tOϳ"�[h��y2��c�bVk+��(K��֒���/_f�    �+�?0������fK�a�(cҶ��f������4�����f�]kz���o�N    �w  ��oUU�����h��y��N�>��*��`�n���d�L&�GG�T<   �]05.\�[Z���� @�JIgժ��OM1��&�N�{|��˧zzΛn    T6.v �C#��}�t ��+r�x����78*���n##~p�:   ���(�?_��d`���R)���J)�^�A09��=R���~b۶�����    @��B �9r��s�58��2\�- �rV�v�{�F�e��Eg2A�駓�!w   �jkUd���jj�kZ@9���W�^�t
P�.5/Y�Wvw�M�     *�# ��G�����ݲP�6��,w��P��#�m��@�q���fΝ+��w   ��s9]8w./�vK�%��|�#)��r%�܁ِ��%-�S/~�t
    �21� ��DS�����J� �R��w�C��+���P�d4���-���z   0Gk�y��o����u9��蟆����LM1���N�||۶ԩ���n    T� �e#����;h��9ҲD��#�n�2��`�%��Аg�   �M_���C    IDATxo��WuuJ���(GRJ{�*6��O�Tjקw�z���L�     *��  ̢xg�^9<��!�� f�pXF������-@1��,���dLL0\    �|_x���Lv{�-�b�;Pn�i�;C��m�����]7~�O��r�s     ��w  f�@WW�58�_��GL� 0CVU����U��Ŷ��I{�
ǿr��ɤ6   ��~��߳[[m��� (7���P���6<50p�t
    �r0� �,�]]Vfd�9�N/1��U_���P����76�N����N��� �y��  `^&�o�Q����yY(7��B���oۦN�����    @e`#	  � 15�o���Mw 0�nn��]]U������{�Ѩ�<��   �Hx��}��׾���@�QJF��+V8�S�R&GF~g�Сݦ;     ���  n��ѣ{�ß�BH�- ���n��������UUJ��*���`�   ��`b"���
Vk���Q�x@9�R:�V9�ؘLM�"p+��D>߇7mz�O��r�s     �w  nC�ر�~<���"�[ �?g�:7�����.�MR��<폌��[   ���٬��x#/"i56ڦ{ �")��z�\�����@z^�:�����i�-    ��ƀ;  �ᓍ���d�� ��ݺ5�������v��mmv0>�`   �������L`���R)�}@���&w�܁[&���Ol��}�����[     �w  nQ|���U��0�`�I)B����}!C�����?0��tZ��   �,����Z�Ԗ��2�`��l�}l���rn��d���]����[  ��ٻ�8�����k�}�[7[2�dI�d0&��l|� _t�`
�&iZrNZ�6��4�$GI?INOj�i{.=9-m� �)���KJBp�M��E�-K��sifϞ�{�u^�$�o��ѳg����|~oF�k��� ���, ��c�w�7�?�8ϒ$��uW�|�u��)�/�R)���[��UF  �9��h:�яNw�|r>tp%I\۽�Qܴ�:�4��GG�����/�N  �?�� g(���c�>��ϯ��G�b\߳�Q|��ˡS��ĕJR���B���;Qn�;  =&ˢ�Ov���x��(I΄~�$q���K�i~�M�p���WMw:��w��C�S   �?���ϫW8?y�Bw �Q�7��6m��H�re!����ȑn�  x!��H�=�-\zi)�T�C?H��x�e���g�y���5��|f�?��7����'��  ��b� ��Ў?k6�v�����ո���7�����+\|q1j����LC�  �ɧ���c��.����\��X�K�yM�����hv֐;��8��ݾ��z�~���>�  ���� ��b���˳f�Cw �O�lYRX�\|q1t,����Vܸ��  =+o���'?93��#�(��B?�V�ƽ�6�/���P<?�,������~   8gl�Ӑ������B� �G�re�x�;ɪU~3���qi˖b�СN�n �7�y�=��FG��-��P�C'�L\*���.+u�Dss�G��sskf&'��w��WB�   �����pb|���N���8?�ի���e���!�j5���ۈ�eCB  ���C���>v*��LC� �\�lYҸ��F�l�o�p���~�����Bg   �����qbϞ�������QX�����hč���Pr������(6� @o��ǳ��~t�{�H't���+V�4�j�)��<�剉��V�n  `� ^����c��c��VC� ��qc�����R1�= ���B\,F�ѣ��-  ��4�>�D'ʲ��qc1�"����ŵZRܲ��}�N��H
�+�v��8~�}G����-   ,n��E�&�o}��|ffC�`�_��RmϞF\,B�RX���OMe��h�  ^Nz�x�OLd�-[Jq�x��E,�ד��s�WB����jm���^���SO}=t
   ��w x�/�Fccw�� ^鵯-նo�G���ŭ[Kٳ�v���<t  ��ll,K���l)ŕ��LXĒe˒Һu��Ot��#)���պ�g��������  �┄ �^t|��[������ ^�u�+U��p;��$���w7���=� �(���i�#9��8���2Ɇ�ھ}��`o��4�����>��*�S   X����0���th�cy��,t��ʯ}�z��(��C��K���aC���c�� `q�v�����+V$�5k|��E,Y��PX�&�<��M�p��Ng���٭<|���[   X|�P���������ׄ� V��kʕm�jQn�E"n4�ªUI���:�[  ��y�=t�u�yq�Ƣְx%\P(�Xwv3���������~��'�2t
   ��w ��;v�è�|g�`a�o��R��zd��d��B�eyz�D�  NW:8�f�fZܲ���Ea�J.���JQz��!w8q�I�}�?�����c���  ��a� ��Ğ=WD'N�z����-��)�xc�r�-����+n�X�FG�lb"�  �+���:G�tK�7�J%	���ºuŨ����A��t�i9Nӛ�;z��C�   �xp�(�������Q�}Q�`�Tn��Zyӛ����l)�G�t�V+  �mv6�|�;�����d�rC�H7m*�33y6<l�N���E?s�u���z�C�   �8xy
 Q�����ԩ��;��Q�o��o��:87�R)���ۈ��8t  �����g?���Ȯn�Z\���Zi����i������ׄ�   `q0���wlϞ�
##�
�,�8�jo{[�|�5��)���,_��v�l��� ���i�>�Pk���Q���$���v5
�\b�NC�e��������R�   z�)  ��|`�<=4��h~~e�`�qT��Z��C�JV�H�+��C��-  p��cǺ��t^ܼ�űۉ`�I��x�e���g�y��
�������ݵ<t��S   �m6���NL|(��Y�X ��a�(]qE�|�5��  p6:���O|b&j���-���+���o_#^��wW8I�y��۷��   ��y������]�����;�`����[�R+n��Zx  ��������O�SSi���ōFҸ��F�h��^F�����}�����  @�*� �&��_�7��%�vk�[�s�p;,Mq��n-v�z���ۮ� `��������ƍŸѰ���RI�6;�?މ22�K����t���#G�  @o��%ivj�����Bw ��vX�*���o_#�Tl� `Q�[�|�f�g��n�\�W���5�c�r��ѻN��yo�   z�w ��;w�'�9tp�n�(JV�*�v�G��]  �n7o����t����)��+\rI��}{=�����GQ�����w�{M�   z�� ,)��������o����-�9d���ʕ��T�ңG��[  ��y�=|��y^ܸ�:83Ʌ
�F�=r�s)��n��Ͳ7�맟�x�   z�w �����ߊZ���;�s(�����f��>�u���L���[  �l�Ǐ���LVܲ���A�b���U�(����qC�����?}�����|�OC�   �;����q|ǎ��''_�8��8��}w�x商ہ��~{��~���  ,j�o}k~���mEi��n�L妛����v�(�����ܵkk�   z�w ���.����~����v���W�H��$���w7���=� ��u�z�3��OLG�v�83�m�j�͛��;��u������3t   ��G~ �^>0P���(Mmx�>R��Z��]/)�Ւ�޽��X�C�  �+�=q"����g��iC$I\ݹ�Q��"7��K��z����,t   ���; }����/G�Nm	��;��n�����p;pZ
k��;vԢ،;  �[>6��x`:��LC� �/.������x�
�f�%d��ox��kBw   ��( ��c�w��� Νʛ�\-_w]5t���n-�o�ѿ  ,z�ɓY����QC��zR߷�W*N_Ë���������_
�  @X���o��@e���>w:+B� �F�曫�n0�
����|r2��Ʋ�-  ��t:Q�;��֭+�+V���D\�%��������<t������:��?x��B�   �� ���o��ĭֺ���Q���J��e���+w�Y/�Yc  �ů��[���L���N���֯/V﹧��ËI���qd��m�;   �G} �����{�E�����]W��v[-t���I�l)u|>� `�����S��ʕI� ',��Յ(���رn��QI)Mo�;?�C��  `	����gw��h����ө�n^���W��۶�"V�s$�T��%�����+� X��<�>܉k��p����9��)n�Pȧ��ld$�=��i4��-�>���)   �I�  8�.N�峳�Cw �\����;�0��s��k����  �<������o|�:8mq��;j�K/u0^�����}���  ��g�; }ex���i����aXX�J�_^��uW=�c���H.�������Аmy  ����n��yq��R��4�q\��Rz�H7o�\1�g��7�{�Ϳ����n�   �� �?���Fub�7�N��xe��7k;w6�$1�,��M�|x8�&'��-  p.�Ǐ���\Vܼ�Y=/.��e��:O>ى�����t��ō�>�P�   Ο$t  �+k������5�;�W��iS��g��v����z�=��< �7�����/}i6�"ò�čFR߿�W*އ��slǎ;Bg   p���@_ܽ{[wdd{���)�[W���m�8�*���w�A  ������|�󟟍�ܐ;,Ʌj�vգ��[x�<O
�����)   ��� �J��顡ߎ:��[��WX��P��q��+p���jR���B���;��  �D62��'Ofŭ[KQ;�	=.Y��PX�,�>��=��Y65;����|�   ��! ����_�[���;����Z��hD��ߧ@0��K�7���  Υ�c�uf?�V�eNr�"P���J��km��Py{s߾[Bw   ����ݻ�-������ً�/Ojo���^���|���__�  �R��!CTo��Zܼ��zM�������)t   �:  �V>0P����Y�8;q���wY�r�ߥ@�(^zi1L��'��-  p�dY6<��.���q�x	q/���9��[-S�{ĝΊ����>���-   ,[2X��&'%n�օ� �N\�ĵ�%\`��-IWw��+Vxf ��t�~�;���36�C�K���wo=�VH�P}����ׄ�   `��X������7���Bw g�X����7
k�nzR\�%�={Q�d�  ��b��x��Bm��F\�
�W���tx�C����   ���! ,:��@afx�������-������wo�p�%��- /%�ד��Յ�OvB�  ���MNf��pZ���R�uBK�/O�+��C�M�{�ϯ���\~ߡC_	�  ���D3 �Ή��_���7�� �BG�;�6m2�,
ŭ[K�n���  �s�������?m�;,�+�(�����zM�l��yｯ�  ��g��E�]��OFF��8;��n�������LTn��R��
s  �;�#G��"Q��jq�VϦ�=�,+eCC�4�   �g
� �t��ّ���ss�n�\��+�n�X���-����n>=m� ���MNf��HZ|�kJQǡ{��qq��Rz�H7o�<��_���`����}O=���S   8w�d`�<y��O��4tp�JW^Y��|��v`�*�ڞ=�x�2��  ��Α#����^+�sC����R)���S��U�Q�{�CCw����Cw   p��0��0t��U���Cw g�x�e����V��ȇ7`Q�����kW=.� ���y�N����C��W�(���mx6�����:  �sǛ z^~�`2��o�v�n_�83�����{Q�n�B�lY��\�t�z��  εll,˧���֭��Au�Y���I�bE�=tȳ)|W<7�槯�.�逸�8t   ��w zޏW��"�3tpf
k��4�RɭA@_I֬)D�n���[  �\�FF�|~>*^zi)t��
k��Nǳ)|���k~��o�̿~���)   �2�� �i���_5�����d�ʤv�@#�T���R��[��͛��;  `!t}tn�k_����ʛ����W�[�O��P�   ^9G �����FiZ	����Z�k��7�z�oM��q\ݹ�QX���h  ��������7ڡ;���qm��z�j��p�]����w����   �2^v гN����xr��;�3P,Ƶ}�ɪU>���Jqm��z\�ơ[  `!�}����G5���RIj{�6�rٳ)|Wwx��&��_�  ��g���4>0��{��oD�n5tp��8���U/l�X
�p�ĕJR\���y��N��s  ��K���/���.*�n^X\�%�/L:O>�	�=!M+����9���)   ���I����{�nۮ�He۶Za��r���-ٰ�Tٶ��  D�G�_��l����C� /�p�e���X	��"������Bw   pv��s�xs::zW����o��R~��}@����WW�ox�C>  ��<��=�J�}�vh�a�[n���lq�DQ�yR����|`���   ���9 zJ>0P898�[�����H����T���ZEq�����6���4;y2�  �\�G�'��7m*&˖Y��).n�\�>�T'o���1Z�鬘.�k�:�?B�   pf�����<�s�������)l�P��uW=2�EI�v�'�Vy� �?u���>5�ML��S�Q�$�={Q��}DQ��w�&t   g�Gw zFs׮��������x��B}��z�$>���j5���ۈ�e�6 З�v;o����d�N��zTrᅅ�]w�Bw@OH�Jiz�_��   ��p�gd�ӿ�i%t���e˒��}��R�{�$\P�m�^�b3�  ���ԩl����gg�C�*��5����{�Qe���5��y_�   N��$ z�;ߓOL�!tp�帾#Y��oI�Qܲ�T���j�  X(��d6�;�3����[�V���jq��b��ݡ����;V��   ��J �?ޱcE4:�OCw �!I�ڎ�d��B��^W���J�u�+��  ��������~v&�2C�Ћ�8��sO=^��7a��xnnե���  ���e �m������^�xy�m�j�͛k���z���u з�G�v۟�|+�"C�Ѓ�j5���ۈ��8t7:�����7��   ��p ��{�ޚ����xy�믯�����`QI���{w#^���7  }���t���ڡ;���^]��uW-t���y�01��zO  ��l� �|`�0�l�V<?o{;���֭��w֢8��	�ťR\ܰ��y�N�e�s  `A�'N�q�.���x�d��B>?�gCCi�j~~��ɓ���z�C�   ��L ����MOo������;v����䢋��� ������������������%�8��7�?zb��KCw   ����О=[������ ^Z�lYR۳����^��嗗�7�P	�  &ϣ��~��uC� / I�ڮ]���𮏥�ۭf��}�3   xq�"=y�CQ���^V.����q��7#�9R��j��J�;  `��i�~�3��x�x��VKj;v4��+?��d|���v�|g�   ^�7 �w'v�|O<1���KH���cG=Y��:����{�֬��+  }+���[���L>3��n��p�%��7VCw@h���?����F�   ��u :h>    IDATΫ?ޱcŊ���/NS/ϡ�Un��Vz�kˡ; �Q\(ą-[J����:��9  �0������n�+�q�ġs��Wܰ����Ԕ�(,]�nm:�6�w��C�S   �~6�p^m�t~5��[�xq�k���������%˗'�ݻq��s  �W�l�s���L��y��y�����x�rߋY�����G��!t   �� Λ�����GF��� ^\q��b���ܰ p֭+V�m���  ���9r�;����<_\�&�]��_���y^(ML�j�   ��w Λ��ؿ��ܛr�QɅ&����Q�6�<)^uU�|�5��  ����5�x��⋋�[o���%-?y���w����   �� ��w�|w<5������ո�wo#�T�>8�*��V+n�T�  i�K_�M�y��x���VJ�_^
�!%���h|``e�   �c�	��G�dt�gCw /"I�ڎ�x�J7, ��$qm��z�j�gt  �W�E��~������S��+w�QOV��\ʒ��ͭ�NM�  �s�� `�m����y�}a���U�m�6m��	 �J%���׈+�8t
  ,������O�䳳Y���ŕJ\۳���KY����=C\�   � ,��.�FG��� ^X骫�嫯���  ��U�
�]��Q�Q ����<������Di��n�_�zu��ַVCw@(y������   � ,����_���fh�A����o��� �o6n,Un��0  }-J�_�B+�"C��c�W]U)��u��d%SSW�ع�=�;   �:� ,��{��O��^�x�d���[�]9�c��]W-]uU9t  ,��w�ә��7�Bw �W��z�zu!t����t����    /& X��@yvp��y��,t�����w,K�/�[�G7o.fǎu�S�l� �o��>�-�Y�$^���8I����c�u�,��_�[?�n_��Ç�:  `����q|j���V�U�;��Q}��zr�>��$���w7���=� п�<j}�s���x:��|n.O����s�/|��~�V�e]�d�##���_�  `��C �N��yi48��(M]�=���7W��__���IGG����OGݮ�  �V�bE�x����ժ�p>��e��D����Y��f�f����Q��������җ�:  `)2��97t���gcco
�|��_]���U��XT�Ç�[��tˠ  ���aC�~�@#J�-��[�,I��f��i�����Y�.X�8ΣM�~b݃���-   K��� �S����9w��o��=%��¤�����T�	���k�s?<�  R��k+շ����<ϳ��,N���4{n���vZ^�z}h�ƍ��<��N  XJ�� ���@�ıc�d�zK\���}������7W��������-  �P:�>:W\�:)^ye%t��������4���neφ��yj�ιVk��'�YE�:  `)1��9s�{~.|��{�qT߿�Qش�:�W&�v����NGGM,  з�B!����
k�Z�Q峳Y6:��V����٧��(��Λb��^v��6>����)   K�w Ή#k+�)�t\!=�r�m��u�UCw pnd�Ne��}�T�j�d  �oōF�x���ǍF�Χ��ʲ����l���p���>7�_t�W�����p�  ��; �������󑑷�� �F���K�;��| }%��~��Ӯ� ��֯/�ｷ%����<ϳ��,N���4���ǻy��03��8��֭��-=���)   K��� �b�}�nI�~���<�Q	zDa͚B�]�Z�~����w�3?�{��
�  �t��[���H�����4����4m6Ӵ�L�n�0;,6˖]w����ݬ   ���� X�ґ�_1��#�V��޽u�� ��x����p�y�ѹ�-  �P:�>:Wxի
�+�(�n�ӑ�����D����Y��f�f����Qn���������'�(�w�S   ���' ^���;2;v�Bw ��Q}��FaӦR� X�����9��  %.���޵,��"K��)y��e##i��L���4M��)[��ߕ���-o����S   ��w �������#G�0��_�xN�[��n��� �<���f�:��0D @ߊW�H����ˢj�-��y�g��Y>>�v�Ʋlx8M�y�e-;,U�z�g��?:  ��p��}��w���� �Sܼ�Xۻ�ű�x KH69��>���|n�p  }�x��ھ}�{���,Ϧ��bN�f3M��4�v=o#�����{.�ԧ�:  �_y	�Y9�s������4-�nl2X��g��>�ə(�� ��U~ӛ���nrs�F���##i::�f##i�l���d�
8�<r�W����   �ʀ; gep۶����7�� �(.���޵,��b� �ѹ�?����  �`�8�8�(l�X
��ⒷZY62�v��4O���,K��bv���q��6����\�  �~d��3vl�g���(�m��P���Z�u����  �������_̇�  ��W�q�=�Y�,_��$ϗ�y69����iwl,ˆ��tp���Z&فs��8��{�<��  �s̖O �X<9�K�ۡ7����l���Rݶ��MLd�c��-  ��v;�{衙ڽ�.���"��,��lj�!���4m6Ӵ�L�n�0;p~��lh~��?E�o�N  �7^�pFN�������_�DQᢋ
�w�kYT(�M�_�gg���}l:?y��0  �V��*�[n���������lb"MGFҬ�L���4I�4�,u���ȪU���s��	�  �Olp����ğ��?6I���j\۳�n���jI}������OG��ͅ  ���?�ӹ�ڵ��֭��-�[y��e##i:6�f��Y�l���X�o��n�ZE�KE?:  ���ഝ�瞟�����8����5
�^�. /*=|x���O��  Я�J%n��������[8y����Y6>�u��4N���n�jy��Ba.}�������C�   �� ��g.,>�?�N����ʍ7V�7��
n ^�������v�  X(�u�
�w�cY�$�y��,˳��,N���4m6�tx8u��/�.��K~��,t  @�(� `qH&&���v��aC�|�M�� ,�o��i�;��n ���L�_�j����X�+��tt4KGF�ld�����i�e�� L2:��Ğ=׭��GB�   �� ��c;w^��c����qm��z�6�p���wֳ���th(  ���sō��-[J�[��������;1�e�f�5�i:6�F����Ғ�y!����(���n  ��� xY�۶}<c�X��8�8�(l��C- g,o����~t:���2 ��W�q�=�Y�,_��n�Wy��e##i��|n+��P7��1��=���|�wCw   ,v�xI��woˎ�p�T�����7�����+�>���<�� ��Tذ�X��n�{��,Ϧ��lx8M��Ӵ�L���4�t�����8���{�<h�   �+P @o�'&~�p;�Uܸ�X���J� �d��b����=�
�  !=v�;��:W��KNS�����X������h���e��P��X���̬���"���  `13���:�k׏��>��;`)�������.��u�kpN�}�������\�  Xq��wY�K,y�y�����iwb"˚�4k6�tl,�r��Υ�Z�Z������o΄n  X������G��ή�KVG���K�S �+�����wB�  �B��/O���=ˢju�.�[�,I��f����P7��1�p��_|�%���?�  �Xp���_����KY�[���`!�N>�_��t::��n ��P���RuǎF��ey65�e��i:<�fcci�l�y�m� �<I�7޳����n  X�\���8��g����⥗�7�P	�@�K���{w}�#�����  �w:O<�)n�4W��ʾy��w:y66����i:6���f�u�ԹU�^gY9o�FQd�  �Y0���'O�r���Bw�R7q��{��v X@�ʕ���Pi��ߜ�  a��_n7֯/&\P�r��V+�FG�td$����SSY�;�
�X䣣�5����O}�B�   ,6��>C��]�?��>�@ q��jI� �_��+� �[�n����k����eQ���"���ʲ����l>7��l���t��W(ϓt|��(�:  `�1�������<��F#��7��R���R� ������k��P�  B�l��_�z�|���o���<����z#���s���}# �jj�;w޻����o�S   ���V��7|���;��f�Da��B}`��7���������??�  LG�w�cYa����)�t�|r2��ǳ��[ٳ��n�:[
���Ɖ�������A�s   �&��k���_0���Jqm����v η�嗗��|����	 @����ϵ��}��T:��^��tb"KGFҬ�L�f3M���(��(�gf�=��GQ���-   ��* �(���v퍟}�߄��cG�x���� ,M�/~�������  �t���w�_��G�je��H�m6�lx8�FG�lj�F^ ^Z�6�nӦ��p�  �i���(��(������T����l����W^Y6� @����_Η�l).������y�MNf��p������X�?���mk�8s��NO ���N  X�5��y_��3�Cw�R�\pARٶ����+;u*��ַ� �$�~���u�q������w�y>1�f��Y:<���f�6�i��f�����~���-<0�  ��pX�������;`)����}{=.��- ,=y���?��\�ߘ�S�c �4��v����Z�M����H�6�i69�E�Yv V�n��r���DQ�/C�   �:�T Kܳ۷�d�ĉ�
�KQ�o�������%����}tn��G�m�   8�J���֭�\��S�S   z�� KX>0P|�	�KQi˖b��kʡ; XB���G��{�����1�   p�u:�٩�E�?�  �˒� �3x��?���Cw�R��q宻��t 8�n7���7���𩹇�3�   N<2��鷿}]�  �^f�;����}��=��L���W��z\�9h������c��}m.���B�    EQ�V�'O�|E?:  �WpX����~>��_�����P.n�\
�@K�y����Wf��	��    =&���k�֋?�á[   z�w�%h���W��<�?t,5ɪUI��[k�; �_��P��կ���ǻ�[    xaq���V��(���-   �(	 ����<�Q�[�KI\(D�;�q��n��d����>5=s��ӆ�   ���ۚ�����   ��w�%�Ğ=��g��ۄ-�_�o�&�z��^ �[�v6�'27��o�EY�   �Ӕ�y!��(�B�   ����V��,+�΀���~}�|�u�� ��4��y�}��>5��#��   ���76��%t  @��E`	yf߾��~��<t,%�R\���Z�.N �\��C�:�����IS�    �Y������EQ�;t
  @/��`	)MM�b�������\���W,�x`���O��   �|r��={v��   �%6�,G��!:z������.��T��r� �lz:���?nw��/�C�    � ��&���:  �W���D�����(����I�lYR���Z� �4��~���O���v   ����:uٱ�;��  �WtXF��3���2t,%�;�Eժ�Z ����g:��応�����y���   `���8?x�w  �(��� Xx�����y�����W��^Z
��Ⓧ���/y6=v��   ��'��Y����,����  �ӿ }nh��=��S��"^�"��v[-t �L���}�˭��|��v   ��)��|`��   4��\61�S�`Ɉ�v睵�Trc �+�>�x��0��Zy�    gg�4���nd�;  �����ǎ�ڵ7:ujK�X*J�\S)l�X
��␍�����}衖�v    �(�򉉿�<h�  X�lp�c���O����#Y�*��rK5t �/����~�=��o�EY:   ���Z���?��(��C�  �P���S�v�|g>=�9t,	qU﹧�q� zZ�}������͓�<b�   �����}[� ���w�>ON����T�o��RX���* ^T61�������رn�    z[�j�z�����á[   Bp��ݹ�������;`)�W�.T���j� zT���<�n��o�2�   �i�q[� ��ʦQ�>T�������ąBT۾�%I��ޓ?�m��ﷲ��,t    �K�j�y��E�
�  p�9��gN������)���<(�pC��fM!t���޽��Y�w޿�u�! PP!�B�A@��TZ�l�(ۖ��ֻ7me�N{ߏ:?�o�{,�� �L*��h4*2:�z9ه�ֵֵN�����-�������_��e�\;�}} #��-�_�z���-�v    N�`~�/]q  ��� &;�i��a��S��tS=v �e����:O?�	�/�   �Դ�����$I���N  XM� �ȶm$�]�&^���v��k�R��$ $I�$E�Yt�~�=��/�[    ��7�����  �2��
`�,.>;�A������  I�$a��������q;    �-Ͳ�ٱ�Obw   �&�,�	�����������n]�~��3�; �/4�����38xа   ���t�$���  �Z\p��c��� /M���|䴤TJc� Q�������M�v    VZ�e޶���   ��w�	ph��������IW���z��<?L�b~~����=:��   ��HJ����   ��w�	P^\���0�Jg�Y��r�L� "�������}Ӹ   �U�e�{�w  `J�@
0�^���'8�!vL�4Mf����RIc� ��\m   `T\q  ��� c.,,�M��t�-[����׋� ���v    FI���жm��  ��� �ء{��pz���!vL��]�*�o�u&v ��X\v��m�1l   `d�?�$�bw   �$��X9���B�&�̇>�&�V��L�0x��n���2n   `�Z�_ݱ��   +�w�1��Ν��WZ��ʩn�T�\rI5v ��h�����������-    �V���_'I�H�  ���;��*?�&�};���^O���kbw �:�?�Y����5��   y���#۷4v  �J1pC�}�c������0�f�c&=�4�J .t�!߻��~�v���    �G�����   +�h`��?���z;������ʕW�bw ���C����>���r/v    ���h\��Ν��  `%Tb pb����N8x�f�Eae��rR�Ї�$I�%�IU������}��OU    ��|~���$���   ��w�13h�?��J�Bj��:S:��r� VF1??l?�p��o�q;    c-]Z��Ў���   Xn� c�q�����?�&U��s˵�[�; X�����=�pk����-    p��$I+Y�cw   ,7w�1�<v�����VB�&3wݵ&)���) ,�����_�:_�j;�m   `b��o:�s�U�;   �S%v  �煻�^[���f�+��eK�t��� &��ȑA�_m�f���    �-�Tm��.I�O�n  X..���w��_�^���0��3�(�o�u&v �(���z    IDAT��w�������   �d����Gfg/��  �\��@x��j��0�&՚;�I��4v ˣh���#�d��~7O
�v    &[+i��w�;   ���;�8z��'y~v��D�K.��7l��� `y�?����ȑA�    X-a~�#Gw�>/v  �r0pűc�.vL��\N�wܱ&v � ��ݷ/o?�x�<��   �U5և���;  `9����gg?�������v��3���*�� �Ԅ,+ڏ>���>O�m;    �)���<�6v  ��2pq������ ��t�Y��7�cw pj�C����7��b�    @T��iG^���   ���`���cǝI�ui��D3��TJcw p�B�o�������,s�    �$I�(����Z  `����F�oC��̪�6U���Wcw prB��/})�}�{�$ض   ����uG�����   8� #굏}lsXZ�6vL�Z-��~��� ���ѣ��s�k^ye�    F���'c'   �
w�5���O������>��]�`^~��y�Vh���-    0�B�y�/�o��  �dw�����������&M���˵k���� �Ą� �O=�u����0v    ��Z��W�   N��;�*�����P��%M��}hM���`������o��~�    ai��C�����   8� #�q���&��w��IS���Z���+�; 8~�����=�p+;�l;    ��4I�R����   '��`�,���g���&J���o�u&v �-�~�����Y���1    0����[^۾���   '��`�|{nnMyaa[��4��n�IO;�s�8(������>�l��v    8Y!�r���  �Dz����CI��6vL���sʵk���� ���,+�_�b���˽�-    0	���]߹�w��   8� #�XX��� �f�w�$�R���7<zt�=�psx��0v    L��`�%!|:v  ��0p���~<�����IR��jy��j� ���嗻�Gi�,�[    `��{�؇   c�/0 #�����`�T*i����� �m���?�����	C��   `%��ιo��_�  ��e�0^���)i4.����~�-��gx�U�n�y��o_7v
    L����b7   /�/�Pi��&M�4vL�ҙg�j[��cw ������_h�n   �i�6W�2;{S�  ��a��/?����������~�k�R�K# #h��+���?�*���-    0-Bi��z(v  ��0p���l~6���0)*�\R�\rI5v �?����җ����1    0m����~�я�'v  �;1p�腻�^���$vL�R)���kbg ��Ð����'��    bH��:�j}&v  �;1p���4}(�����IQ��z��˱; �5y^�{,������)    0���an��  ���DTZZ�/vL�tf&�y���; ��B�1̾������A�     I�^�]���S�3   ގ�;@$���q_h�ϋ������$33�m FD��k����V��P�n    �������   ގ@,��'c'��(�[W�]}��������=�H���    ��B�y��ٻcw   �w���yUXZ�:vL��;�X��Ji� ������Od�``�    #*m6��   �V�"�6��1	��A��+�.���  	���t�~���v    e������m��  �1pXe�ssg&�����TJ����� S�(B��S�޾}��)    �;KC(�{��  �1pXey���d0�����z�u�Һu�� S��-ڏ=���~�    �������X�  �7���tq���0	ҙ�t����� �f��f_�Bkx�� v    p���5G^���   ���`ڶ���>/vL���7�$33�e ")^{m�}��b~���    ��tqq.����-  �H�K
�**�Z��� ��t晥��͵� �j��_��G�B�b�     ���y���}�c�3   ~��;�*9�s�Uai���0	��>��Ji��i�{��n�'�d00n   �	�O�n   �u� ���j�M�A.���{�S�\vY5v�4���y��;IQ�N    �IXZ����][bw   �w�U���w�Mo����v�mk�$���
���t�}6�    ,�4IҢ�|(v  ��0pX�T�"�����qW��j��+�; �J!��N�����N    VF�������   Hw�ձ����	0�J������� �*E�j�_|�;    XA����7����   Ib���^���&Y���0�j�^[+�}v9v��C��_��?�i?v
    ��J����   Ib���*ͦKp��մv�ͮ������c�e�_�r�    X%���C�����   � +���ܺ��xS�w��n��k�xnX!ϋΣ�����   ��I��S�   � VP��x(k�;`����^�n�Z��0�V�h���oc�     ����xs���ύ�  L7w�����=v���[o���J�`�������*��-    @a8���2v  0��V��;fC�}A�g���.U��ҷ  ��b~~�~��,4��    0����{c7   ���`��f�`���v�L����������/~�Z-�v     	��y�����  �^� +���܅aqqK�g�.(�7l��� �d�Ç�#�d!�C�    `t�f�S�  ��e��j���IB(��qV��f�$q�`��w{������    ���..n=87wa�  `:�,��gO�XZ�;v�����W)�_�z;�
<��<�x���)    �
EQ�6���  L'w�evd߾?y�.v����n��� 0���   ��1�����+  V�_D �Y�����0�*�]V-]pA%v�$2n    �W��ux߾�bw   ���`-�ڵ�XZ�*v��4M���z;�
0n    NT�����  ��1pXF�,�i>[�$U���V:�r��Ic�    ����t��;.��  L#L�e��j���]�;`\��rR���z��Ic�    ��J�<���  �t1pX&��Z�Hz��cw���l�\O�8��v�ed�    ��tq�#����;  ��a��LB����`lU*i���\oXF��    �r��G���  ��0pX��ڵ�h46��qU۲���Y�`��    ˩h4��   LC2�e�o6J�$��c�ZMk7��z;�2<�o��?���   �e�h\~t��kcg   ����}{nnM��p{�W��[k�̌g�e�/��d0�[    �ɑ&I�f�_��   ��1�)��v���`�&v��Z-�o��z;�20n    V�pa�07W��  L>w�ST,-}4v���֭���v�SV=:h����    ����׾�e;  �|e ���ݻ7���e�;`��zZߺՕ�ST;6l?�x�����    ���Zs�  ��g�p
���CIi�G�믯'��g�SP��ۏ<�
yn�    ����t��]bw   �ͨ�$�={J����;`��zZ��:��NAh4���ˌ�   �UB��e�g�  `��������a��g��qT��&��NA�j٣�f��*b�     ӥXZ�;����<  ����I�f��n�q��̤�͛�; �U����c��h�    �.���׾���;  ��e�p��]�,.^��Q���i���� K�n�y�Ѭ��7n    �ɲ?��   L.w���.-�e��ƍ�� �`8�/�=|��a�    `��o����;  ��d�pʍ�ݱ`ծ���v��Q!��lx�� v
    @Z�����   &��;�	:2;{wh�Ϗ�c�VKk�7�bg ���?�t���_�    #c��4�  �L� '�Ȳb7�8�m�ZO�u� '���o�����    �ץYv���[bw   ����|{nnMiq���0v�մ�e��� '���ۿ��    �j�?;  �<� '��,�D2���㦶eK-����p/���>�\�    ୔��n>X��  LC3��l �&-��ږ-�� �dx�@��u�b�     ��^��#��;  �,� ��ȶm�Fcc�7�뮫�����8��>h?�d;)��)     ��n��n   &���q*��!�܄���I���]o8N���<K�}��   ��P,,\wt���bw   ��P�8���ߋ� �z�t�Z� �!�y��җ��n�    �#�r��|*v  09� �á{��ph�Ϗ��$-�������� �aȿ��XX(b�     ������  �� ǡ��>��M��+k�3���NB��Of�#G��S     NJ�u�+��7��   &���;ss���ts�+i��n��;`�O?������     ���n"v  0����v����?-v����WKg�U��0�z�����^���     8U����ܜ�  �����FcW�7��w����^�����     ˢ�{��Ngw�  `��������[n6����r�ŕ���Wbw ���7�|���;    `�d�}�  ��g��6���?Ea�'�v�������,ڏ?�%��u;    0Q����s�=��  �7w���j�~�'�w��\^��K! o!��!���B��    'k����   ƛ�;�[8�m�šټ4v����7ד$Icw ����?�c6|��a�    ����Z��  ��f�����ϓ|N�q*�uV�|��� �*��7:�_�r�    `E--m:87wa�  `|n���ټ+v���M7Փ4u�����G���/�bw     ��B����g�;  ��e��[��kזR����0.ҵk��W�bw ��������vbw     ��V���	  ��2p�-Y���K�p�j�__O�e?3 ��XXv�|��E�    �U�f���;w^�  O� �Eh4~7v��Z-�^}u=v���v�Η���n7�N    XM!��Ȳ?��  �'w��ptǎ��N��0.j�^[K�u��~]�󕯴����   ���l�;  O� �a���Q��RR��Z��Q���7;��;     ��t�9�c�]�3  ��c��k��\9YZ�5v����W�3�(�� %��^��~��^�    ��  N��;��9���N{��cw���m�Z�� 0J��G�7�щ�    0
�KK���9ǒ  �b���Z���N�qQ~��*��ϯ�� ��.�O>��a�    ����z�����  �x1p��o�ͭ	����0.j�_�z;��(��?�DZ�"v
    �()e�#c  �	1p��K��O��`&v����g�*��;���J��ot���t;    �o(--���j�;  ��a��+����xp������4v�(��b��⋽�     #��_s�w  ��$I�ؽ��R�yu���LZ޴ɕ�$I��G�g����     e�NgW�  `|�$I��v?��J��뮫��������v�~�,��S     F�pqqkx����;  ��`��$Ih4�� � -����ͮ�E���?�C���)     �.kG���(v  0܁�wdv�������AeӦZz�i����}�|x�� v    ��(�Z;b7   ��@�z!���$��p\oH��/~�������     �$4���[�  }���K��ñ`����J��*�; b
KK��W��NB��    0V�pXI�?��  �>w`�ڶmch����Am��ہ���y�v��Y�    ��J��~�  `���m0x M�4v�����K���; b�~���ocw     ��F�ʅ]�Ί�  �6w`��Z�;c7�8�m�\KJ%/� S������܋�    0��pX����cw   ����Z��vm���bw��K��z�5�� �����3�tbw     L�f��	  �h3p�V���D�$.R�;�l�TK׬�� L�0�ΓOfa8��    0�ͫv�:+v  0��Հ��l�;�Am�f�ہ��}��v1?_��     �a8�tz�?��  �.w`*��}����Z�F]��ﭔ�;�� ��K/u����cw     L�4���   �.w`*z�O�I���QW۲��v`*����3��;     &R�q�®]g��   F��;0�J����`ԥ��^�l�P����B�:O<�%�A��    0��pX�v�s�;  ��d�L�׶o�4�Z��QW��ZR*��`�t��N��P��     �h����	  �h2p�N1>��`�o�TJ�W]U����?�I���˽�     �n��t�w��]�;  ��c�L�f��	0�*�^Z-�q��`��Fc����;�;     �AZ����\�  `��S���܅�պ$v����ͮ��%��?�T;��B�    �i�f��n   F��;0Uj���I>��m��:�T^���`5u�>92��    0U�k�ܜ�K  ��a�	L�a�uW�u�͛�I���; V��ȑAo��n�    ��3�β]�3  ��b�L����3�V���0��r9�^ye5v����󕯴���]    0������  �h1p�F�e����FYeӦZ:3�� ���uB�e�    IXZ�!����S  ���05J��ݱ`�ծ���`�^z�7�����     �j���o���o�  ��2p�B��g����ձ;`���=�\���r L��h;��f�    �$t��c7   ����
���gK��z�e�-[\o�C!�v���)     $I�l�?v  0:܁���l�� #�VK�7�S����wG�cw     �+y~�k;w~ v  0܁����I��%v��ڦMմZMcw ���o{��n�    �k�e��n   F��;0������kcw�(�^}�����+��}�v:�    0rZ-� �$I܁)P��{c7�(+�{n�t�y�� +-�ַ��oZ�    ��v��;w^;  ����xi�uc�e�͛]o&^q�P���ucw     ��jy~_�   >w`���kז���FUZ.'����; VR��C{��NB�     �F�e��  ����hE����0�*W\QK�u��D�>�l'4E�     �^�ټ��{�f  0�ڀ�Z��n�QV���Z���T:���R/v     �,�Pnt�s�;  ��܁��ˏ~�=!�.����t晥�{�[���RB��{�v�b�     p�J��]�  ��܁�Ui��OB�9o��ys-I�4v�J�~�[��h�;     8�Ƶanη �3�&V�ݾ3v��R)�n��?��5<x����{�;     8A����<�;  ����Hߞ�[S4��bw���\zi5=�4��D
�n����IB��    �I�d��;  L�J� ��pI��N�Cש�-Ԯ���0���=�	�f�    ���e7�N   �q��Hi����`T�kצ�.�0��G��/�ԋ�    �)�t�9�}��;  L)w`"�����`TU�����i�`��!߻����    �ST��?�  ����8������{W�U�M�j� VB�;�ɋ��"v     �.d�-�  �8܁����;FU��ʥu�ʱ; �[q�ذ��vcw     �<�V뒣�w��  X}���)e��Dŉ    IDAT�`TU����v`��{�a8�]    �2IC(%y�3v  ��܁�Ҹ��s�,�(v���\Nj�_^����z?�Aw��k��     &��]�  ��g�L��јKC���EeÆj23���(aii�{��<v     �/4׆={�}  ��_�����n�QU���Z�����0t�    `"��k��w��   V��;01��\9i4����(=�r�E�� �i�ӟ�bw     �rJ����  ��2p&ƫy~W�﯍���z啵�TJcw ,�n�ȿ��N�     VX�}S�  `u��#Ϸ�N�QU���Z����[yh�C�     VX�����܅�3  ��c�L��jys~���K�S���\���:���ǽ�     ���j�},v  �z܁�pdv��$���FQ媫\o&GQ��׾�I���     �"d��  ��c�L��߿/M�4v��4M�7Vcg ,�����p��0v     �'4�W��9�X  S���i�s{�E���+�ڵ��&Bh6��}���;     Xe���W����  ��0x�^س��6��bw�(�n��z;01�g�ɓ� ��      �N�b'   ���{�|��J��bw��I��|饵� �ax�`��cw     G����  X��ثv���n�QTٰ����i��SV!���;�3     �'�Z���}^�  `��c/Ͳc7�(�^qE5v�r����-��     DB��v  �<w`�5v�>'ɲ��;`��ji��܁�W�ZE�{����      �R�sg�  `��c-�v�!�cw���n�XM��4v���>�L'��C�     �Yvm�  `��cm���� ��v���co��+��?�s?v     �!���Gfg���  �,w`��ͦ7��7���^*]xa%v�))��?�L'v     �%��gc7   +��[Gw�6�vϊ���z��$M�� �����b~���    �h	Yvk�  `e�c+����0��7Vc7 ����E���cw     0zB��ᅻ�^�  X9����tn�� ��t晥�y�cw ��������;     =iQT�]��A�  `��c)<�`54����QS��j�$i���U;6��R/v     �+�v?�  X9��Xz�С����FM���k� NE��g;IQ��     `�����  ��1p�Ұ����0jJg�Y*�{n9v���������     ����~��ݻϋ�  �w`<����N�QS��j���V!��7��     ��J���;  X���	<�6�Z��QSݸ���d�^x�[,-�;     �۽#v  �2܁�s�ر{�ʱ;`���>�T:�?�x�v�޾}��     ���j]�  X��ةt�w�n�QSq�c�}��!�C�     �G��{h۶��;  ��g����e�c7���n�X�� p2B�9�����     ��R�b7   ���+Gw�>/�t.�����n]��n]9v���>�\���     ��<�@�  `���%�w&!��3`�T6n��n 8�k�����cw     0��ͫb'   ���+�n���`�T/����d��>�'!��     `\�z�ؾ���  ��2p�J9˼���t�٥Һu�� 'j�����bw     0�j����  ��2p�Ƒm�.N�|]�%�ہqBȿ��<v      �o��   ,/w`l�!̆��0J��^j����O~�ǎcw     0�B�yyس��  &�|`l�y~K�%�g�J�_��pB�"���N7v     b08����  ,w`lYvU�%��.�&I�[���{�^h4��     L�r����  ��1p���]�<_�FI��K+� ND�vCo߾<v     &�o��   ,w`,4�|{�%��LZ��Bw`��~��n���    �����Þ=60  0!<�c�����FIeÆj��i����������     L�������?v  �<܁�eW�N�QRٰ���Dt���&����     ��r����  ��0pF��]�<_�FF��V.��;�x�V1����v     VN��;  X���k����0J��^ZI��4v�����ycg   ���ޝ5�u�w^�n���Z�,K�d y����WQU��>� �9�;�ӥ����Y6�<)��{�5=�I������꽮���~Z�� Xb�ѣϥ�7�`  `	���r>�Vt���gW� �V��qW��Ut     K�i�����  읁;0|�۟�N��(�l��3����U�����     ,D1����  `�܁A{��߿��f'�;`(&�/O��U�7p t�u��/��    �B����  ����6�N��Rʣ;`(���W� �V����    ��<y�\t  �w����U�������'� O#}�a[ߺ�z;     �W��{7n|1�  �w`؞<�RtEq�D�?^Fw <��/̳���     `d�����  `o܁�z��m�����ɳϮD7 <���a[����     ,\1��et  �7��`�m�|���S��&ׯ����?v�    �����  ��1��N�.��"?|8//\(�; >M��q�ܺ�z;     !���ԝ��K�  ������ӯF7�PL�_�dy�Gw |��'?�����     `�RJ��ɓ�;  ��3p)�������������+� �&mow�/~�z;     ����o�  ��3p��W_��Զ�����&W��� ^��s��    �����  `�܁A����`(&�.M��Uo60hi:�^r�    �x��>��:�  쎱0H�|����������OS����iRt     �)�����;  ��1p)=yr-��br��$��OI�y�]o    `@�l���  ����������Y]�Ew��Eq�D��Կ��<�箷    0i>�rt  �;���4��?D7�P�\��z;0l]������v     %��t�]  @~���Ͽ� CQ>��Jt���ܺU�Ǐ��     ���9�����  `�܁�)��?� �PYy���p���/�8��     ��s���1�  �9w`P|�{�i:=�CP^�8�WW���OҾ�Z�=x�z;     ���f߈n   v���Y]�s���M�e���5�ہA���'��    0Xɷ� ��dD
J���&���|晕��Oҽ�V�޻�Fw     �'�NO߻q�7� �c�J�Ͽ� C��������i`��/��z;     ��gY^����  ��0���"��jt��ڵ�,������}�A�ܾ�Dw     �����_G7   ;c�Ɲ_�f�4G�;`&�<3�n �$�O:�R��     �O��S�"  ��;0������<��+W܁AJ�Y�ܺUEw     ��ȟ<��n޴� ��/��`t��ף`&�ϗ����h`���^�R�Fg     ��i��;/����  �����oo6����v`��.�/�4��     ��(�ڷ� �b��ϟ~��N�Fw��W��D7 |��W���I��     ��(��?�n   ���;0&��O)��-/ˬ<ޟ`���?����     ���f��  ��g�B]�� CP^�<��2�� �C�;Mz��6�     v���>���_��   ���;0E]9����zu� �q��t�      ��R*/=��;  ��c�B���Lt���w`p�Çm��Mt     �V5��Vq  8 ܁p�n�8�f��-?|8/N�.�; �P��KU�Rt     �Z;�}5�  x:�@�j>��<����6�zu��?���m���*:     ���N�G7   O��7����n�!�\�:�n �C�+�Ti6s�    �-��N޻q�lt  ��܁pyU}!����r����g?s�    �/��M��  ��3p�mo_�N�h��cE~�X�𿵿�mӾ�^�     �����*�  �t�@�����gRU�Gw@��ի���S�����     �7U���  ������ot���w`P��v׼�j�     �f:���  p �����ztAq�;0(��[Uj��     �7i6;����9�  ��܁X����c��͢X_�&C���^��#     `�u���G7   �1k:��3z��ˮ��Ҿ�f�>�;     `��M�[� `�܁0�����YU�Gw@���;00��    ��|�8  ��;&ϲ��n�!(.^4p#=y�5��^Gw     @/��g�  �?�����߈n�h��cE���=���/���3     �EU}k�|t  ���0��~�lr����p���_����     ������өo �3p�t��W� Zy���;0���Mz���v     �Z7��Et  ��܁o}����Z��h�K������z;     cPV�o �3pB����n�h��F�ol���f��}��:�     ��M��D7   ����V�ף ��ʕIt���oݪS�Fg     @��lv������  ���!��~.��M.]r���嗫�     X�<��v{�o�;  ��g���g�����x�w`��������o    `4յo ��2p�߿��c�l�����������Pߺ�z;     �R���  ��gX,��VW����Gw@��ҥI�e� ��6կ�RGg     �"u�ٵ�  ���7�N�"���/�� Y�eͫ��i>O�     �Hi:=���|f  d�,\�4��n�h�ŋ���,˲�嗫�     X���V��f_��   ���;�pi:�� ����3g\� ¥��s���     �y��ut  ��܁�J7oi:=���s�&YY�� ��~Ue]�     !���+�  �3p���ϯ�m{(�"�/��B���ut     D���g�  �?f�,T���o�^y��$��{���}�6�     ����rt  ��܁���W�1z�.���[���     ��W�����K�  �G��5���7F���,�#G��@�T���ut     D�L��   |���P�|~1�"��.M� �;w���Q�     ����	  �G����_��|~"�"M.\(� �W^q�     �,����E7   e�,̛|+K)��H���.���.տ���;     dY���W�  ��2pf��� �&��8y���j�x�Ϊ*Ew     � L���͛>� ��:�8��� Ry�|��o1 Bտ����     �?�v�������  ����SUע Ry�|� �[��T��Z�     CR��_F7   �g�,L>�]�n�Hw X���u�4)�     �$��_�n   ~��X�{7n���z=�"�g�N��q���:�     �&o��D7   �g�,F]�uJ)�΀(�ѣy�������]{���;     ��4�^�n   ~��X��i�� ����]oB5��V����     ��)��3ik���   ~��X�|>�ltD*Ν�b@��׿v�     >Fj�ɻu���  �w܁Ũ���	irႁ;&�穽s���     �������  ����f�s�&ϳ��w L���uj��     �n>�Bt  �;�@��ݸq6����R?^d�{s�0�o~SG7     ���Ms-�  �c;�w�i|��V^��z;&5Mjn�n�;     `��|~)�  �w�u����T�=;�n ƫ}�:k��     �6��N7o��  � ���]^ן�n�H�ٳ.�a�����n     �������/��m   w�w]U=� a�<+O���1�.կ��Dg     �Ap�,�<�  0p �f� Jq�X���zo����MVU)�     �����   �=����#yU��(���et0^ͫ���     pP�U���  ����3��7����a��3g܁(�y�w     xJ�|~9�  0pzV��E7@���Yw D{�^��<I�     p`�fg�   w�g��>� ��ӧ܁�믻�     ;Q�k�om���  ��3pzU������ol��#�Z D��Mt     4���7�  `��^u�����R�=�z;"=|ئ��o�;     �Y�/F7  ������OD'@���R�����     �u}=:  �������|�3YۮFw@܁(�k���     p U���  ;w�7�����T�>m�,�|�5o��;     �BQU�  `�܁ެ4�� J~�p^��{g��k��i����     ����N��7}�  ��B�&U�g� Jy���@��7\o    �]ʻn�ß��zt  ���;П��� Q�ӧ܁��}��     �`����   cf�����E'@�����X`�w�m���]t     dE�>�   cf|�"mm��|~"���N��,\�曮�    �^����  3w��7�s��&�"ϳ��Iw`��^3p    �=Ju})�  ����E�4_�n�(���E���Gw #3�w�{�     �G�|~>�  ����E[U_�n�(��Ӯ��ܹ�d]�     ^1��H[[>� � �@/��y&���N��.`�7�p�     �AJ�|��>�  ce����k_��hMΜ�׼���;     쓕��bt  ��Џ�:� Qr܁�<hӣG]t     ,�<��F7  �X���f������eV?�}�y�-��    `uu}5�  �� �w�����y������e��yt0.����     ��ʺ��   ce��Y�})���O���Ȥ�Z�    `_�Uu6�  ����w�R�ltD)N���ݿߦ�<Ew     �2ɫ�dt  ����&Ms-��'O��,Ts���     ��������tt  ���;�ﺺ�� Q\p�y�Mw     ���G���   cd��4���n�yYf����V`aRӤ��]w     �A޶��n  �12��]WU���q��,�<ϣ3�����mR�Fg     �Rj����  #w`_����ײ�Z���S����B5o�m�     =Im{)�  ���W'VW��g�֌R~�D� �K��[Mt     ,����G7  ���jҶ��n�(���"�m���3p    ���Uu*�  ���_m{-:���,Rw�n��6:     �V^U��͛�5  �`~	�W�^�N�y����U`a�߶n    �����}�+�  06�x��Ju}>�"�E>����x�o��D7     ��+��G'  ����*����ar�7X��K�ݻ�     г�m?�   cc�쫼�ND7@����2���޽6�mt     ,�I�^�n  ��1p�M��:��z-�"����T`aZ��    `!����   cc���M�\���+�Ra�,P����     � y]��n  ��1��MWU�E7@�����`4Rs�n     �PU��  `l܁��ҵ����eV�����8tti6K�     0i>ߌn  ��1p�ͤi�D7@���2�sw`!�{���     ��]}�����  �11p�M[�� B���=���o��     ����s�  0&y���k��:�T�����.�    �"uݳ�	  0&y�����DtDp�p��    IDAT�X�٬�<�3     `Lڪ��   cb�쟪ڈN�����S`!����,��     ��m�G7  ��������=����2�����6�     Ʀk�s�  0&��������n�yYf��z��Cw�~�      cS����  w`_�������Yfyn�,Bj��s�     ����  0&������jtD(77���B���4���     ���֣  `L��}�������;�-����v     �ж�o�8�  ca��Զg� Ba�,H{;     �����n  ��0��E�4�ouF�8~�[
,��;     �Y��k�  0Fy�����	�w`!�.��c�     AR�\�n  ��0��G]�N������]��A�5M��     ��j��bt  ��Q�g�?\Mu}$�-_]����<�X~�;�4�     0fE۞�n  ��0p���o\ϳ�ȗ�)67���B4��E7     ����=�   ca���jY^�n�����Q`!�����     ���7�  `,�=���RtD�76���"���w�     P�4��  0�y����3pg�r܁H~�eu��;     `Ԫj-ݼ��A  X �x{׶g� B�;� ��    @��Ry����Ew  ��{V4ͩ��P;�zg�     �0��k�  0�y����=� r܁��y��     ���D'  ��{���ft,Z~�p�������s�     ��Ȳ�  0����u�� �V��{C�ޥ�KO���      ˊ�9�   c`��I�y���z-����p��]z�}��    ` ڶ=�   c`����^:��TFw����P�w�t�     ��Ms2�  ��8ؓIU]�n�kk�P�w�{��     C�4��	  0�y���Yv)�"�yt������    �@��9�   c`��IS�� B���������#     ��V�k�	  0�y��L��TtD��ּ�@��G�RVU)�     �om{$mm��  ���iwF���[���mt     𿤔��e��  zf��I׶'�`�����<:Xn�     0@���  Xv�����9� �V�����<�     ��Jy~1�  ���;�'e�nD7��ǎy?�ޥ>p�     �PӜ�n  �eg��Ig������O�w���     ӥt.�  ����'y]�n�E+�ͣ�喦�.��)�     �Ms2:  ���;�k�_�u%k����p.�=�<p�     �(%w  虁�kw�޽���5�S�����Uz�n      �X�4ǣ  `���֥t)�B=��zպ�     ����Xt  ,;=`׊�.D7@���܁^�>p�     ��mף  `���Vtݩ��;г��\p    �JM��   ��@ص���D7��M&y���;П�KݣG�     0Du}$:  ���;�kyJ���h�ښq;Ы���.���    `�R*����>�  ���ص�m�G7���kk�N�W��C�v     ��y~>�  ����{)mD'����.��j?���     ,�L�D7  �23pv-o[wF'?z���U���2p    ��S2p ����4k�	�pG�x;�^u�     0lm{::  ����{mk���kk.��j?���     ,����  Xf�����X8܁~�d�     ��u�  �##=`������ɏu��Mz�$eM��;     �O��t,�  ���;�+���u$��Jt,Z��j���{���v     ��m� �G���<��}!�"G���I~h�     ׶�Ft  ,3w`W�8� ��Y�;У��#w     ��mף  `����tݩ�X�|u5�����Mz���     ��#�  ��܁]9����X����v�W�Ç�     0pE��n  �ef��Jj���h��;г�ѣ�      �i�mW�  `���R��Ft,����M�W�w     ���  ze��N��N�E�]p�4�uY]��     ��n�o[[G�;  `Y����n=�-?|���M���q;     W��Tt  ,+w`W:wF�w�O�ѣ.�     x:+y~2�  ���;�+eJk��h��@��<1p    ����>�   ���ؕ�uG�`�\p��>~��     ��S����  XV���4��;㳺��z�\p    �#ϲc�  ����]��Ht,���@o����     p@�]�;  ���ؕ��V�`ъU���I���     ��Y��   ���ؕ�m-}�|e�w�7����     pP���;  ���ؕ�iE7��:d����R�N]p    ��H�ht  ,+w`��͛E��Jt,�d�gEa�����NY�o    ���5p ���;���h=K�ЗQ���<П'O��     �饮;�   ���ر���ft,Z~�Pt�ĺ�m��    � )��pt  ,+w`Ǌ��Xt,Z�;Ч��w     8@R׭F7  ��2pv�m����p����S�    � i[� �'����4�Ft,Z��j��&mo�    ��R:�   ���ر*ˎE7�¹��(�f�     p�t�jt  ,+w`��,[�n�Es��S���     ��Wt�Jt  ,+w`ǚ�ۈn�E�]pz��S�    � Im{(�  ���;�cyJ���p.�=��    �`i[� �'���)�n�E+&��`���mw     8HR*�֖+�  �w`�����L\pz��&eMc�     ���ٌn  �ed��X�����1pz�f3�v     8��f-:  ���;�c]��F7���++�	�����    � �ő�  XF���Y�;㳲�;Ћd�     R�u.� @܁�k[w�g21pza�     S[��  �w`�R2pgt����`Y�    ���V��  `�;�v��;��;Гn63p    ���2� ����Y�5��O&�	��JUe�     ��  �w`��3pg|VV\p�1��    �A�uG�  `�;�R2pg\�"ˊ���E2p    �)O�w  聁;�c�w�f21nzc�     S�e�  �w`��&��H��C�@���     ��m� ���������e� ,��6p    ��K�Ht  ,#w`Ǌ��}w�G���     �]H)�n  �ed��X2pgd�ȣ���U��     p ��$�  ���;�s)����L���#w     8��]�n  �ed�
�X�:?;��t��O]�    �4�s�� @���X�g#��et��RJ�m�+     �]hRr�  z`�
�XJ��ƥ�<Џ�4�	     �.)M�  `Y�;�n�,2wƦ,��`I�u�N      v��2w  聑*�3��+���,��e�4�     p@Y�D  聁;�#��;� 7����"5Mt     �[)��  =0pv�j���X��s	�#u]t     �K��� �{��4y~(�-/}� Џ�iRt     �K)�   z`���z׹����e� ,'�    ��*���  z`���R�zҶ.�    ��R�D7  �2��v��:Ag|܁����N      v)��;  ��bؑ"����ɣ�����        a��HӶ~n0:)�m܁^��     W�V  ��Pؑ�����oz��.:     ح�|�  =0pv���2����I޶)�     �5$ @܁����F'7p����    �J�  �CU`g|�cTx.�~t�     p`�>? �^X�;���       ૠ ����������3>�]
��     p`%� ����<�N'��p�@_�.�      �=$ @܁9<�og�����    ��r�  za��H�eet,��@_��;     Tɡ,  腁;�#����\=�o    ����  z`��Ȥ,�       R��9  ���          �A0p          `�          w           ��          �A0p          `�          w           ��    �����-�m�gF��!�iYm����+JUbo�8%R%��  [�rve�>(vs�y��=�J��     � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           � p          �w           ���=       �r�<��45�w�i�z\�0��   �M�      ; �0��n�ǻ����5�����Ƚ   ([�{       p=~l�7�u�ɽ    >��      vDa>N�aȽ    >��      vHa:I�4V՘{    |*�;      옶��')����so   �O!p     �tc�,�W�w    ���     ��z�Փ�y�{    |,�;      찣�y�0�U�    �1�      �㞵��a]or�    �E�      ;.�0�t�B�so   �?#p     �=C���˳XUc�-    �G�      �'��')����so   ��     �9���ҫ�;    �C�      �g�x��i�s�    �$p     �=��i.�Y,V�w    ��	�     `O=k�7w�z�{    ���      ���^���;    ���      ��b��ry�j̽    �      ��Ɠ�NCU͹�    ���      @uc�SJg�w    ���      @UUUu?��QӜ��   ���      ��I�\|�X�r�    `?	�     ���Y۾�[���;    �?w      ��<O�lY�}�    ��;      �O���=�U5��   ���      ����"��uUM��    ��      �Z�8��ҫ�;    �w      �Oݏq�]Ӽɽ   ��'p      ���M�z�X\��   �n�      凶=��U�    �.�;      �Ѧ�(�    IDAT���e]�    �&�;      ��B��ry���1�    v��      �$M�IJ/몚ro   `��     �O��q�1�W�w    �[�      �g�����y�{    �C�      |�GM���bq�{    �A�      |����^�W�w    p�	�     �/��m_-�˽   ��M�      |���"��&�m�-    �^��  �?7�s8�n��so  `���&�1�n��tܶ���u�M�m   ��  P��86�5�7����  �~9j�sq;�c��<���v�ӹ�B�=    �.�&  @�Ά���w���v   nړ�y��i.r��������y�{    ���  P�a��}��j����   ���qu�4�r���{�4�y^��n��   ��!p �����ߺ���kK   d� ���Rru�k�}۾�����8�ɽ   ��A�  ������  �\��x�SJ�s�`�<k��]�-6Ӕro   �|�B @f��q�o���v   r9����}�{��a~��i{    �� @&�<������t��XU1�   ��2��$��:�9�vWa:n۳����[    (��  2�NS��������[   �_mË�R�΍H1�S:U��    H�  7�rқ���0ϋ�[   �_M�������ܘ�1n�o�7�w    P.A  ܐi���fs�O��p   ��U5�H�e{��QӼ��y�e;    >DX  7`��6��?��9��  �~��j:I鴭�m�-�����v����N�-    �E�  _�TUa��t����   ��擔Nb�so�gm�z�x5M��[    (G�{   �~�����  (A������c�ro����:��8��6�!�    �!p �k6WU��������<�!�   ���z�ҫ�1�s�ߋ!L')��U5��   @�  p���T���w�Ðro  ����i^?��*�������)����    `�	� ��\Cz�^��NS̽   ��iӜ?j���w���c�,�W�w    ���  ��4��|��s����[   ��/�6�E��1�x�x�x�{    y-r  ��l��6��?��9��   ���b���m����⻶};�s|7�wso    �;  |����j�9�Ʊɽ   �у/����;�s�ضo��[\M���    �P�{   �6�8.^_]��  P�;u���m_���+�0�tֆ0��   ��� �G���Z����fsg��{   ��e]w�)����[�K����NcU���    p��  ���T���w�Ðro  �I!�/R:���숶���)����    `O� �_���f������{   |H��b�<�!L���u:��{�ҫ�;    �9w  ��<�����e�/so  �?�j<I�t{|c�z�4os�    �f,r  �m��f���<��[   ���U5�%��m]oso���i��ߎ��[    ���  �;SU��fsЍc�{   ��PUӋ�^���[�&<k��뚫i��   ��s  �Rt�x}uuO�  @�BU��)�����7%�0�tֆ��:    v�� ��7WU�������<�!�   �3���R:��&��i1��d�<�U5��   ��!p `�m��>_�ﮇ!��   ㇦y}?�u��K��$���    ��;  {�rқ���v�b�-   �1�������̽r;���1�W�w    p��  �i���z}��   ��z�4o�4�E�P�1^=i���w    p��  ��vۼ^��ӴȽ   >�7���i����9j�w�u�ɽ   ��#� `/LUV��A7�M�-   �)���Y۾ɽJt>w���+}    ;D� ����qq�u��<��[   �S܋�꧔^��%�ǃ��ǹw    p��  쬹���}�\Cʽ   >�a]o����;�D��q�k�=ɽ   ��'p `'m������4��[   �S-�;I�4�0�������]�d�*��   � �;  ;�r�e�/s�   �ϑB�_�tZ���lƱ���NUU��   ��!p `g��T��&߹   �JMۓ��4�0����i�s���   v�� ����n�U����ij   n�XU㋔^6!���@i�i�?w��XU1�    �.�;  ��TUa��t����   �����EJ/ۺ�������뎆y��&   ��@  �Z�8..����v   n�PU�qJ����[�4�<�?o6G�<;n    �'�  �:sUU��~���{   |�PU�O)�݉�˽J3�s���l�ͽ   ��#p �V�NS}�u��i���   ���1�W�c\����{ܾ��e�-    �,�;  ���0�˾��&   ;ᇦy� ƫ�;�D������t�{    7O� @��i�W]w�O��W   v�QӜ?j���w@����]���;    �C  @�6�m����y�C�-   p/�4�E�P�����o��^�    �#p �HSU��fsЍc�{   \�ob\}׶os�������w    ��� ��t㸸�CW�  �%b�|�қ�;�Do����0<̽   ���  c���}�/�Ðro  ��t���?��*�(��q<�m�ͽ   �2� (�0�q���i���   �u:�����r���q��]�8�    �!p  ��aH�}�̽   �۲�������[�4������Uro   �w  ���^u�A?M�K  �9m�IJg1�)�(�zۿ��   � !  Yl��f���<�  ���j|���Ec�-P�~��t�ө���[    (�� �5UUXm6�86��   ��PW����^6u-n�0LS���滱�b�-    �I� ����qq�u���  ��ꪚ^��2�8�����s��뎶�v    ��� ��n���}�/�Ðro  ��%T�|���A�}�-P�q��_��i?�^�   �O	� ���q���?�N��\   �PU�O)�݉�˽J3�s���n��ͽ   ��	� �j.�!]��2�   �ڞ���~���;�4�<��vݓ�4y�   ��"p �ڍ�T_t��0M�7  �y�5͛�1^��%���_N�A�    ��#  ��f�mV}0�sȽ   ���Ms��iV�w@�~�oW�x�{    ��� �k1UUXm6�86��   �M�v�x��i.r����߼ǻ�w    p�� �b�8�/{�����m�$�����HJ��������'�h�$�*��?�d�I�;�$�I�s�!�-pq:�^m  স�-��Kw@��{��l��    �j2p �O�M�|���4��-   ��	���ߔ��Lӝ7�ͽ�    \]�  �)SJ�|�6�J�   �ײ�u��˓�P�w�t�izX�   ���� �?�b���8�Jw   �״��y�Gm���-P�Ӕ���ǥ;    ��� �di���aؚ��w$   7Jl�q?ƣθ~�CJ����   ���0	 �O��l��q��9��[   �kZ��Z���K�@m>�_�nngF    |�  ���iڳ�zkL�/�   _[h��|�:Z�m*���Li�¸   ���� �kLiq:�^m  �&�fޏ�pٶ��-P�q�/�awn��t    ׋�;  �����0���i��[   ����q�*��t�f�9�^j�P�   ���� �_�R
�㸵�g�   �Hm��g1o�0�n�ڤ����zo��=#    _��'  ���4ŋq\��   ����xr;�u���/��1�t    ח�;  M���l��y�}  ���m߿����P�9��`v�9/K�    p�0 �p�ͦ?ǭ�s[�   J���w��C��͜s�rv��K�    p�� �PsӴg��֘�_J  p�������?+�5z5��/�y�t    7��; �4��8�m��  @�<X,�����t���0<:Oi�t    7��; �s>���i�;i   h��^O�˷�;�F����iJ�Kw    p�� �SJ�|�6�J�   @nw���OJw@�~��o7���;    �y� n��i��*�   ����w1���Lӝ���^�    n&w �k,�ܝ��[�<��  ����vx�q׶�t���fs�izX�   ����	 ��Zo6��8n���-   P�e�N���Qh۹t��4����q�    n6w �kfn��l��S�K�   @MM��W�C�v���V?�q;    �� \#CJ��a��j;   �Zh���a߶�t��"���0��q�   @q�  ���8n��iY�   j�5��<ƣ�T�js���q;    1p �⦔��0l����-   P��i���BK�@m�y^��ݹi�+   Pw �+�b���8�Jw   @�ڦ�Oc<��P�j3�s8���4�t    �_�  WPʹ;[���y�=   �Ɠ�?��e��Mʹ;��)ggK    Tǡ ���l��q��9��[   �V��7���c���/��1�t    �+�  W��4��z�5���   ~�^߿{��Jw@m��ð���e�    �w� ��!���0l{�   ~����t���Jw@mr���aع��X�    ~��; @���qk=M^�  ���~��,��Kw@�����U�    �w �JM)��a�N9w�[   �v�B��{�oKw@�^���Kw    ��0p ���4ŋq\��   ��`���O��7�;�F�����fs�t    |*w �������z{��P�   ��U��c<��6�n��Nӽ�����    �G� Tb����㸕snK�   �U��q߸���i�s<M�Kw    �e� P��4��z�5�ԗn  ��bٶ���B�Υ[�6�6�[?M���    �g� 4��8�m��  ��M���VG��M�[�6�)m�8��Kw    ��e� P��8n��iY�   ���i���m�)��9Oi��0�   p�� |eSJ�l�S�]�   �Jڟ����-P��)��a77�?   p�� |E�/�qU�   ���i���BK�@m.SZ�0n   ��0p �
R���z�=�s(�   WM�4�i�ǷCX�n�ڌ�x1�s��[     ׂ�; ���l��a�.�   W������.Kw@m����0쥦�    ׆�; �27M{�^o�)��[   ����w��C��Mʹ;X������   p�8� ���gð�snK�   �U����w���t�&���ޘ��    �v� >��q�ZOӲt   \eB8�����P��s�rv����	   �k�� �3�R
gð�r�J�   �Uv/�Ob|[�j�sn_���y^�n   �/�� �3���x1�.  �/��ǧ1�)�5z5��.�y�t    |I�  Aʹ;[���y�[   ����w��I������,�[�;    �K3p ��֛M6ۥ;   �:Xu��<ƣ�ms����q|�>�;�;    �k0p ���i���1��t   \˶��c<���7������n�    �Z� ��!���0l���-   p�m��_�C�Υ[�6'�t�x���    ���� �����z���;   �M��c<��6�n�ڼ��[?M���    �� �SJ�l�S�]�   �.�����x��M���YJ[?N���    P��; �︘�x1���   p��M���x��X�j�!�իa�)�    �� �i���a���s(�   �I�4�i���!�[�6S���Nn��t    �b� �O֛M6ۥ;   �:z���.Kw@m�)�/�awn��t    �d� �iڳ�zkL�/�   �ѷ}��~Kw@m�y^Þq;    � 4M�4CJ��a��9��3   |�}��a�(����9�^j�P�    j`� �x�ͦ?���   p]=^,Nw���t�&���ޔ�;;    ��� 7^��7   |!��o����;�6?��wǜ��-    Pc.     ����œ��m��Mι}1;�y��[    �6�     �gw��.��\�)���e�~9ϫ�-    P#w     �Zu��,��ms��ͫq|t1�[�;    �V�     �g�v܏�3n��x=��R�U�    jf�     |˶��W��жs�����������    P;w     �/M���x�h�T�js<Mw�l6�Jw    �U`�     �%]�����p�u��-P���t�p���    ����     ��ڦ��c<�!L�[�6�)m���G�;    �*1p     ���i���BK�@m�SZ�0�Kw    �Uc�     �am��1�a]�js�R�~vsӴ�[    �1p     ��o����.Kw@m.SZ�4n   �?��     �C�������t�f��ŋa؝��   ���p     �d;}��qߟ���L9��Z��IMJ�    �Uf�     |�����^ߟ���lr���Ƹ    �2w     �?�o��w�;�6)���0�9��[    �:0p     ~ם>>��M��͜s{0��y^�n   ����     ����n��ryR�j3�ܾ���<��-    p��     �Ҫ��1�m�K�@m^���y�*�    ׍�;     ��m���:�v��W���<���    p�     �ҷ���ju�v.��y=�NS�]�    �+w     ���I�1�m�J�@m~��o7���;    �:3p     ��i��i���]�)��9��;'�ͽ�    p��     M�4�Y�G���-P�w�t�izX�    nw     ��ڦ���xt+��t��t����ǥ;    �0p    ���1��	a]�j�!����    �U�    ��m߿����P��)ŗð���-�    7��;     �P{}��a�(���Li�¸    �0p    �h������Y���8ϋð;�G   �"�    �� ��?-���rð��&�n   ����     n�{!\<��m��Mʹ;X�����[    �&3p    ��v�]>��t��q��s_�    n:w     ���n�]�ǥ;�6s���0�s^�n    �    ��[u��,��ms��ɜs�rv��K�     ���     ��e�N�c<m;�n�ڼ���U�    ���    ��
M��c<\�m*��y5��S�.�    ���;     \C�i�?b<�θ���q|p����    �o�    �5�5��<ƣ�T�j��8����-�    �k�     p��M���x��X�js2MwN6�{�;    ���     ���i���o�0�n�ڼ�ln�4MKw     ���     ��'1���t��4����q�    �?3p    �k���{?���;�6�)�~�v    �"�    �����w����t��"���0��iK�     ���     ��ǋ��nߟ���\��|i�    W��;     \Q�B���r��t�f��ŋa؝݅   ���P     ��;!||��P�i���0쥦	�[    �?��     ���[�\���ڤ���a؛r^�n    �w     �BV]7<��m�\�j�˸}̹/�    �y�     pE��n܏�3n�_�9�/�ag=���-    �_c�     W��m��1���K�@M~�_��t    ���    @�BӤ��ѢmS�������b��Jw  �/K    IDAT   ���;     T�k�y?��e�nJ�@m^���Kw     ���;     T��yܾ
a*��y=�N7�ۥ;    ����     *�6M~��Vc����4�{���-�    |~�     P���xr;�u����4�9����;    �/��     *�m߿����P�w�ͭ���a�    ��1p    �������}��t��,����q�    ��2p    �J������?+��9Oi�jvJw     _��;     T��bq�����;�6S���nn��t    ���    @a�B�x�\�-���Li�¸    nw     (�v��xR�j3����0���    �Fq      �lw����Ҹ�ɔs8���4�t    �u�    @����xܵm.�5I9w��ޔ�t    ���    �W�l�i�:
m;�n���2ns�K�     e�    �WԷ�f?�C�v���s�rv�9/K�     ��    �W�&��x�w]*�5�9�/�a��<�J�     e�    �W�5��<ƣe�mJ�@m^�㣋y�*�    �g�     _X�4�Y�G[!��[�6?�ó�n��     �`�     _P�4�i�ǷBJ�@m^���)�)�    ���     ��'1���t��p���l��     �b�     _ȷ}��~Kw@mN����4�/�    ���     �������?��ڼ��[?M���    @��    �3{�X����Y���YJ[���Q�    �^�     ����o����P�)�^�Nn��t    P/w     �L�p��ߖ��|L)~o�    |w     ���n�d�|S�j�N�1��{)    �8H    ��h�u�����ͥ[�&c΋�a�3n    >բt      \e������7�yð��&�n    ��e     ���l��y�G�m��-P��sw0{S�[    �w     �BӤ�1-�6�n���<n�s�K�     W��;     �A]���1.�nS�j2�ܾ���<��-    ��d�     @��}�T�j�j��U�    ��2p    �O�6M~��Vc��ͫaxt��v�    �j3p    �O�6M~���֥[�6����iJ�Kw     W��;     |�o��7wC�,����q��v��[�    ��    �?���w���P��i��f��W�    �>�    �w������?+��y;M���A�    �z1p    ���bq�����;�6�)m���G�;    ����     ��{!|x�\�-��9Oi��0<.�    \O�     �O���i�oJw@m.R���nn��t    p=�    ����u��˓�P�˔�/��   �/��     ~���y�Gm���-P�q�/�awv�    |a!    �i�e�N�1u���+S����oRӄ�-    ��g�    ��׷�f�:m;�n��lr���Ƹ    �J�    ��BӤ���M�[�&)���0�9��[    ����    ��k��y�Gˮ۔n���9�ð���e�    �f1p    �Fj�&?��h+��t�dι}9;�y��[    ����    ��m��4�����-P�W���b��Jw     7��;     7ΓO�pY�j�j���]�    ���    �Q���7�C�X�j�z��t�t    p��    pc�����}��t��������n�     w     n�ǋ��Nߟ��ڜLӝ7�ͽ�     Mc�    ��`�8�f�|_�j�n�n�4MKw     ���    �k�^O�˷�;�6�Ӵ��4=.�    ��    pm��˧1���ڜ�����    ���;     ��V׭��x\�j�1���0��iK�     �3w     ��ض�����ͥ[�&�)-_�    3p    �ZY��Z���K�@M�y^�����    P1�     \�i���m�J�@M�yð��&�n    �=�     \]�����p�u��-P��sw0{S΋�-     ���;     W^�4�~��1��t��q��s_�    �S�    p��M���x��X�j2�ܾ���</K�     |*w     ���i���o�0�n���9�/�a�r�c�    �?��    �+�۾s7���P�W���b��Jw     �Q�     \I����}Q�j�j���]�    ��0p    ����������t���8>8M�v�    �?��    �+��bq�����;�6?��������     ��;     Wƽ>|�\�+��9��;'�ͽ�     ��;     W>>��M��ͻi���4=,�    �9�    P��[�\���ڜ����4=.�    ��    P�U��c<j�6�n��|Hi��0�    ׊�;     Պm;��x��ï\�_�nn��t    ��d�    @�����VG�m��-P�˔���    �ue�    @uBӤ�m�J�@M�y^����    pM9�    �*]���1.�nS�j2�s8���4�t    ��b�    @5~��B�J�@MR���0�M9/J�     |I�     T�m��4����-P�_��c�}�    �/��    �*<���N��P��s�bv��,�    �5�    Pܷ}��~Kw@M~�_��t    ��b�    @Q{}��a�(���~_��V�    ����    �bv���Nߟ��ڼ�G�)m��     ���    (�A�{}Z�j�z�n6�Kw     �`�    �Ww/��'1�-��9��{o7���;     J1p    ૺ�u�Oc<)��9��;��t�t    @I�     |5�]��.���P�w�ͭ���a�    ���    �*V]7<��k�\�jr��֏���t    @�    ��m;=��8��\�jr����0��     ���;     _Th����mS���ǔ��ð���-�    Pw     ���4�1�]g���:���q;    �o�    �EtM3?��(�0�n����8���=    �o88    �k�&?��h+��t�d�9�^j�P�    �F�     |Vm��1�
a(�5I9w��ޔ�t    @��    ����xr7���P�_��c�}�    ���    ��������c��Iι}9;뜗�[     jg�    �g��������P��s�bv>��t    �U`�    �_�h�8�����P�W���b��Jw     \�     �%�C8��r��t��axx�ҭ�     W��;     ڝ>�=Ʒ�;�6��������     �j�    �S��n��ryR�js8M��n6wKw     \E�     �a����xԶm.�59��;��t�t    �Ue�    ���q?ƣθ~��4��i���     ���    �d˶���x�v.�59Ki��4=*�    p��    �IBӤ��ѢmS��ɇ�V��a'7M[�    �3p    �?�fޏ�pٶ��-P�˔���    |6�     ����q�*��t�d�R0{��    ��Ɓ+     �V�4�Y��[!��[�&c��v    ��oQ:     �z�=Ɠ�!�Kw@M�yð��&�n    �n�*    ���m߿����P��s�rw��="    ��    �{}��a�(�5�sn�aw=���-     ו�;     �����w���t�dι}�?��X�    �:3p    �=�|��OKw@m^����*�    p��    �4M����I�oKw@m^ã�Kw     ��     4�C��4Ɠ�P�����4�ۥ;     n
w    �n����-����O~��o7���;     nw    �lն�����ͥ[�&��t�d��W�    �1p    ���m;�V���O�N���izP�    �&2p    �������x�v.�59Mi��4=*�    pS�    �0�i�~��}ץ�-P�)�~�ǥ;     n2w    ��k��y�Gˮ۔n��\�_�nn��t    �Mf�    pC�M���x��X�jr��Ҹ    ��     7@�4�i�ǷBJ�@M�y^���ٝ	    @�    � Ob<��e��ɔs8���4�t     ���    ��������c���&�p�^�M9/J�     ���    \c�}��a�(�5I9w/���1�t     �f�    pM=^,Nw���t�dι=��u���-     ���;    �5t?��o����;�&s���a�Y�s,�    ��f� �?v�"���[U3Y�$��h� ���3m@ԍ��Ƭ֡��g�VT�f�繱�4�?�Û�?_   .�k��\,�=z���������F�     ��    \ �9�����y�����էG�^�    ��'p    � �伺�X��Rꣷ��|�Z}�փ�;     �cw    �`����b�c���w���ߵ~4z     oG�    p���{�ʏ%�6z�����������     �=�;    �9V"����)�:z�ɓ�f��fs}�     ��;    �9�#ڿ�vsގ�s�t����f���     �yw    �s(E�����R6�����z�[q;    ��%p    8gRD��X��W�z����Z߬V7zD�    ��F�    p���~k��頔��[`NNkݽ/n    8��     ��W;;?T���0'�֦��Ս�    ���    ���bg��';;ǣw��lZ+�V�/jD�    ��O�    p|�������2z�I�=�[����>��    ��!p    ��O��苝���w�����׽��    ��#p    ��k�,������;`NZ���ju㬵��[     x��     3uX�ɭ����;`NZ���j��ik��[     x��     3t5糯ww��s�p��층��;     x?�     3s%�՝��ǔR����j��Q�WG�     ���    ��"������,n�7|�^�փ�;     x��     3����Ε+?����-0'������~4z     ��    `JD��X���R����fs�x��6z     ��    `���.?������f��h��>z     ��    `��o/?^)e3z���Z�~��|6z     ��    `��o-?헲��dY�oW+q;    �%$p    ��b���RNG�99�u�`���#��-     |xw    ������Z)'�w���ֺ{_�    p�	�    >�/vv�\��Y��s�nm��Z�h�]     \j�    >�Ϧ���;;���s�i��[���e�     ��    | �L�ї���7z�I�=�[����>��    �xw    ��Z)�������0'/��u�;��     0w    ��l?��[����;`Nz���j��Yk���     0w    ��h/�ۋ�O�w�����O[�2z     �"p    xO�伾�X��Sꣷ��|�^v����     ̏�    �=�Misg�����Fo�9y�^zT���;     �'�;    �;V"����)�:z�����'O�ۃ�;     �/�;    �;�#ڿ�vsގ�s��fs����G�w     0ow    �w$G�����R6����<�l�l>�    ���    �)��^,~�+e=z�ɓ�v��fs}�     ·i�     ���띝��)պ��zO�ED��"Z��Go��Z��[�?�    ��C�    �7�,eyѣ��_W���_�
�s��SD��z�����ܞ�}Q<��Q�W�V���    ��"p    ��Q���9o������Dk�A������׃�H�G�=��zD{�c]Ϝ�Ժx�Z}����     ��'p    ��n�|�iΫ���WyĿ�����u��{�=�_��g!���]:�u��ju�E��[     8�     ��9��(�l�׼q��s�u>���������󿾈�?�l.�ukӽ��q;     ��    �O�$�՗�����W��
�{yv��e����^xv������z��^�/����˽��QFo    ���    �	��������?zޥ�H�ڛ��_�/B��_^}���Z�D�B�=�;;�bӻ�     �-�    ��~J�[�t|	����"�Dk�zŞ�G������%�)��,~o��grμ��׽��    ��'p    x{)mo�����=�����o�^�g���>�������Ӄ����wGo    �b�    ��ED�3M�<z���?��Z����<x=�O9���Y ߃az���j��IkWFo    ���    ��݈vwg�<����RD����<~�GN���zzv齥�[�xq��?����z��qk{�w     p��    ��)��)�h��NJ)zDN�G�^"����Տ��R�)���[DK)�Q�/�oW��Ժ?z     ��    �7��~���ݜ��-�%)�^����)�E�-E��{����w��������_���w     p1	�    ~%G�;�-�����9Z�/����s��{J-Rj=�ų�����a����v{m�     ..�;    ��|]�r/�:z\����_��=��������%�o6�?m6��    ��&p    xͭR�9oG�`^RD�֦�5���%|���?�l���    ��'p    x�R�������2��Ժ��f���     \w    �������9�G��b����)�9�x��H����f�/k��p���G��[     ��    ���yΧ�����-������ߏ�.��T{J/���;_8�u�q;     ��    �Ԯ������;��^�����}�)����{��"|���׭M�W�-"��O    ��#p    .�k)��*�d��/R���KDD�="RD��[���뻌�7���9;��F�w�g    ���    ��aJ���t<z���_J��2z���=�\SD���\SJ������˽�ꋭ�    �A�    �������iZ��C�I)Z�^�qO���)��R��kv���?����V7ֽ�|��     ��    ������뜏��\)z/�����{D��R�)��/���ӽ���Yk�#    ��    �4v#��iZ����?RJ/��xv�G�oj=�    0w    �R�"ڝR���^��p�=X�.n    `��     �[��wK9�͹��s�#����/�v     fD�    \h9��)�h!n�7��v���/F�     ��	�   �+G�ۥ,�r�����<�u�߽_�     ~M�    \X�JY�����qk�ǭ��    �%�;    p!�*ey(n�7����G�^�     ��;    p�����k9oF�9y�������     �G�    \(7r>�4���0'�֦����     D�    \��|v����;`NNZ+߈�    8'�    ���IJ�/K9��䴵r����Fo    ��!p    ν�RZ5M'�w���Z��k=�    p��   �sm?�ͭi:V��+���Z��      �3�   �sk/���R��vxe��o�[�  �[�    IDAT    8���     ��ED�3MK/�R#ҽ��pQFo    ��·    ��ٍhwwv�JD��Gă��`%n    �s�    8W��v���I�/���A�'�{�    �\s�    87JD�[��n�m���k�_��3z     �]w    �\��N)Gq;��#�����/���     ��    ��ѿ.e��s����v������     ��   �ٻY��A���;`N~���Ͻ_�     �%�;    0k_�r�QΛ�;`N�������;     �]�    ��e)'�s^��s��G�^�     ��;    0K7r>�,���0'O[������;     �}�    �s=�ՍR�F�9Y�6=��`�     x��    ��\Ki��i:��䤵�    �K@�    ��AJ���t�F�9m�ܯ��E�W    �O�    ��~J��ӴT��+����Z��     \w    `�����vxӦ�t����-    �Kģ8    0�nD����c%��}�o��    p�x    ��"ڿJ9�r�\Ԉt���uD�     >4�;    0D��w�����ۃ��    �Kj=     �|JD�S��"�6z�E�=�zpһ�{     .-�   �*G��KY��\Go������e�;��     �Hw    ������~���;`.zD|��^�����[     `4�;    ���*ey n�7<�u�I��;     `�    ��RN�����Z���ڕ�;     `.�    �{w#��Os^��s��O���     s"p    ޫ�s>�Q���0'OZ�}T���;     `n�    �{s=���vx�/��|W���     0Gw    ླྀ����RNF�9Y�6}+n    ��J�    �s)mnN���0''��oj=hi�     �+�;    �N������^9m�<��P�     �O�    �3��z;�eN^xa�Z�_�A�    ��    ��nD�[�єs��b���zX��    �[�    �mSD�#n�7l#ҽ��p�-     ޚGu    �o)�n)G�9��[`.jD����#��-     p��   ��,G�;�-���R�������     �4�;    ��~���^�u���q�I���-     p	�   ���f)��9oG�9�v��_��3z     �W.�     ��R����G����է���     ��    ���e)'����j�{��b�     8��    �[����g9�F�9���+?�ve�     ��    �[���ٍR�F�9y������F�     ��B�    ���SZ�����;`N�����֫�w     �E"p    ~�G)��9M'i������|W���     p��   ��j?�ͭi:��+��&q;     �w    �7��=MKq;�r�Z��փ�_     x�    �XD��9/= �+g������    ���}
    x���r4��Go��X����zP��     �^	�   �����/q;�a������M     �;��    @DD��~���ݜ��-0ۈto�9�zO    �<    9��.�h!n��jD����#��-     pY�   ��U��j�u����l��g�v     ���    p��*ey��v����ۃ��wFo    ��F�    ��W�_�y3z�ɷ���R�     CL�     c|�����ףw�\���֫O{��     .+�;    \B��|�y)g�w��<�n�����     .�<z     �a]Oi�����c�W~����     p�	�   ������i:�����?��7z      p   �K�0���i:���Ik��[���;     �g�    p	짴�z��i���ek�w���     �"p   ��JD�:�cq;�r�Z��փ�;     �7	�   �ۍhwJ9*9��[`.N[+j=l��     ��;    \P��}��K����Z��     fI�    P��wK9�͹��s�n-��    ��	�   ����N)Gq;���H�k=�z    �Y�F     ޝ�o���˹��s�m-ݫ�pQFo     ~�K5    p��*e���v���Z;X��    �\p�    .�[�,���R�=�zpڻ�p     8'\p   ����\�y3z�E�����/{��     x{w    8�n�|�iΫ�;`.zD|_��_z��     �s�    p�}��ٍR�F�9yT�ޓ��w      ��    ΩOr^}Y���0'�j����+�w      ��    Ρ�RZU�I=f�qk���v     8��    p�짴�5M��vx�Ik��j�:z     ���   ��Ki{����^y���w���     �}��    ��YD�;Ӵt�^Y�6=��`�     ���-    ΁݈vwg�D��[`.NZ+߈�    �B�   ��M�N)G��^:m�ܯ��E��[     �wG�    3V"��R�vsn���\�Z��k=�    ��#p   ����N)Gq;���=߫��z�    ��     ���o���˹��s��H��ۃ��m     ��|    ��g)��9oG���fs��(��      ��    f查_�y3z�E�����J�     �4z     �ʗ��|��z����{<���w��     p	��    3�yΧ����G��Z�����     |w    ���9��(�l����o�W�}w�     ���   �`�RZU���0'��۽'�/F�      >,�;    t����4��s�C�W~����     ��'p   �A�S�|=M�4z����?��7z     0��    �Ki�u���vx�Ik��j�:z     0�4z     \6���4-KD���ik;�պ?z     0��    �M��4-'q;��lmzX���     �xw    �@JD�[��nJm������7�v     �9�;    | 9��)�h����;m�ܯ��E��[     �y�   �{�#��R�{9��[`.V������    ��	�   �=�U�r?���0��ҽZ�7j     �W|<    ���V)�Cq;��}�o�O     ��    xO�Q�ɵ�7�w�\Ԉt���uD�     �'�;    �7r>�4���0="l�+q;     �;��    ��,�����s�{�����M     �].�   �;�IJ�/K9��G��Z�����     ̟�    ޑk)��9M'�w�\��~���Kﻣ�      ��    ށ��67��x���G��=�}1z     p~�   �o�Ki{��e=f�Z���ڕ�;     ��e=     γED�3MK�$��ǭ-~jmo�     ����    ��݈v����Go��x���Z���     �Ow    ���v���)gq;<�Kk;�պ?z     p~	�   �O*�n)G�9��[`.��Mߊ�    ��I�    B��wJ9Z��ᥓ��7���4z     p�	�   �-��u)˽���-0������    �wA�    o�f)�9oGX����zP��     �;"p   ���U)����b���zX�3     �    ��,��z���;`.���fs���     �c>>    �︑��g9�F���fs��(��      ��    ���)�n�r6z�E�������     xO�    ������4���s�"n?�}�     ���    �+���9M�i���o���e�;�w      �K;    ���6����R���۫O{��     ��\p   ���R�ޞ���^yT�ޓ��w      ���    "b7���y��^���+?�ve�     ���   �Ko�h�*�hʹ��s�ŏ���     \.w    .5q;��'��>����     ��#p   ��*�v)�ݜ��-0O[������;     ��I�   ���#�ץ,�r����\,[���     �Hw    .�[�,�sގ�sq�Z��փ�Fo     ./�;    �έR���vx鬵r��Cq;     0��   �K�R�����b�Z�_�A�     3 p   �Ҹ�����ףw�\lZK�S���[1     0>Z    p)|���R�F�F�{�v     `f|�    �»���q;�T#����pQFo     x��   ��Z��J9��G�7�����     �!�;    �AJ�����s�#��v{p����-      �E�   �������4-��!0#�n��Kq;     0c��    �-"�����\���۫O{��     ����   �����r4��Go��x���=�}1z     ��   paL편��c�W~����      oC�   ��P"��R�vsn���\<im����F�      x[w    ν��r���KO[������;      ��;    �Z��KY��\Go��X�6=��`�     �?K�   ��v�������w�\��V��     ��   �s�f)ˏrތ�sq�ZyP�a�H��      �w    Υ�r�^Z����zP��     �9&p   �ܹ���9�FX����zX��     眏    �+��|v����;`.��~�[�     �0�     o��V_�r:z�Ŷ�t���uD�     �]p�   �sᣔ�����4z�D������     ��;    ������4����{<���wo�     ���;    ������4-���L�����/{��     �]�   0[��z;�G,x�G���^�����[      ��   ��)��-�hʹ��s�ֽ'�-F�      x_�    ����%n�7<�u��֮��     �>	�   ����r��s���qk���v     ��   09��.�h!n�������֫�w      |w ����	  <�u)˫9��;`.����]���w  ��wߧ  �?� �ܶ۝Tk= ��[�,rގ�s�lmzX���  �L�;Q�UGG   ��#p .��s�lv��  �Y����k9oF8i�|#n .�֦�nR�;��    �4�  �Z��Z飇  _�rr=���0�������M��*��v/r�"�H�s-   �� �4z�9m�S�  ���9�~��j���Uk�~��v �Rhm��6�i:�����    �G  �R�S�lvB$ 0�SZ}Q���0���Z�w[ �I�o6WS�W�w�   �� ���b���)�o#  sq-��W�t2z�Ŷ�t�փ�� ��RJ�[ۍ֦>Mg�5w   ��|, .�����n�� 0+�)mnN���05"ݫ�pQFo ,�k�   p�� \D)m����������]{��9sΥ)�,K�H%.
�E���rR�q#�%Ҭ�ʲ7P��j�p�-��iP�j��m�4Ha�H� TFI�D��%)R"E�佤$�"M���g��sESI�眵g�������9��g�γh͏�  &f?��;f�3�*p�Eĩ�O\4n ����}���B�Tz7   ��� �,��i��7�v ��ٍ(�����p���r>q�5�  �������   ��� `S���6��%  ��ED�y>q<���^��'J�?�ڼw �T���RQ����H��n   ���M����� 0i��z�8�83n��8�����^hmѻ `M���~���;   8znp �Y��gɭ�  �5F�w�㋋ap�"\�T)��Z3� �:)j�i��b6;���   �-� �zjmH��<�� 0YCD�y_�1n��<]����  XW)bL9���[   ���w `�Rf��ѭ�  �5D�����rJ���gj��n���   ���1������   �A��u�b�����; ��v�8���ܻ��ZO��׻ `��:�Zǘ��GJ~\   b�  pEJc�Z�q; ���8�gn0n��<_��[����  �PC�y?պ�;   8� �����r�G��< �~bϽ~V�;`*��:{���;  6Y��V�N�V�њ3p   Xs�� ���0�V��@ `-�y���a�ػ��\��i�v ��4F����y�   �ڹ	 ��Tʬ�:��!  \�7Å7���0�k/�zp�(  �'���1������   �f���I�Z͛ ��x�0\��q<߻��b��㥜0n ��y�:�lv>R*�s   �+7�  xI)cZ��a �6^�ҥ���9���U��Rn(�� L��r�O���   �����RD������]�  �c?�Ս��Y�v8�/�۳q; �d��h����6�#%��  `��  }�6�j����] �F�)���q;(�Rn�1�n ���Zg���ڼw   ���� t�J��ZG��  ����r�lv�/�@��S9��h� 0u�弌a��0\p�;   L��; �C��j�� �YD�w��/��^�z���kͳV �uQ�<j�lv!�Tz�    ��E[ ��j��i���q; �ڙEԛ��řq;D��?�'r�?�ڼw  WmL9�Z�C   ���V! �ؤRfQ�h �~ƈ��q|q1�wLA��o���BkQ  �+�Rv��1��B���5   L����R��V��; ��7D������vx�S�,��u�w  ���y�y���6   L��; p�Z�j5o��� `�q<��һ���Rv��u�w  �'E)��ڼw   l;C3 �ȤRf��E��-  \������aȽ;`*��u绵.{w  p$R�y�,[k�k  @'� �QH)�y���\ �������aջ��ZO��׻ �#V�<��Z�   :0p WkCZ��5g  �����7å�0/�:�V)��;  86c�y/�6�   �f�;  ���Y�ul�C  �.o��o���;`*��:{Ҹ `���2�a�p!R��   ���; pR�y��v ����a���q�л��\���RNԈԻ �Nj�GkC���H���  �Mg� \�ֆ�Z͍� ���S���q<׻��|��Rn0n  Z#���ڼw
   l:C4 ���Rf��{  ��)��>����Sq����RN�w  �S��L�����   G�� �)�<o���C  �~�)�n���Xg��UDz����  ��V�"��ͦ   p4|� �NkCZ��� l�eJ��pָ���juC�� ��6���[k��!   �i�  W��1r���' ���(7�fg�ah�[`
JDz|���R��U p%R�V{Q�n�   �$~M \�����v ��1����g���N�|�q;  W!�Q�"Zb�GJ�c  �u2R ~���¸ `s��������:n?ךA  �6��"��֚L  �u2T ^]kCZ���z�  p8��v�8��3�wLœ9�im޻ ��7�����-  �� ���1V�y3n �CD�i�,���n�)h���omѻ ����j��Zw{�   ����] ���<�ֆH��  ���xfr����JY>��N�  6KJ)��E�6�0���Z�&   X'np ^.�ju�� ��r�8�9a�/��Rv�u�&  G��Y��Z{�   �:1^ �6��j�m �0?1��^?��0�Ժ�G�.{w  ����^Ժ�   Jm��    IDAT��� �vp�̼� l�7��?;{w�T<W��R�zw  �UR���J�!   ��� @g9�Sk~� ���4�<�zw�T<_��[����  `;�Z���x.Rj�{   `��� `{�X�a� ��ސ�ŷ����0gj�� �]kc����S   `�� `�:��j�w
  ���)]z�lv�wL��Z�ӥ��� 0C��.z�   ����I�̢�Y3�  �H'RZ�}���P��x)7� 01)J�M���  ����  �O�y�Z�7 ��L)�cϤd��j/�D1n `���-�C��H���  �)0p��b�Z� l���r�lvf0n���X՚-��(  SW����  @D8����ڐV�y�� `c-"�;���1�m9"=f� �IC��Z�v   �� �`��1r�7�v ��5��7�㋳a0n��(���W�.E��[  �*��y/j]�  ���`C�Rf�V7�  l�1��s_\C��S�"�t���� XS)"���T�n�   ��� 6P�y�Z�C6 �6D������v���q���O�mm޻  �W;��}�a8)yc   [�� 6K��ja� �ن�v�8�YC��S�"�ۥ�1n `��:k9�g�   l_�`S�6��j��`
 ��z�8���ܻ��;9/��u�w  �1D���5og  `k��h����� l�����êwL�wJY�qk��;  ���y/j]�  ��`� k.�2K��� `�e���vx�3��<[�q;  /ED���J��/   � �X�y�Z�5 �-��a8��a�ػ��ZO��׻  �S;��}�a8)��=   p� `=�X���  ���p���x�wL��οU�~�  ��Y�y?�   ��|��5�Z�j5��o$ `��>�K?1��{w�T��u�D)'zw  @O)b����ػ   ��; ��ֆ!�Y3n �
�K���g������jO� ����y/�6�   ��� �E)c�<7n ��)�n4n����u<U��w"  x�TW�e�u�w   w X��Y�:�� ��X��o���X�����r�� �I)E+e'JY�n  ��`( S���Gi  [bQn�3� ��Z+��  xm��#"�a8�Rj�s   �Z9�	K9�ø `k�"��g�`� �#��9�Ȟc ���u�rދּ��AZ�^���>���  �i�4�X�nn �����r����Kc�  X3c��8���ع�~���  �i|���Ii��G��U  ���n�3�a��[`
ZD����E�v  �V�呻����O������7zw  �&1p�)imH�ռ� l�!��c�,���n�)h�ũ�O�omֻ  �\���Rk��!��Ƈ��'~�>׻  6��; LE)c�l� �en�3�Ð{w���x���38  pXR]���֝�!����]�����w  lw ��T�,ju;! ���q��`�q0n�v){/����  �$����T�n��dCk���Ώ�����w  �;w �-�y�u� ��z�8�}�0�zw�T<U��9�J ��i�.���֚7��I���_�˿��G>r[�  Xg� �Q�y��< �2?>��8�zw�T<U���Z�&	  G��Y�y/���ȤK�R|����'>�3�[  `]�@)V�E3n �:?6�l/�x�֝g�� �8���x�褳g���������-  ��|a���j5���  l�7��7n��<W��R�zw  ����}��j��?޹��nw�1��  ��� �SkCZ��͸ `�~.�u��x����J���  �*E��y������o��������  �uc� ǥ�!�<3n �>'RZ�}��8S��RN��   ^��a����#7����+�;  `���1h������ ��~J��f�3���jO� �����^Ժ��jv����c���N�  X~� G��1�2�d��b�R;���"��q(�- �i�R�q6;�/A8�kMO׺\D��- ���)��&)ED�y7�c�q�ػ6���o{��[������w  L��; �V�,�:���Rjo�����|�z�|�� �f���9gzw  }|��ݧk]�� ^YJ)�֝H)�0\���&��/|�~����s�����w  L� ���Rf���w     �+e�J���(]���w������'�|�  �2w 8��Y�ո     X;��E+e/Z�Z8d�����]w�l���N�  �*w 8l9ύ�    �u�j��Z�F�p���|�ĩ/}��;  `������њ�W     `�Zg������y����~�{w  ���!h)V�E3n     6��r�OF�p�ҽ��������  Sc� �/��j�     'E-�}o���5��;�����G�Z�  �_>���     �`�����;6J�i������O|�gz�  �T���jmH�ռ�     �!E�{F�p�ҹs������O}�M�[  `
���ֆ��̸     �2)r�k��z��&���w�_��ý;  `
��j�6��     ��J)�e�á�x����]��  ����j��      ��&w#w8d���'�����  =���jm�����      �Z�{��y��)"��_�����ڻ  z1p�+qy��;     `JRDԜ�Qʢwl�TJ��{�W��{�  @� �#�Zg��      �,ED�u7j5r��r�ܘ����祐|�w
  7w x��E[�<�     x)"Z�F�p��yf�z衇zg  �q3p�W�j�i����      X)���{);�[`S�<���/�w  'w x%��4_     �JJ)�֝��p��:�����  p\���Zw�V]     �Q;8o�\8����7���n ��`� /�J�us;     �!(ea��#]���w����v�[z�  �Q3p��R)���E�     ��Q�"�b��`x��=���  p�� ��     �J������江��{{w  �Q2p�R���      G�����������  G�����JٍZ�;      6]�uF�p�Z��K_��S�����S  �(���J�us;     �12r�Ñs����㛷�~c�  8l� l�Zwø     ��պHF�p��/�<p�  8l� l�Rv��v     �NZ��T�N�Xw�O��������  p���.���     `Z);�#w�N�}�������w  w �F�uǸ     `:Z�F�p�j������?�я���)  p����4G     &�պ�q��\�8��������^�;  ���; ������CQ     ��j�9���ax�ٝ�����;  �z���R��v     �iK)E�y������#o����  ��a���uQs��     ����Ƚ#w��{�y�o��?��  �����T뢕��R�]     �J)E�u7�6���*���_��O}���Z�  �� l�R��;      �j)"j�K#w�v�ܹq8y�K�;f�[  �j��QRk�V�q;     �3r��7<����?��{zw  ��2p`c���5�q;     �����=Zs5\����������w  \w 6Bkm�rvs;     �I9/��;\���X|���ѩ�n{W�  �R� ���Ɣ�2.?�     `��tp���;��ŋ�p������E  X� ����9�q;     �&K��^�f� �`x��S���}�;  �J����J�%7�     l�9�5#w�&����������  ?�/} ���R�y?|�     l���M�.@���Z̿�����m���w
  ��@ �Ok)J��c      ['EQ��;\�t��0�<���g>�ӻ  ^�a  륵�X��S      褵�������3����so�  x5� ��Z�ɸ     `륈1j]��u4���������Ի  ^��; 룔e�:�     �D�:�R���j��w��}���w
  � w �B*e7j���      `bj�G)��3`�\���w���O}����S  �����Rv[���      LT��T�N�X7��gw.=��=�;  �����T�"��     �Z�;�V#w�J���+�}��w  |��; �Uʢ��u�      \���˓�*������O}�?�;  "����f��ݔR�      �DJ)Z)��ڬw����ᮻ�y�  �0p`�Z#�i;      W+ED伌���-�N��|�������  � LKkC���=     �5H��^�fW!�<���n��ӽ;  �n��0��f�     �������\�Tk�����ԧ�Ի ��e��4��"��	     ��3D�{��������ɓ'{w  �����Z�1��      `���,
�B�#����_����w  �����JٍZg�3      �P�΢����V�������ʿ�; ��c�@_��D���      l�ZQ�N�Xi�J����Q���� p���&�6o�z�     ��h����;`]������?���{w  �]�袵6k9��!      l�-��hm���b�����?���;  �� ��ژr^��3D      8N)rދ�l&�J��]w����o��w
  ���5 �Wkɸ     �ξ7rwfW �=;�|�w��  `;�p|ZKQ�^��     ��������?~�~����  `�p|j]Fkc�      �l�Z��#`]���߸����� �f3p�x���Zg�3      ���:�R���J\���<���3  �l� �T�N�:��      ���y���;���䓯��#w  ���; G*�6��z     ���Zw�5o$�+�8y����Gn�� �f2p��6��wS�      �RDD����ػ&��Ծ���ÏB  8t� ��R伌��     `���2Zs�?���3�O�����  lw ���}/|�      �~�Vʞ�;�h�����c�Ч{w  �Y8|��F�W7     ��Rk��3/����'�O>��7�N `s�p�R);Q�w      \�Z�֝�0u������{;  �� ��f�C>      6D-e'Z��K=���>���ݻ ��`���hm����w      ���6�n�Ik-Ɠ'��o��-�S  X� \��R伌���      `����2Zs�!�93{���ٻ ��g���9���      6��J�kF��o~������V�  ֛1" ק�݈�JF      6ZjmLgc��i-fw�����_k�  ֗�; ׮���u�;      �E��(e�wLY:{v<���_�� ��2p�ڴ6k�zx     �Vi��Dk��0e�o|�������� �z2pવ���y�z�      �1K9/[kc����b��W��ß�ԛz�  �~��:����2.?�     �-tpf֚33x��g˯~���  �w �N����      ��3�U�=���>��;zw  �^�r��F���      0	��R);�3`�Z��=����O��w
  ����+�ڬպ�      SRk݉�\�"���셓'��� ��0p�Gkm����w      LL���y��`��~�'������ �z��
���Z���q��      �CR��l�9S�W�Z������O>��7�n `��xm��F��;      &��1���`x�ً_��zw  0}� ��T�N�:��      k��y�u�;�j���~��[n�d�  ����W���J��      �B-e7Z�dx%�F����; �i3p����R�ˈH�S      `���h9�Ek����g�Y���_�l�  �����J�k>#      �����J���S5�{�O�~����  `���>���䕉      p]Rkc*e�wLQZ�Rz��ܻ �i2p�%��y�uѻ      6A�u�Z���)�x�������w  �c�@DD��Ɩ�$      ���w�7(�+N���o�~���;  �w "ZK)�eD��)      �aR伌֜��H�΍�G�|�  �����Z��3      �D�R�ަ�`��#�8���f�  �Ø`˥Zw��Y�      �d��y�uѻ&��H'O�WO}����S  �w�m���J�      �A+e'Z{w���'�N}�w  �`���ZK��2"R�      ��弌֜��|��8}���� @� ۪���9       �*E��ꀗI������w  �6l�T�"j���      ��T�<j]�΀���N��=��w  }�l����J���      [���h�n~�x�}���'?���  ���6i-E�ˈH�S      `��ݵ��^�������w  ��l�Zw���     �T��Vo_�0{��<u뭿ڻ �>��Djm��{w       �պH�9ǃ��5����  �a��ZZλ�3      ��rލ�l8�e��O�?����N�  ��/G ����,#"�N      ^Q����5gz�r��{��گ��w  ���`åZw���w      �ơ֝�0%�a��#��w  ���`�����E�      �G��,��Y������y�[���  w�M���r��      \��RD��֚=|O�1�����; ������y�w      pUR*e�;&�g�����; ��a���R�;1��       �Akc���;�d<y���?�?߻ ��g��iZ��]      ��j]Dk.���xqH=����  ���l��Z����w      p�R��9����#����������  �h�l��֝��v      �c:8""����{w  p�� 6DkmVKY��       O�u�Z����{�����  w�M�Z���)y;!      l�Cλњ�@�l�կ�������w  G��`Ժ��m      �EQ�n����f�����;  8� ��E�:�      �Z�5�p���?��G>�ӽ;  8|� k��6D);�;      ���r�m��z@D��*�G���;  8|�� �����zg       �"�Zw{G�T�������O��  �p���RvR��;      8F�μ���b���C�  ��;�j��Q�w      �A��֚˰ "��O�?������  w�u�ZJ��FD�      t�R)��5g���������zw  p8��M�;�6      �n���֝�0�����O~�w  ���`��6k�.zg       ��Z.ǂ�׾�3O~�#?ݻ ��g��&Zk)r���A       ""ED伌�#���j�꣏���  \?w�51�^���     ������0���O�~����  ��J����Z�w      0=��E�6���R�Q|��� ��1p���R�띂      �+I���+���'�xã��ٻ �kg�0u��D��      �W��8x+4D���׿�7zw  p������y      \�V뢵��,�����.O��}�g�  ���;�����      �J)���0�W���������  ���LT*e'"ܮ       \�1�a��^������w  �2�    IDATW��`�ZZ���      ��u�ل������蓟|K�  ��/3 �JYFD��      ��g���҅��G�l�  ���;�Ԕ��Z{g       k��1�5����W���ZU�w��v��l�I"d 	A�@0�0c�顙�p��bP��%DG	QB"R��"AJ�H�3�� "!{<���az�O�ϻ�֛��V��O{�z���<R��.vZ����]e��+�s�_���  <9w�U1�	      ���l_��aئ�:~��?Ύ ����Bjk�K)5;      Ѕzg	�6~����x�9  x2
� ����hm�      �G�6q�4��Z��_���  <w��2����      th6�W"�$͠��{ߑ~%;  �����\�      ��ܞI M^y巳3  �x
� �"&��Iv      �c�m�sI�����9p�+�1  x4w�DQ�tjS      �x����fi��R�/���9  x4w�D5b_�,      �cT#6�C@�����<������  <�R%@���l��      �41�m�}m���_��  ��ya�2��w�      �d���?;�z��w{���ώ ��)�dhm��2Ύ      Pk���2կ���3  �`
� �Q�l�/;      0\m:�_"\:�`�.\�<��O�Qv  �2w�%���+��P      ����;�K��׿�\:4�� �_���L���fv      ���f�g�,�K�6N|���� ��H�`�f��V�      ���R�t�?;d����OǗ��6 ����,��>�      �3.��[��z����7��s  ��)�,CD-��(      ������Q3X�W^��-�  �C�`Z�_���      �bꝙ&R�rer��W�gv  nSpX��Iim#;      ���l����e���?��?  ��)��tj�      ��j��N���s@������W��߳s  ���X�mV�Z      `=�kkJ������8tȌ  ���D���fv      �'��f���9 ��ҥ���'�5; ��)�,Jk�K)>�       ���ΐM��͟��  0t
� �1��6�c       �Tkm3"��9 ���ō7>��?�� 0d
� ��~��     �uTK)#[����/��� `���Fl�Rl3       �V�6)���a|�������9  �J�`�"��tj�      �����%���R}��/eg  *w�9��m�V      ����2�s��~����� 0DJ� �Q��;      @b6۴ŝ��x���� `��極��v      ����ھ����=�����of�  w�y�Gk�1       歵����a����� `h��a6�ou;      УZJ���@MN�|����� `H���Fl�
      ��Ek�1��KQFG����  C���5�S�
      ��M��K�˭�ё#:���?�� `(�����Y<K     �aՈ���t��v��e�  
�L�݊�q��      01�m�����^�맟���s  ��;�.����R|�      ��ޙ� �[��ӧ�Wv �!Pp؍�Q���      `٢����9apꫯ~��/|�d�  蝗�ݰ�      .[����룭7����  �Spء���      ٝ-����l����q��$; @��v�����v      `�j)e��fvX���59����Av ��)��Dĸ���      ��Ek�wh��+�eg  虂;�N�f��#       �3T��;����>��9  z���"&�       �#bn�fp�����  �RpxR���       ���ff���������3?�� �G
� O���R���       ��׈���T���g��^v �)�<FD�2�mf�       XU͍�����?����� �w�Ǩ���{^      <D-edqCS����o}�d�  ��&��DԸ]p      �jk�Q�s�2�_{��eg  荂;�#Ԉ�Z�0       ����b��ҥ�ѧ����  =Qpx����      xr�m[�����Rv ��(�<Lk����       ;Q��Za0Fgμ�������9  z��� ����      `�a�;�Q�����1  z��� ��v      �ݲŝ�>����/���  =Pp�_D��      v�w�f:�����  =Pp�_���       {Sk�fvX��k��@:4�� ����Q�lf{;      ��l�i�;CR�^����sv �u��p��lo      ��Z[�ŝA�8|�`v �u��pWD-���      0'њ-�J=s���z���d�  Xg
� wԈ�b{;      �<�b�;R#���''; �:Sp(������*       �f�;3:|��g���wf�  XW
� ��v      ��ŝa�yst��7�Kv �u��`{;      �BEk�a�;2>z���3  �+w`���M>�       ,H-�V[����Oy�/d�  XG
���E��      `ᢵ�b�;QK)�';; �:Rp���v      ����������>��=���s  �w`�"���      �g6�ŝ���n��+�� `�(��5���      `�F�wd��?; ��Qp+f3M       �,f37m3�s���x晗�s  �w`�n0�      X>[��v��gg  X'ʝ�0�X      �&�S[���c������ �.܁���I�g�       ���-�1��w^����1  օ�;08�5�        ���/;,������  �.܁A��q�f��       C�٤D�0o���Ƀ?� `xI ���Yk͎      0x�V7p35�LO��w�9  ց�;0��f{;      ����6J�-e����OġCz  ���GľR�#       ���[��k�����O'; ��Sp�!���l#;       Q�f���3�ȑ�3  �:w`Z�,��      ��Z#,,cF'O���/}�oe�  Xe
��0��c      ����l3;,Cm�\;r��s  �2w�{w~��y      ��F%b��at��eg  Xe
�@�b:�K      ��پ������~���s  �*w�kq����       <Z���]ar��W�3  �*w�k�5��      ք/C1:z����K��� ��܁~E�b6�d�       �ɴ�6"B���ݼ9:���!; �*�B t���Yk͎      ����a�;�0:~�@v �U��t)"j����      ���6J�mft��:���{��G�s  �w�K�v��      ��Sk)���hu:�������  �F����       k+����������  �j܁�D�K)��       ������6:{�]'�{���s  �w�?��%?      ��3�eZ+��g�Sv �U���%���&�1       أ�&%�fǀE;�w�3  �w�/���      �����3�ܹ�Ǟ���9  V��;З�6�#       0'f�@-����;; ��Pp�1)�k       =ݙC�FǏ���  �B臫�       �f�@���8y����s  �w��hͯ�      z��$"t\�^;q��  ����Bmm�f�       `�j�=���V��Xv �U������md�       `AZ�(��ѵz�����>���9  �)��/b����>       }���IvX�ӧ��  ��;��f3��      :��fvX���?�  ��;��"b\Jg�       `���q��u�k�ڵ��<���9  29�kmԚ��       Pk-�5[����ԩ_��  �I�XkM�      `8Z�dG�E�8��  �܁�1����       ,ͨD(�ӵz�����_�� �E�X_��      7}3 qꔂ; 0X
��z����qv       ���I�p�7]�'O~Wv �,
��Z���,       ����N�F�/O?���9  2(�k)Z�dg        ��;0:}���  ܁��1��      @�q��{�k��'?��  ��>�v�_�      ��it������� `�܁��Us       �lfvL��o���  ˦���Q)�RJ��      @�ZJ-���H�ӧ�;; ��)�k%lo      ��j�L���N<��g�  X&w`}D�hͯ�      (���MJ�[��WDi�����  ˤ����6}�       ��F��N�N����  ˤ���p�       ����,���Μy������k�9  �E�X��      �_6��qvX�:��o�����9  �EYX��      ���IvX�z����  �E�X��      ��lfi]�:���  ˢ����W�y^      �0�;�e�R�qct�g~�W�s  ,��(��jk~i      ��E�-ӷs�~%; �2(����Iv       V�lf�L�N��Dv �ePpV[�$<�       x�Q�g��E_��y���$; ��)�+���      ���mdg�E��=���3  ,��;����       �PX�F�Μ���  ������I)�f�       `m�J�8;,����wŋ/>�� `�܁�e{;       ;e�LϦ�z�ԩ�ʎ �H
���ru       ;
�t��;w ; �")��)bRJ��1       X/��zg�]�9��  I�XM~Q      �.U7�ӱz�������  ������Z|l       `��R5zQ��ʎ �(
��*�Rjv       �V�����ٳ?� `Q܁���       �Q5{�c��7ߟ� `Q܁�Ӛ_�      �7f�t�^�>:���(; �"(�+��q5;       k���qvX���ۿ�� `܁�R��      �y��Ȏ �2z�����  �
��jQp      `^f33h���[O����d�  �7w`uܾ�s	      �y�sh�Tg�z�ԩ�� `����Qmo      `�Z�Ȏ s��g�#  ̛�;�2B�      �93��g�����  ��������c       Нq���!`!.^�<��ߝ `�܁�P#6|M       `�����ӥQn�?���  ������1      ����̤�V�;���  �I��QKk��       t��I�p�8]�g�~8; �<)��`\n�
       �P��l�3�ti����Wv �yQp򵶑      ����&�`jke���d�  �w ]��       ���Mӳ���Tv �yQprE�k)5;       ���qvX���o8; ��(��Z�Ȏ       �0�[���ŋ�^��_�Xv �yPpr�u<       K���;]����s��yv �yPp�D�hM�      ���R�%�f�E������  �����Lj��       �娷���N�Ξ�Hv �yPp�Dk>       �Tf��jt�¾#/����  {���im�      �a�f����R.^�Jv ��RprD��g       K��"Bɝ.���"; �^)�)j�+�       HQ[3��K���#; �^)�)B�      �<6�ӧ��ʎ  �W
�@��|,        Gk�Q�c�����z����g�  �w`�"ƥ
       �R�w:Uϟ���  {��,]��dg       `�jkf�t�^��3  셂;�t�G       ��f�;]��ν/; �^(��QK��       ��R�%�f�y�[[�>����� �[
����}        ۝ٵmt�F���˿�� `�܁���M�3       @)�3l:.�Dv ��Rp�*Z��w       VC�6]���ǲ3  얂;�<5|       `EDk�Q�s�ܝ?���  ���,M-eR��       ��Zk��L�s�����z��g.; �n(�K��(       �ji�M�t���K�8; �n(���        +&̲���Ofg  �w`9"jDx�       �R��q���9`�.^|v ��P6���2���        VK-wJ�Йz��f<��� `�܁�p�       +jd�M��tZ��f��� �S
��RD��       �$��U�|��3  씂;�xU�      ��e�;�]����  ;��,øf'       �����6zt�·eG  �)w`�Z�dG       �GRp�C�K��eg  �)w`��Un       �:w:Toݪ�<�Lv ��Pp�z�       ��,o�S�[[/dg  �	�S`�n�½f�       ����m��.^���  ;��,Tu�       �c� �mt���3  섂;�P��      ����̸�N�x��  vB�X(/�       �3n:4�y���쳟�� �܁ŉ�%�s      ����KD���y��/dg  xR���"�k��      �z��N�:S��~ ; ��Rp�Fx�      `���̺�N\����  ���;�0��      ��ѧ�?[[�ʎ  �ȁ�	�j      `ݘuӡ��˓8xp3; ��Pp#��Rjv       ؉(eT"̻�J�V����9  ���;�(~�      �ڹ�lש�;uk��  ���8��M�#       ���yӣ˗�Nv �'��,��       ��̛�ԭ�eg  x��b�6Ύ        �ҚNݩ[[���  �$Ɓ���Q)�f�       �݈R�%�ܛ��+W&��K��� �8
���U�       �؝f��7]���7����  �� �]�gg       ��0��G׮�tv ��Qp�/³      ��f�M�.]���  �� �]��W�       �5�o�t���#  <��;0_5��      ��7����nm=�� �q�P�y���      ��W�n�]�:�C��] +�a���6       �`Nof�z����d�  xw`���=       ��Э�;׷�?�� �Q�j�s      �.T�:4�r��3  <�C80o�+       t���s�3�z���  E��QK)5;       �C-��۳p�Ǖ+�͎  �(
��ܴR�r      ���Y8��r��  E����j6       :S#�k�����q:�� XY*�<y�       �w�3����g?� �a���i�3      ��D����Nm���  F�'�       �b�;�]���  �����B_�s       ���aNW�W�~4; ��(���y      @����˕+�͎  �0��\TW�      Ы�qv��+Wޑ �aR��Pp      �cf�t�^��G ��r��"<O       蕥ot�N���s�}ov �q��5�       �f�th����3  <��7�w�w       zUK��`ަW��Pv �QH�,Jy�      �c�D��Еɭ[��  � �����:       �gCW���fg  xo`�ZgG       �����δk�ޓ� �A��=��      ��Uw:3�v
���    IDATmv �q��,<K       ��8ݹvm#; ��8x{ךg	       }�p�9}�ys/��Tv ��)���%      ��E��ЕQN]���  �s��$n��+�      лj�;��u�Əeg  ���;�'�s      ��0#�+q��'�3  �ϡ�W�      0��ћɍ��  p?�n`OB�      ��h͌����Wߟ� �~����Rjv       X3r�2�~���  �Sp�$�:      ��]zs��fv ��9t{b�;       �њ9]ݸ1��  p?w`���      0�6�e{��4 �rP�݋�E�      ��wf�Ї٬����3; ��܁��      `P¬��lߺ���  ����Z�      ``�����͛ߟ �^ʩ��Ek�!       �Y9��y��  ����^�~�      ��T�r:3�~�#�  ���^��v       �Ŭ��ܺ���  �Rp��K;       ��6��ƍwgG  ��7�{�)�      0,f�t�޸�Tv �{)�{�      ��(�ӗ76�#  �K9ؕ���      �A	}:3�qc�� �^��n�Z��      �ZJ)�ё�uK� X)'��TW�      0P��ӓ:�ַ���wg�  ��a�-w       ��̜�ܼz���  �Rpv�Fx~       0H#w:Ӷ��'; �]
���D��u       )Zӹ�+��>�� �.�m`W�_�      0\f�te|��G�3  ܥ��JxY      `���M�y��  �Rpv��:       CefN_f��eG  �K�؝ּ�      0H�sCW���{�3  ��얂;       �f�tet��;�3  ܥ�얗u       ���ә���?; �]
����5:       C
�t&n�ڗ� �.w`�"j���      �Z������Fv ��܁��      ��)�ӓz��8; �]
��nxI      `����h{[� X&���:       CW���HL�zd ��p0vl�%       �u6� V��;�s^j       4��ӕ�J:4Ɏ P��;���       f�t�o}�C�  JQpv���       �2)��  JQpvA�      ���֌��ʾ��gg  (E��/�       ����y�և�3  ��        ;V��p������  �(���-      �A��s���  �(���       �/���fg  (E�؅hM�       �#m6{Ov �R�       `7,��+u6{Wv �R܁����ػ��F�,=��8�KDV��=�G��XcdR���"�� ��� +KU]y	�q?��Y������       Б� !p.�w       6����Lӗ�  "��xI      `�2���.�; �w        �T)��ѕ�ֻ�  "���#�       l����V- �J���Ru;       @gjݵ�  !p.4Ex�       菖 X%�E��}�	        \Y֪% �C	p��xt�       �3%���  !p.Tw;'�       "J�ӏ�; �J����s       ��l= �h�	 A�        �q��]�  w�B;�       �S25! �"�        6�F��E�).�       tgp� X�;p�����       @ojՄ  �����n�z       ,Cq𚎸� ,�����e       �?� `!�� ���bl=���a���Vc(%[o    X���r����-�)|� �&p B�\����<��C��+    0�/�0}��Z� �k�10})~��e���׺       �n ��܁��K�{       ""2[/  ��U��LӮ�          �$p.R]p      ����z  �H�
\�n�;       ���  �K�\�m��       �z   tH�\��7        ��  0�*p���          ����Ȱ���       �w�R�< �A�
\�8���7       @k�� `w�"%��       hM�  ���2Zo       ��2[/  �.	܁K�{E      `��wzS�H � p.�9x�      `��  0�;p1/�       l]I�N_�D K!p.Vjm=       �� �,���Jq�       �#�� ,���\��      �M��� ��        p�R��  f p.�;       [Wk�  �%�;�w       ��g����� �A�\,��      �u.�ӛR�� ��;��
�      �:���?� �R܁�e�w       6���Ng��A �e���      �q�g�  0�;�^�      �4��� �B܁�yI      `�|v  ���Z��       `�j2��
  �H�X��wR      �Y%��;  �B�\N�      ��e� o �y܁�MS�       �L�:�����u ,�����       lX�,w  ����XN��      ���L�� �L���J��'       @Kw�R�H �!p>$k�f      �6��  ��2�kt       6�Q8  �������      ��*w  ��@�_�      �F	��N�# ,�����u�z       ��w  ����/�       lTN����� ��܁��      �QC��'  @�����      ؠR�w:��  ��;�!9M��       ��2b()�3ŝC `9���LS�       p{�C
� `6w�C�8��]       6'kB�  ��3���:       [���m�Kq� X�����      �M)�>+ �	܁+~�       �1w��; �0�T��2�      `Sr}V  3��|X�u�z       ��49w  3�Vj��      ����M�# ,�����&�C       ،���4��W�w `aĩ���q�;      ��"���z\�� X�}�����w       6�ֺ�;�q� Xח���y��      �fdwz�' X�;�a�V_S      �v��cr  ������u�z       �B���З�o6 ����|��w       6"��g�  03������       �0��]������Ӵk�       nB�  ���R���;       �+�1M�g�U�� �	܁�9��      �{�+��g�U���%�������      ��M�.���w `�����q��      @�2u6t'U �y�>�K<       ����q  ����e���       `Neu6  p��ϛ&�;       ]K�;�)�� �_���<_�      @�ql=�K� ,�(��<�]p      �[��]��z  l�������       �Uk݇��Τ� �B�R�O+�s��l�       �Pj����; �P���ˌ�2      @�j���  `+��U�L/�       t�����; �P����iڷ�        �G�  ܈�o�*r]p      �?��8�[���r� X0�;p�t��      ������ ��	R����y��#       �ڦi�q  ��;pe�z       zSkݵ� ז.� &p��dz�      �+e�5t���� \M��u       :�糾��� ,�p�jr��7       �5��Y	  7$p���N.�      ЏZ�1M�W�u�� ,�����q��l=       �!�i�cp  �%�;p=�X"�      ЇZ}�9�q� X8�;p]^�      ������?w `�<�W�Ӵo�       �B�N�� ��y�k]p      `�JD����;)p N�\��(p      `��4��4��  �#p�*ܳ�       ��R�o���v `��U�Z#�n      `�r���G� ����iڷ�        �r:	� ��;p}��      �U��IWCwr�c ,�'��N'�;       �U�~��+  `�����CDd�       �9M�L{ӡRZ/  �Cw��Ʊd�7"       V)kݵ� W'n VB�̣�}�	       ��t� @#w`�(p      `�N'���� �J܁Y��$p      `}jݕ�Y	Lwr�� ���Ey�ED��       �u���n��6 ����8�Kz7      `e�8��r��E� ����M�&/�       ����k=�N� ����M��w�7       �%�񨧡?w `E<�����_�      ���c[�  �M��y{�gD��       FN�>���th�� ����M�5J��      `��7�ӥ,� `=���r�Zo       �?�x� @cw`Vy:	�      X����񨥡?�� +�����>[o       �?P2�1M�g�ե� X�;0�r<%B�      ���4��r�T� ��܁�e��'        �v:�ZO�Y�����;���'       ��:u4t)� ��x0f����      ���Z�y:��鏸 X!�;0��a���3       �WM�^L�� �
	܁ٕZ#3w�w       ��G�iӥ� +$pnc�ZO       �_���o=f!p VH��D�w       ��:��QL�� �
	܁�8���g       �߫�t���l:$n VJ��D�ޜ       X�qܵ� �� +%pn&���       �{y<�[o�Y����7���]�       �7��xT�'�; �Rw�v�}Fd�       ��E��W�,R� �����2�^�       X��}�0� �bw�r��[o       ���x��'�; �bw�����      ��j��]L�r�� ��I���p�GDm�      �m�i����3`.� +&pnkK��      @c9���  �&2no�[O       `�������� 	 ���ps��v�K�       h%k���XZ�9d� ������ᮔ2��      �6�i��t��N	����7Wj��ܷ�      �F��>��_w `��@y:=��       �F���ZO�Y���܁6����}o       ��4��tR�'�; ��;�Dy�EDm�      �m��t�z�%9 �~�h�62#�O       n����`6.� ������       6����^�>���Nx`�9�JDm=      ����>����� ��h��ϥ�=      ����y�z�F� tBX
4���C�       lCy{�ӭ�` @<� m���ED��      @�j�����5}r� ��h�翎��g       з:���7�l� @G�@S%3�V�      �Y�����`6w �#w�����![�       �g����d�V
���xp���R��z       }���>km=�#p :"p��R3��g       Ч<��Zo��0 �/�n�exh=      �N��:�F�\o :#p��p���      �u�zWƱ�
�M
���܁E(�㐭G       Н<��Zo�Y	���܁�Ǉ�       �Kw�5ȿ ��x�#���p�      ��uW�G���� @���b��a���;       �C��}�0+��y��#3rZ�       ���]�	0�R"[o  ���X�<�|      �Y��!�޴1����  f�!X��׻���g       �n�o�w�� 蓧`QJf�i�q       |Jy��3]K��N	܁�����l=      ���u��AC��� @�<���//�����       �)��>�i5:&p :&p��1M�*      �ɷ7�9ӵd_ @�<� �T��#�      p�����a�z��w �cw`�����0L�g       �2���s� 蜧`�J�Q���;       X�����`V�� ��������      �?���î��S�� t���X��r���;       X����Hw���� �܁�*�����z       �oo��7��� �܁E���1"�y=       ��֡Z�6� ��X����O�;        ��>����-]p 6@�,[f�8>��      ����'��\o 6�S�x�����      �J�C:��z; ���+oo;u;       ������ޥ� �Fx�V!O���       X�|}�o�f�z; �!w`���}D8�      �?�Z���]�K�\o �ē���N�      �?9�\o�.� "p��x|l=      ��y}�k=fU�� ��;�//Q��z       ː������o�v `c��z�NCd��      @DD�����`v�T �O?��Loo_��       ��Z����o��.� #pVex~��al�      �Ʀ�>jm���z; �A���u��R�g_1      �u��ώ�� � O@����뗌��;       h��]������  ps��)���"p      ج<�\o��v `���*�����       yy�k=f7H� �m�����c�2��      �m�4����5�K�; �Q���u:�KNӾ�       n�pxh=fW� �]w`��/��g       p#����k=f�z; �a����ʗ��(���      �m�8>D������$�VɌ8�[�       �6�����])�� �4�;�j���K�p�      �w�tW���z�-]o 6���j�x��2      �������	�; �q���իoo_|5      @�j-���o=fW|I ��X���t_�al�      �y�4=�Z[π٥��  w���<�}      @�^_�[O��� ܁>��˗��Z�       ��j��ۛƅ���z �"x��P�}��      Н|l�n��v ���=9�FD��      �Ք|z�k=nB� w�#����0��      �u��鱤;gl@).� ����F�5�x��z       ��Q���[p� �o<]�?�f)��      ��4���TZπ[H�; ��x2�R��R���       >'__[o��(�� ��	܁�L//_��o�      `�jݕ�W]���]�	  ��E �����o�      ���ǣ��l��  �@������       +Tk)��w�g�M�- ���Х|zz(�L�w       p�Ǉ�|��F� ��'$�K�����W�      ����}�	p+YJ�	  �#p���Ǘ���g       �'M�]���Y��� ~��$�_����Z�       �Oz{{h=n%�  ��Sе|}���z       ��!_^��g�M���?  ����Zyy�+���;       �}y:=F�_�F�� ~���^=~
W�      �������ݮ� ����+OO1c�       ��<�b�Zπ�?{��    IDAT(ŕ> ��!p�Wk���C      ��Ɉ�����;�V��v ��%p������w      �����!N��z�L�� �{��6�c�����       �Qy}�Y.�1ȵ  ��'&`3�?e)S�       �U�w���_a3R� ��<1�Q��!���       ~V_^��� 7S���  �]w`S���OQ[�       غZ뾼�jW��� �OM�������>      ����[O��Zx���d�  "O`�������R      �H�u���}�p3�,?T��z @��ؠ��r�z      �����K���p=�]��� �R܁mz}���       Z(���0��������Rt �"܁M����      �\�_���3�v��$Z�� X��<=\WɌx{s�      ��2#���[π���Z/�S�pe ��;�Y������      �v���2��W�픲��{EC ,��جRk���e-/�       kW��Zo�[ʕ\o��Մ� @����}��e�s�       ��q�/�si�n���G>�A� ,��ش2���N���       �OO��w�M�K�� �"��)
�������a[�       ��4���Sa[����z @�� ��\�tz�g�       ח?~��ζ�YJ�q X
�;@DTW�      f����z;��۵^p��; �^ ��+�y:=��      p=�������]o��(�ݩ� ��;���o?��      p=y>����+��/��z @���o�8��      pE����v6'w��>f�w� X�;���o�~\q      ��:����=k��e� �"���
`eK=��d��      �����v�gŁ{�c�  w��߾}-��+�       �z;�TJd)�W|X� �E�(�X�w      ��p���Z�����2o�7  D�~ݷo_�0L�g       ����lT�<p�axo=  B���~����;      �e������������� ��;�o����0c�       k���P���z��꯷GD���o�  w��6�����      �Y?~������������ ��;�������;      ����!N�*_��n�z�u���  !p�}�X�x��      ����xzr���)%��������O�  w�?����p�      ෝN����E9��_������ ��;������_�w      �_���C�	�DG��������  "� J~��%K��w       ,M���ir����(n/�]��w�n ,B?OY 3*��//��;      �_e�%�p��M�ݮ������o� C��'���os       �_�_Ku'���z{DD��I" ����I`^���/�;      @D�P~��k=��-p�� �bt��0���r�~w      D}}���3TJd)�W\����z �/D� ����_"bj=      ��Z���y�z4�۵^puywwn� �w�K����4��=      `����k��D���#"��N�'  �B�������a��\      ���4���9a��N����ZO  �E�O\ 3;��<�3��      ��zzzl=Z�N���� �����o?���w      `3�|~��w�	��i��wwϭ7  ��ߧ.���c���O�;      �?~���f�n�z�|���'  �B��?~|�a�Z�       �[=���\Z������/_��� �_���0�Rk���_"���      0���ZO�VJ���#b*�?Zo  ���ೞ��0�     �n����R},�FCd�3����n� �w��ʌ�Ǐ���L��       \]�C|�~�z��C��������  ����� n�����4�3{��m      `K2"���O�w@3����s���� �_����?���ײ������־���3���!Eʒ)Q�2,+p�H2$Y���YQ-ܦA�(X�@�]((�-(3R,�I��i#������k(��N|��h�\���s����#�C�C���ۗ��'5|�2:k��ٿ�����z\�      ��L&�tpP�΀b����n��G�x�F� �0p8)��U>:�ǭC       f���R�(&��pz{�zM� ��������U5)�      𠚣�~/���`No��ȝ��� S�����������      ̬�4)����;��E9�="R�7*�  p;w��6ts�b|�      ����Rj���[���#"��;,�  p;w�Ӱ���S���       �gMS�`�.��,���M��_� �v� �a8��x��9�.      �k9"�`�\���lR��n�N  �݂]���fss%���t      �]��qxhO��J)�ܛ^o�t ���j���85+q�      ���#R���l�Qw:�)�  p�Ż"8Ci{��      �,�y4J�3��E;�="�i����  �[�+2���s4����Ҥt
      �5M�۝�PT]�.(����t ���NY��k�ɤ����     ��#���[�4Yp�xz{���^��Kg  �n�� �^��\Ku=*�      �C�������j������G�ۤ�^;.� p;w�3�F���Kq��      ���#"���Kw@q�xz{D4KK��  o��Wf %ln.GUMJg       �i8���q*�%-���KKG�  ���������E��;      P^�T���-��-�����=(�  �v�{uP@��m7�I;�      ]΃�rdO/Yp�|z{DD��S: ����X��\����       W3���p������������W: ���
���8����єN      O�H���/���E?�="�����	  og�P@���5�t      ������dR��J)b�Oo������  ��U@!ys�\��q�      `�4M+�v�(θ=""�n��n  x;Wj �����9:�GD.�      ,�fkk�t�Rd�Hu�������  x;Wj %mn.GJM�      `���q*���.�0���I� �wb�PR�D3�E��;      pz���[[��P\J�~��tT: �������y2i�K�       s(GD3��g�����4����  މ�;�4��\����/      ��F�txh#No�����	  �ć�i0�|p�M�      `~䈔����;`8���r����  ���`J���^��      ���9G��_J/�����~�_�N  x'� �ds�\��Q�      `��J�A�tL���������  ���`����j2.�\�      �q��˥`*T����&G�vοY� ���L����H�)�      ̮��p9F#�^��5p����#o�q�t �;q�0eR����SU�J�       3�i괽�.�S��";������N  �w�i4����R�z+      �]��lm���i��t�tZY�+�  p'� S*ol,GJM�      `v����t|�j���L��$���,�  p'�� �T�9������ƥ[      �闛����ۥ;`Z8����KK��t ���L�ttT����$      pGyss�tL��wW/-�^� �;1p�ryss9�d�      �Q><\J�Q*�S�2�z7���_J7  ܉+9�)�r���q>�j\�      �BMӊ��N����*�0���|��ם� L-w�����8:�G���     ���[[˥`j�t�w�WVF�  ލ�;��h66�#%w      �M��p)���y��t��kVVK7  �w��r�fs�|�4)�      L��i��v�tL��";��=嵵��  ���`����GG��p�;      ,��#om-�΀i���~W���*�  �n�fL��\����      @9�p��ǎ������ߕzy�wK7  �w��r�fc�TU��-      @MS���N��*No�k�^�WK7  �w��������rD8�      L��\)� �$�u��3"w����_�f� �wc�0����R���}L     �E�#���_��(�n��R�@ݵs熥  ދ�;�Y�s����Tף�)      ��L�i0h�΀i�[��	3%��J7  �w�Yv|\5{{k1)�      ������r��*)���]�kk�)�  �^�f\����ɤ��H      ̟�wvVRӔ��t��I���,�  �^�����ZT�S�     `���~:8���U����ø��ǥ  ދ�;�<�LR��}>�d�      �i����΀����{��*z���t �{1p�i���݈ȥ[      ��#"oo/G�n��ڃ�����FO��/��  x/� s$ol�4�#      �����ȶn�RD��}9~�t ��p�0GR��"�I�      ���ɤ���ۥ;`��.�0��s�]� �n�̙t|\僃���      3*���R��:)����YY���	  w��`mo��i��m�     `��ȃ�J��V��6No0���_/�  p7�����ZU���      ����ǽ�߷ⅷ�*��?�V+_{���t ��0p�W�q��윋�I�      �.�\��f�tL#��?�|��qz�5�� 3��`����v�;q�M�      ����lo�����]n�J'̼|��v� ��e�0�66V�)�      0�rΑ��ph�o�ҭ_<�ɹsV� �n�`0�&���QU^5      Өi�i{�S:�Q���	s�^]�?J7  �-w�����fww5Rr�;      L�Ԭ�/���i�����'d�����  w��`A���;�:�K�       ����ժiJw�trz����~�~�wKw  �-w��66VsJ�     �h��ph��ĸ����K7  �� Hj�����"b\�      Y�L�i{�S��RJ�+����z軥  �+A�Es|\�����$w      (#�����0����OTu���]� �^�,����q'"r�      X4ykk55Σ�wTU)���+yu�WJ7  �w����W��     �l��å�5��������n秮^���  ��&��r���8U5.�      a2i��v�tL+����<��0���]  0S���q���E��     �iʹj�חKg�Ԫ���JW̝|����  ���`�������ND��-      0�����8w
����"�?�/J7  �+w "���dw      8��p)�6p'u��)�Ν��  �O D�9bc�|Tոt      ̓<��c{�S��VJ�+�S�j�'�}�(� p�\p��q����&�'���׿     ��)��/��i�=�>5���k���  �W� �)�4u��/�z��T�t      ̪yss55M��^U�R銹�.\�^� ��a��[�kk���W��ou�_o��     �Y�#"����ё]�IJNo?e����t ���A
����r���^���~��[�W��      �{���{1xc2����W]��F� ��a����G���Ո�$彽^�����g:����	      w�i괱�+�S��"��Ч)w:����z� ��a���:/�q�.�hT�ᰓ������N�h      L��4�Y__)�S���y����  ������H++��Ї����ѨU_��z��L�7�     ����;;�i2�P�M]G.ݰ.^�v� ��e�@DDt�_����ٶ����z�����?�:�2      �n9"���r�0�ݤ����L���n� ����H�v�?��;��yw������J����{W      �&���N�tL��r��Y�;�ߗn  �_� D�������U��Ij��zQU���O���V      ""��N����0�r]G.�(VW'�~�+��t ��2pXt)E祗�����f8�D����S��F�      ,��4)ol�D6ۅw�R��L�4/n�n  x�\�����Cw7V?<lE�T��s��S?�7       X`y0X����P�^�t�B�/�a� �a���:��rO}�9"�W���O~�}JY      0�rΑ���������|�,MΟ���  �-�V?�xԗ/�󝄼��M)5�_l�_|�um      0��hԋ��A�{I)�7���v;���~�t ��p	��:?�c��/�LR��׋���'?�j]��}r      ,�����f�t̂\{�|�&/��^;.� � �Tu�\��{���Ѩ��a'�:�?�v}钟)      ̵����J�\:�^��t�/�A]��g�  �1"����rDz��	���<שӉ���v��w'      �K9"bkk5�c��ཤQ�%��/^���  ʕ$�J�n�?������n7"�Z^����I�����      0Er��_�����B���	�)��}����  xP>x,���/Ft:'v�D3�"�\_�T�>�َo�     0/rΑ�å4�J��,�u}�w�\s���ʗ��G�;  �"�����\�~��gӤf0�GJM��պ�?�w      �C�tbk�[:fBJ�@��.]�Q: �$��X0�| ����]~2Iyo�)5��~��~�E'X      0ۚ��7o.�΀Y��t�Bky�wJ7  �w��y����G�*���R���'[�k�ܽ      `&刔76VRΥS`6����)�:�˥  N��;���~:�G=�;
���<������ϴ�K���     `�ln��xl�w#�ȕG�%�s�FW^��Kw  �W� �{����&��ur�)u:���N����      3!GDV��Ȧ�V��ޥ�G�Y� ��0� ���~�3��5�A/GDZ^N�/|��:�3�{     �};<\��}k]�[u99󬸋���	  '��`At^~9"���*��#���""ח.U����N�}      �X������&�[)E�̏��������  '�&�HKK��Ї��o<�����M)5���u�ӟ�o�     0��ɤ�76��;`��V�t�WW�׾��,� pR�@����V�̲|4����nJ�i?�\����h�      �;ɹ����s����=5�#�l�n  8I� �Պ��/�m�����󱏵:ׯ�?      S!G�fcc55M��U�2;��.�~� ���J`�u^x!��r���o��ߎ��RD�}���?���      �#"��W�hT�y̐����rx���(�  p���YJѾ~�tś����#"R��_�K�֕+~     PJ����qxh�����ӤY[?���s� ��dX0�Z�<�ŋSs�D��<�rJ9WU��s���%?�      8S9��GGKi0h�n��RU���<�&"���t �I3*�c�W^)��Ú&���U�D�����ک���     ��������0SR�\{����\��OK7  �4w�9U?�h�W�L�p|2I��n?Rj��r��j'z��l     `�L&����/��Ƹ}
������t �I3p�S���t»J�q����H��.\��^}��Z��Y      ̳����7WJg���u��Y6m�GϾ��?/� p���PZ]��>P:�W��Rj���z?�S���h     �4M���WRΥK`����N���cV� �4���C��_�������pX���vD��3���O}���      �����%s�    IDAT�jL&D�=���=������  ���`Τn7:�H�{����y<�SDn}���'>�.�     �|�[[�q|l��ȸ}z���;��Q� �4�̙��?����͹��N�4U�ȝ��[��^r�     �����#�^UUx���j.]:��o�(� p|��'U���KWܷ<tsD�������:/�P�n     `6�����i�3'�W)E��љf�c�}�t �i1p�#�矏t���~�>ED��Ӌ��SJ����v����5     ����p)�v��E���or���X� ��̑��/�Nx`)�Ȼ��F�U����t�}���W      ܵ<u��V�t̤��H3{��B��~s�k_��;  N�� ����z*�'�����Ij��z)�&�u�}�s��O��     �{ʓI;����;`&���hv�5O<�^� �4�"��pz���x���=Z�����;���ǀ     ���4u�ys�t̪�j�N�n<���V: �4�́���h����3N�hT5��ݔR�~���zm��     ��4U����r.]3ɸ}F����Y� ��d�0:����|��ú;)�&���ޗ�ԩ�����+      �%G�fcc5M&�S`6UUĜ>r�7���_�f� ��d�0�R��^(�q�[��q;"ru�\�{��N�tJW     0rD�ki<�΅��R�.]�]ʏ?��J7  �6w�����"����Y��ߎ񸎈\?�H������.]     @A9�ț����x����ii�Jp�G�j� ��f�0�Z�h�c�+�L����dR��\?�x����;�I      )GD��YMGG�p�r��tw-w:�����7�;  N�y 3���FZYY��(��n7rN)"�W�Խ�~��g      �&����C�!������P��gߓOn��^;.� p�,fX����	E4;;����{�ڵ���O��x     X)"7��+�����WJ��-{�L{�J7  �w�պv-�G]�Uw����)"�����_��F�      s.G���`%��-0�R�q�,��Xz����t �Y0p�Q��_.�PT�[#��u3��`���B�l      �%�1.��τ�4�V8<l�4�>�����[�*� p�fPu�R��{_��RΑ�7G�_lu?�q�u      ̣��~lmuJg�L�*���<��7K7  �w��y啈[���4)�������~�ݹ~��     `�4�ǽ����R�.]�}j~���n  8+� 3&-/G��,�1]&����{��D�����      ́<u��F�t̼�s�fU>~t�_���  g��`�t�_��k����d���^/���R�'��~�y#w     ��'�vll�Kw��k�n��Lj�|�OJ7  �%w����h�c�3��x�&{{�H��U����t���sF�      ��iZq��rd�\x U99Cm�=���.�  p��fH�������.�h���^���{��5#w     ����nn�X1n��R����Y���|�G~�*� p��fEJ�y���a4���A7Rjr]���~�ݾz��<     �Y�4U�ys5�Ãk�J���˗o��^;.� p��� fD�����CNo�[GGu>8���{��\���S~�     L��4us��Zj��)0�Z��5�ٗ�|��n  8k�~ 3���+�f��Q�|�$�h�R�_贞|��>     �)����7o��Ã�u99?m�۹�r寖�  8kF~ 3�~��/_v��~|�$��G��c���     0Mr����q;���"*�D�A��[O���m��  8k�ff@��/�0۾?rO)5�餥/~�S?����      ����ɤt	̾�"�Z�+8!����*�  P�q���Ν���ϗΘ}GGusxxk���W_��/:     �����͛�1{n(ED�u�NJUE��c�Q� ���\祗"RrC�$�>r��S�K_�֗.�Y     PB�Tycc5&���4�Vd���F�����Ϳ�ǥ;  J0��b�ۍ�G>R:c��6rO�~����t��     ����Nn��QU��s%?��7J7  �b�0��/���q��i�~���     �B�Ta�''��u]���S�������  ��L������+���G�_�R��     ��}���l�'&�Z�8i�>����)� P��;��j������;M�a�;F�      g���v'���1n�O����� �B3p�R��^*���pؚ�Nr     8])on��I�����I)ң����  %�L��駣z�qw"�H:<��p�$w     �ӑ�����<��RU�+��y�}t����v� ��\�L���/�NX8��e�     p�rӤ��͵d�''��u]��S2~��+�  P��;���~8�g�-���~0r#w     ������Z�=o���R�V�t�$��K��j� ����L����n��[����I�?�3���y�}      ܋���͛��p�>ߚ��{�+_��Jw  �f�0E��R��GKg0��������Rj]��.     ��j�*ol��q;���jE$��ڕ+�S: `�L���>�j�#1�����N     ��i�f}}͸NXU�ϻ���C���  ���`Z�Z���GKWp��������     ܅������4��.���R��K��]���Ͼ��?/� 0��D�G4���O�Ѩ2r     xw�iZ͍��x�'*�ȭV�
�@~�Z� `Z�L�����K�+�#w     �;�LZq��Jʹt	�'�/�T�9]����;  ���;�h=�LT/:�}��F�dw�o�     ���d��7o��q;��V+"y��&�/o_����t ��0p���_.��]H�qjvw��-     ��ɤ7n,��)�������|��n  �&� �U�<��O���n��)�����     ,��n�X*��(WU�ʤgQ�N'��z��/� 0M\����#"|�~�L&���     ,�<u�͛��pR����������}��~�t �41p((��F�G~�t�c2Iyw��k7    �E�s�||܋��~��K)En�JWp�&�/�R� �ic�PP祗"����j2Iy0�EJ�     �\������-0����N^Y�\�����  �������F��Kg����="�[�v     �M���R��4n���jE$g�-����uz�q� �ic�PH��"�]w(�AӤfg��sNF�     ������J�����Uב��ӓO�ץ  ���;@	U��^*]�	J9G���妩��    �y�#���[M;;��-0��*re��������W�t �4r�P@���"�?�+�s(�f<���     �a9"���j��m�n���R�.]A!��O�t ��2p(���+�8M{{�||�N)5�S      �U�H����-oᴤ���#��b���?[: `Z�R8c���Q=������A+���;�9�B     0�&��͵4y��ȸ}�5O<1x�+_�g�;  ����sz��ȇ��|x�u�;     0�������pʌ�IW����  ����U��G���/����a=����     �,7M+߼���q;���jE$�Y�t���O�{�;  ���;���rDr�bѤѨ����#"�n     x�<���ƍ�h���)׵q;�\��g���o��  �f� g$�z����KgPH�S��u�;     0U�hԍ7�#;�NS����L��橧���  �Ε3�i����/��$5����    ��rΑ��{���/�s/���.]�h.\8~�׾�s�;  ���;�Y�JG"n��wv�NA     
�y8\���^��{)En�JW0-����/�  0����7�ǿ�;V�D�9���^n����     �����W��v�t,�v�TU1y����t �,0p8CG����7�a�L��������
#w     ����`-�v�X���._�����~�wKw  �w�3v�[����}�f"""�<�RJM�     `~5���\����t,�V+"��L��k�\� `V����c����?�#wn��o��F�     �)�)����ё� ���jE6n�v++����ϖ�  �>���s��?�����;�[y�g�     �������w.�Fֶp�������3�����kǥ;  f��;@)M���1�ַ�ܹ���ʻ��d�     <��s�ɤ�o�XM�Gp&�*re��ۤ͓O���  ��U5@I�I�������ȝ[������	     �䈈Ѩ7n,G���DUE���L���'׾��,� 0K܁{Rյ�N�F����.r�d����~���     �9"��`)66z�[`a�d��姟���  f��;pO�Ng^�v��h���F��3)��;;�f<���     �Ky0X���N�X)En�JW0�r�ߴy��-� 0k�T�{��:��O^>:���=��~ט�?����GG픒�'      w�#R��\K�����3d�λi�y��{�~�t ���P�K�눔Jg̝|t���F���a�9<��     �$�\�͛kqtd gȸ�w�#b����t �,���o��2r?F�n��zF�     �[4M��qc-�c��,y^�{y≽g����W: `����t��F�����ǭ/�     .�F����D�|8K�Պ�99�a�쳿Z� `V��k�NǛ#��o���s�qʃA/r�d�     �*7�a?����C`�ԵC�xOyee��/�;�;  f��;p"��OG>:����w��y��I��N�i���     NnV��V�t,���\���ޚg��fz���  ��U7p2R�0r?Nr睤�������:�佣     � rD�����.����۹;U��'���  �̕7pb�����á�;�(��u��î�;     ̷�i���~.��-�p�*r�w�y���+���{�;  f��;p�rJ>؟�<����J47n��V�a������    `NM&�t��Z�R�X8��ܫk׾\: `��'.W���)��Nr7r��F����ӭ7�     �/7�ǽ|��J4ι�3��q;���p���/��^� `���"WUD��bNC>8���}-��~׈���LR���o��2r    �ٖ#���_I��-��R��j��`�4�<�ۥ  ��)pjr]���<�:��;�1b�-RD�`�ͣQ+��(     �Qykk-�����۹�N>�x��*� 0,O�Se�~z��Q|��1������!y���F�     0cr���7ϥ��C6(!��v����g���_��o��  �>�.���� ��|t�_�zL��O���!y8�'{{}#w     ��I��qc-���A!��
_�g)Eu��X: `^�g"�ZF�$���ZL����gᇤ�(5�A?�)܋    �)����^�qc%5έ�R��۹O�˗w�������  ����1r?=y4��_���[����$坝^n���  ��g�^c-��3�?��־�SW0U`(�
0�.P��f���T<�(��vҶb;،4���H��hZ�h$^��h�%;�Q:qbn����)�!]��6q����c���U眪s�9g��Z�߼8U6v����ߗ�G*��T��bW�����g   ��%y������ ���}6�O���/��   0N(�(�Q��}�����3����˕��̌�        ���`���I�˥�Y�I�=6·o�����C�:v  �qB���q8�~�B�GU���Qr�k�2o�*��       ��=�ɓ������ȳL��5�Cx׻�c�   �e �<Mc�_�K��?O�oȻݴXY�Qr       `�\���䳳���j��g�y�J�+�]���9   �w q�����#���u���J�xC����j�d���       ��so��|nnZ��<��X�k^����h.v  �qC�@<���W������_�+��xc!������g��       ��|ii�����9�I�i�r;�_��/���  `Qp%����_���O=E�o��,�v�"J�        ���0?�Y�V;
0��TJ������/_�rf�b�   G��@|f%�u�{�u�qI���:��WVj,�       �v\��y9��m�<g.�-I�۱F®]�6v  �qſ����zG����%w��<��^��L|N        8_�������9v�Ky�K�F.��y��~�   ㊂;���frJ����o��I!p��7d���rŻ�k�        ��,,.n�z�; Qnǚ+�����   �w Å%�u����W��_����;�\���F�J�       ��B���M��p��Xc�ys������9   �� ��Sr_w�K/����R�G�o��O��rM���g       �����W|vv���b� ��X�u����qG;  �8��`(������*^yE��w:����B�^�Qr       �My��A'N�b� p
�v��j5�W_���1   �w ��L��a]ǎ�}���f��2ޔI���w�%3��        0L\2_Xؤ��R�, N�܎u���������/��  0�(�j�$���Y17��̌|a��;�Z���F�J�       �UB���M�v�{��v��2�/��3�s   L�=J��/��j:�0;K�o��O��rM�L��       �T�^U��T;�S(�c�k�y�ꙙ�b�   ���� b�y������x�UJ�xkEa^�WC����       &QXY٨�'��s x��D�s翌  `RPp0:Xr_w�����ʿ�=J�x{�F9�ZQr       L��p��fk4��Q ��v�3����+���s   L

� F�Sr_y������쳔�����ԗ�k��$>3       �q�!��>7���}���Pn�:sIv�5w��  0I(�9�� u�|R�������W��z��<5��       c�h46������`�Pn� �;�.��;  �$��`$Qr wu�~Z�#G\,s�x�Q�v��;       `l���'6'++Y�( ~�v�_{��  `�Pp0�(�F��Qu{L
��;�^�����$7�       ]�y^ss��߷�a �������<���  0i(�i������j��R�SX��+
�z-�y*J�       ������2�:��1@a��/��   0�(�y��#�%���Z���m�$5e�t�fb�       ���'~��f[Y�bG�(�c��t�x��ߍ�  `Qp0(�Fq�Z33�J�83�N��k��Xs       /�</���&�z;�7@�f�w%v  �IE��ؠ�>aqQ�C�����3S��Z��T��       C(4�4??%�J��1`�ys��n�\�   ���;��B�}0��T���U����8#&I�F�;���B�<        �b:yr�-/�b�&(�#�p�uawܑ��  0�(�;�$�,�c�y���W�����M�g��I}e�&ɍ5w       @$.����������܎|�Ƣt�%���  `��`<�Qr��y�Iu�z��2�\�[��k^�(�       "�fsZ��S�SC�r;"�ݻ��_�b+v  �IF���2�(�D�g����]!p
�3b�|e��NYf!v       ��!�'6��r)v o�Ӕr;�����֭��  `�Qp0��T��b� ��|G�/Y��(���u:�//�\���       X?z����nR���0�<M��:"ٽ�?^<3ӌ �n��    IDAT `��D `칙K�����Z< o�(*����^��n�d��       �AX^�h'OVc� ��(�#���m�   �L
39%��(�SkfF��IJ�8;�v�*%w       �ZpI^���m�f��"`�QnGd�u���Ew޹;   (��$��&,.�53��G?�䎳��'E�>�L�w        ��VkJssT;����r���k��^{�?��   �x: 0Y(��w:j=���瞣���b����w:e��       8K!�D'On���r�, ޞg�vDW���̎�~!v   ��	��1�(�FQ�����9�b�g��I}y�&ɍ�       ���z����w���,[��"�Z-,����  �L$7�J%K�w��:�KyNIg�(���Z��3c�       �&\RX^ި�'kr�#��@�C�����ff�b�   ��Pp0�\,R���z�y�ũ2�^�Y
�F��;       ��\���i~~�5����e��d@d>5��k?;   ~w ��������̌�ɓ��q�����ק�i��       0��;��fg7(Ϲ�F��*��=���_�   ?��; �C�A
��j�̨x�
�8k�._^�x�Sf�       &����f[\����q/�a�7�m�Xo  B��S�;�zH���Srǹ�tҰ�R3ɍ5w       �$�</���7���f��b�={��;�\��   �� �:�eR�_���j?��zO?��s����Z��3��      `2���>??e��02(�c��M���Xo  R�8�x�Rrwu�~Z�G��h��f�T���Ě;       �+�</���-�lf�� 8�����	��=fw�ы�   o�' �O�բ;"���Ժ�^��2�d�c�       ƕ�Vk���-p����R�ys����+v   �9
� �f�D��>0�ܜ��ޫp�%w���f������      `t�$/������R)v g)I(�cx�����   Í�; ���e���P��!��?O1��O�z}��<e�       F�{�5����s��YJޖ��.��w�7|.v   �5
� �v�$J�j?���O=�b�����F9�ZJ�       0\����'���R9v g�Ӕr;�Zػ�O�;��9   ��(��p3���]�g�Q��a)�)���u�iXZ�)_�       �a��n����&��YmFQ�J	5/���?����  ��Ǔ �)J�����W��L1�.��劷�e��      `���$��<����J�< ΍g��r;�\�{����   g�� 8fR���3���S��{������ay����>O       �{�W�c�6����UY��)��_q���?��;   �� p�\���7j����~�R2�OQ�/-U��)�5w       �&�����f[X�����y�ɹ7Ős3����wc�   ���� 爒�`y������{䈟~_)p�:��Ys      ��󼬹�M�v��F���~��?�u��}�s   ��q`  ���LJ��t�zG����/K�.�d���k��n�5w       XA2��7i~~�زF�v��4�p�U�;   ��L 8O����,��P����9���k���k�ƚ;       �������7��Nc�pN�ہ���\93�W�s   �����5�i*���RX\TkfF���O!�5w       X!�$,.nf�IB���\�ގ�<v   �=
� �F����^O�GQ���\,oc��5w��g
       ΙK�ݪ��m�N�{i`�%���0B��{�^=3�\�   8{$ �Z:�J>��c�����3j�+R�K!�(L���t�ƚ;       �w��-,l����XmF��)�v���d��_�   熂; �53��.�%5�W��INʱ6:�4,-�Ě;       �)W�[���7���.�eR�g�������/��  �s�S �3�TZ�N�TkfF��/SF���|y���vY��      �rI
!	'On��b%v k$˸��H
\н|��O��  �sG� ։�Ԣ�>坎Z_��zO?�buk��M}i��y�Ew       x=W�]���M��q)�3y�ɹ�Ĉ*n����;��c�   ���� ���E��O?���K�.%w��L�F94�U3�(       L6��p���묶��v��bǎ��=��c�   ���q	 �iJ�=���ռ���y��X;�^��)��T��      �LZ����h�>-X`\$��r{��9r3�����9   p�h[��x�Ji;��	j��(���v��F���$g�      ��p/������R)v k(IV�3��W_���C�   珂; �'��+�0P��}��:O<�
�"2�N���z����Xs      0Ƃ�bee���6(�Ym�I�Rn��+��ع�7c�   �ڠ� �frJ�Q��}V��7��ܱfL���R��Rk�       Ə{��5;�%i4�� ƌg��H0��޽��<t��9   �6xJ�̤Ri�gT��j�}���^���5eyn^�׼�-�5w       #���y��I��S8��N�q_���6�۷�j�   X;� ��"�F��++j:��3�Prǚ�v;󥥚B0��      `�����t��f��i�< �ة7N;������33s�c   `�Pp��<�$^�7x!���S�|��<�莵���r%4�U3���       v��H�ĉ-��X�s�	��S�vF�0.¶m��<��9   ��hT��4�������wԼ�n�'8������bqq����5w       ��%�Fc���m�~��+0��d���3ٍ7�^�   X{�`Xp�M8qB�����.%w�9���f)���N��9      04L
��%���b++��y ��$apc'\}�Ov�w���  ��G� ���Wb��U��G�y�	W�����|i��NY��      ��WX���E���8��o��8*��ع�7b�   ���� ��L*�V����}V�{���ܱ>:�ԗ�j��Qt      �K�N��c�6[�˝10�<��	�1~�{����=;   �O1 0�\��M���(�W󮻔���ܱ>B05��hT%����      ���^���o��b5v ��L�c*lܘo޽�Wb�   ���� C̳LbQ!
�v�~�u�q�@���O�^�y���5w       ��%�������`yN�gf����1�n����_�B=v   �Z� 0�<M�4�c2��w��Z< o4(�c�x�Y����%��      �!3��?���,v �,IVG��1.�l���l�   X_�`x���BQ����w�x�e��X?Ea��T�N�,�`�      �WI8qb���O�s��;O���,`\%��ݻ'v   �?
� 0"�ԫū��VK�/Y���k�c��N'��T��Lf!v       ��%�fs���nR�ǝ00<ˤ�?�o���/�:t��9   ��x��Qb���N�=����7պ�~y�A���ܥF����5���B       �^�^E��[ly�;�`$�k���^����  ���� #��Cl�+��y�*~�J�X_Ea��T�f�̂��        o�B�'On��'k
lf �r;&H���;��~;   �v$ �(OS)McǘX�j�����{�+J�X_�^R,.N�^�$� �#      @�ճB����ݨ^��_`R$�j�� �}{��Ç#v    0�<I$��qW��Q�ff��:�c�+��V+�����̘`      &[�^���j++��a P���a��L�={~/v   w qΫ�+�S󮻔���ܱ���|y��ͪ̂I|�      ���BN��j5㍏�dɲ�,`B�~���z��?��   ��S ���%w���nW�GU���]y�m�_�����T�vKb�      {~�GXY٨�ٍ��|L3�T�3z�IR���kׯƎ  ���b  �OS�$�����{N��j��']�	#�_��y��jj�o�R.w��      ���:�)��Uہ	tz�
�0�o��λ�~!v   ( 3������m�"��La~^����=�-#S�Q�F���9      q&/����jq�*����I��H��[;������  �8(���׭8L}��*�rK�D��{=�\�Ç]�.7�~?�z���nIf�(�      ��]����Yss-�yc(0�<�Vǭ�I�$�o���1   w Wf�RIJUn��j���T��j��_xA�;�T��S4��ۙ/-�B��2��       8s.yh��u��fu:4[�	�Y&�m�d*������{O�   ���; ��4�̔��cS����͛c'�8aiI���W���\!Pt�`�`j4ʾ�\Sf�     ��f<�K>;�Ֆ�ʱ� ��L*�(�cb�ƍE����`�   ���; L 7�̔l�nS����+��i��3Ϩu�}��EJ���0_^��F�*�O�       0$L
^Y��ߪ��ilU +I�Y�A>&��tӟn��?<;   �� �ͤ$�U�V��'T��ؑ&R񓟨y��ʟ��IV��x�^�N�,�`�     ���%+7knn����5�,M�i;�_q���_���;   �� �%y�HfV��V�}�#�R)v���ݮڏ=���în��1��IC�>��LfLA      v�P�C��Aǎm�N�F+0�<�V���	�Y��={~+v   �,v  ��y��ܕ��mS^��GQ��cǚ8�^Pq옪����]�2�ܥf��Nf��=�i!wN�     ����L�z�j��	0����@����ˮ{����9   0(2��r3�L���6���*۹3v����Ժ�~��~���f`���|y�VVjr���      ���E����V-.Rn %	�v��p��������9   0<(��s��5�j�j��_�|�-�1$>p!����j=��|i�[����R5�Z3�ӷ$      8O�!XXXآ���s�ȳL���c ��La����_�b+v   
�  y�HfV��V�}�#�r9v��T��wީ���R.F�nZ,.N�n��$��      �;���Fc�fg7[�˽, �lu���)৊����>���s   `�p� ��Ӓ��뮳��nSrᅱ#M$�v�y�	���U�N�r1�$��μ^�y��2�u�      �qw�Y�v{ʏ�j++�ؙ 	���?�7�={~9v   
� ��r3�LɅ��m�)��ؑ&V����'���i#�������$If!r"      `���*~����+G 8��t�����o������   Ç�; ����{�l��\�[oeI"o6�~�au���s�8��|i��F�$��       ��/�,��o�����" �N�I	���v��z��;   �OQ �7�I"�Y��[�����*�ؑ&V�����җT����O���z���vY�      Ir!�'�hnn��9k1 ~�L^*��A��+�=\}�Gc�   ��� xSn&7S��w���+��ؑ&V��պ�~u�z��b���^�׼�)�,Ew      L�{⋋�4;�Q�w� ~^�ȳ,v
`h�n���w:�L�   ^�  ޚ�<Id�7�ԧ?���M��{��ffN��T��:�4,.N�n�D�      �%yh46����餱Bi*O��x3~�%�]�=���9   0�(� Έ'���V9x�j���\�ibǎ�u�����ߺ(#"��v;󥥚���%I;      ��N�zh6��ر���R��	�p�,[�S�Ʋ����>;   �OV �3�I"�)۳Ǧn�M�EŎ4���W�?���O��H�q�`�l���Ҕ�<�Y��     �hswɬ�N��Ǐo��e�_ �13�TZ�������ϗ�}���9   0�(� Ί�II���m��[�ݻcG�hŏ��w��(k(�������nfbG      ΉY��(�����b�t �f�du�=v`�����+���[c�   �h�� 8k�SkU?������J��5���9rD��//s~����|y�R����]�     02�
��,��]���i��3�7�e�4��z��n���;��cg  �h�� 8g�$����{m�ӟV�eK�H-�e5��%��}��;���ii�Z��VK�|6     0�B!�'�j~~��9�v o�L*�V�|�m�����W�{�}�s   `tPp �7�̔l�nӷ߮��kcG�h����j?����
eb�n7���)�t��     0d��`����fg7�����[�4�g��
^ؽ�}�{�   -�  Λ������V���T=xP�u�Q���j�韲����a��^�Y0��      ��]RXY٨����t8����LJ�Y g,I�8��wtbG  �h�� �f<I$3+8`S���lÆؑ&�O�ܿ��F�"1��IR����ũ��Rt     ���.�oбc[��(�`�I��ꛍ��|߾�/��;   Fw ��r3�L�6}���v�i��/���w*���(ch�$��?-�[��     ��V���v g'I�Y�6p�|˖��{9v   �&
� �5�f�$�MMY��P��[W�-��Zj?��?쾲�,���{��8]Pt     ��sI�++��1�2y�Ǝ��$�����c��P�   �)�  0�<Id�V����\��}M�lƎ5��_T�WT����?�:��0�բ{��Y��[��3w�Sx      �,���i[^.�`ĘIu
�\���=�}��A�   ],� ֕�IfJ��¦o�]�Ν�#M<�v�y�	���e��e��1TN�C�>���Ew      �%���ִ;��r;���$���s #ʷn�m޻��c�   �h�� Xwn���>=m�O|BՃ%^�]�����/����1���K�f��;      ΐ�Y���;�5YZ*�9Np��L�p�D����_�B=v   �6
� ���$�̬t��M��J�l�i�y��Α#j:$_X��'S�Y
KK�     �F\?+�_`�z�b;��f&�J�o&p��n������c�   ��� (7�̔\r�M�~�J�];$����]w���3.��C�(~Vt���Ҕ�;     �ds��ݮ�S�v�h�9�4�g��y�/얯��c�   �x�� 87��D*���яZ��]V.ǎ5��W���Ժ�>�'8��p*
S�Q���EB�     `�����Ǐ_h�z�b;�s�e�wV ΋���o��|��؊�   �'5 @.ɓD2S�w�M�v��m�bǂ���Լ�n��1܊�|e������g�$�     ƛ�,�v�N�B�L F���TZep�����ͮ����9   0>(� �r3y�(��B���6��8L�/��}�)5�K�'?�4��U�f����B���,Pt     +�R�N�������Qlp>�T�e�S c#l�־�[���9   0^(� ��'���V9x�j���V�	��ܜ�33�<�ף4��u���KK5�     Ƃ��C�5���/��b�x�$��a&ϲ�;) k�Tr�|��;��Q   0^�Z2 `hx�H����.���bo?���W_���?���^R�C��]�bb�+S�Y*Z�RR���Z�)��%>�   ���� �ug���i[Y)��^_kg� �9Iy��N���K����w�}8v   �
� ��b&7�m�dS��[����Q��ߔ�"v��獆�_���k���>$��    IDAT۸�R����[�Rh�JV��V��l�2��-   p���~��)v ��J����%%��N����a�KF����,[����
;v,]��c�;   ��� %O)I�|�-6��O)ٲ%v$���������=��"	C�$������T�tJ2�s     0<�D.)YXP��?T��(9�7 ր��T����j5���;;   �w ��r3y�(y�;m�s�S��bG�)��s�Z��/_X�	C�$���|qq�;�2Ew     ���T��z�_�Zl�я�.-�N`����r;�u���=�\}�=;   �Ot ��$R�bՏ~T�UWy��'��~�T�T��wީ�����[n����N'�NgJ�ja�Z�$�;_�     �䢋T=p@�m�d�E��ѣ�cf�4e�XG��k_������9   0�(�  ��K�$��)ۻצ>�%۶Ŏ���\����Լ�.���"6FG�����Th�*2���     �u�^v��~�״�WU�-[d�����<��G>"+�cG0�du��r;�n¦My{׮���  ��ǂ; `t��͔l�fӟ�����-u��-)�Ia~^���Si����*������M�۝�J��Z�'3��      ��L�Ν��ۧҦM�<���휥ݻ�n߮�#�(�8!(�QG��$Q~�Ϳw���;
   �w ���$��Y���W�s�w\aq1v,H����=����Ty���t��$q��ѰZt�y��MM��,�=�4v,     ���$*]{��{�(�VeE!��[��/��g>��7������3�2j� ����]�g�.v   L�) #���I���Km�s�Si��ؑ�:��s�Z�)��{�<�ٰ<7-/W����,I
��     �+�T޿_�~�7��T*�V��g��+�>�QU�Rv �5OSy�qx@ؾ��������  ���W� #͓DV�X���3e;wz�'��v�X8�x�U5�[�o��> �J��ct���J�Ӵ�j5O*��BH��      ���T޷O�k�Q�.�K!����T>p@���j>,o6�6,��g&O���v �Tr8�)��^�(   �� #��d��k����.��7�����b��iE��ѣ�_zIՃ=��jN�1Z���l��V�d�jn�jO�&��     `���ͪ�ۧ�ΝJ���K�o ݱCӟ��ڇ�x�5��qI�Zn00����.���ñs   `�������{?`/����9p�*7�,���_�4���J%+�ޭd���"���o����Q���^avV٥�ʪ���\b��$�y�N�$)�R)73�y݋��$���v7�   �z2K�4�Ď �/پ]���G��y��6(Y�b��Y��Ҿ}RQ�������w0��L�$�S %\s��ˏ�9v   L� c�%)Id�Vڿ_��y�1Ǐǎ���_|Q��P������{��$�Ga�t:�w:S�\vMMn&�?˅Y��)w XgY]���G   �|�)ݹS��S��dy.�����&�*�ުd�6u�xB����	`���D�6���{oѷ�;
   &w ���Sk�Ʌ��m�y�o�F�o~�5�!����O?����W�C����(�c$Y�g��2e��Ԕ�e����&���� Xw�=O(�   ��J%���Q���Vz��#����{�ҋ.R�G�����Y&W��%���ϫ���WbG  �d��] �����k*��ʷ�bӟ���.�����S��!uܽ���y�sey�tyY�Ғ<��5!.]     ���iU��^m��'�a�efg�����\t��o�Mٵ�F�` ���@$�7��>���s   `rQp �57�'��w�Ӧo�]�86��?������=��+��YVJWV���R�O�     �����T��Vm�����UW)�s)�ر~�*�>�1U�x30��lu�@�⋛W��}�M�   �l< &�'��T�����v�������ш�㽞�O?��w��������I+�+%ͦ�j�+�jU2��e0     �O�)ݱC�={T޾]I�+�z�S�+8�d�vo>,o6c���(��y��a����w䱳   `��� �����]�l��ە]sM�Hx��I�|P�v_^f���]��(�ו4�r�~�     `X���޽���k�>��-������aӟ���K/���JS��@d.�x�{�rf�bg   xo����������c�����|�T.���zf�R�J�]g�ƍ*^}U*�ة����w�,Sz�%��c�4+
%ݮ,�W/kJ%%ժ��Q��%�� �^����?� �|�%E�Vb�  ��d�VU��M����nۦ4IF��sV�Xi�>��Qq�X�8 ����v�A������+�񍃱c    ��W� ��df*�p�eW]�'�T�⋱c�x���_��z����z�k%w�<�sY�!%�ljJS����R��U��x�6     Xf�.�L�}�T޾]I�#���S��$�ʯ���K/��O�{�؉ �OS����\�ݸ�=�T�(   �$��%�G�o�N����m�;ޡ�?��<v,�o���y�ɓJ/�TV����s�幒Ng�M;v�|��J7nTh4�V� 06Xp�5; �$�TTڷO���jW_�R�����1�\t�eW]��G?��۱� x3��åT������w�ɟ|;v   �4
� �
��C����$%�x����UX\TXX��
o �8����J!(��R)I�lc,XQ(�veE���U��z���B�s���{� 0�(���� #%ٲE��n��>��E)u����b����}

'OƎ�%�j��8������^��C�&v ���ޝ�u�w��=�9�^l$H Aw$�k��HN�I'�d��I�;q��+3U�L��j��K=USSS���Ju�����m'q�Φ$vK��ˤ�E�)S�
�$ @,�lϼ8HٔD�8w�~�P�i��S�s�{��� �V� ������!c�Нm�/M��;���wde;;����a�T&��}�2��7��m�l(�z��$ �K� P&� P����۫�GU������"�$2�v��`�6ن�gϲ< �lm*R�u���o�Ѽ�    ~���   Tg��s�n5�==n�;�Q|�d�c�6҉	�<���c�\�SO������Ԕ4=-[,���
{�*�я���Ѽ'     �44(Tq�V���L�$MO�=V�L��lG���˿���k�<v��&mk���{��Ky�   ��EX6�W6����Ww횢Ç��������QSL����H�k֨04���_����Ii�� P�� e�w �8^g�x@M�>��U��T&�[�[�+L08����&'��/lm*W��������W~��(   ���X��C�~�ɂ��v�ءtlL�իyO�O���(:rD���Y#��{��$���Lʶ��߰A��A�bQ�Ą\�=" T,w (w ���`�5>����Thh��"n��D�X4�ΝR�(�{�>X��휪*Rr��;��3�{�s    ������W�{�6��ǊO�R|ℼ+d������c����,v�}y��*��%��K
C�׮�=" Tw (w ȕmmUq�>5=��֮���1�0^[��ӧ%6�����@�K7m����߽/�9   �O��=   ��Y+���[MsO����w�<��X��+���?��i�kx�)�+�Q{�����7;+��
�����*�vM���
�C��ټ�     ��Z���*��)��C�̌T*�=UU�M���n���\��h�� ��Z9�{@%K��±���W�   �T��� lp�>lp/#cd��)L�m�ܫ@z���Ç�(���-y�j�IS�0�-�d�[��А�erׯ�MO�=" �� P&lp�%c[ZTػW�O>��u��#E�sy�VLS�)l߮���W��=P���T� p�����_3�Q   ��B�`Aܫ��"0F2FުU&رC��A*Y�*Vt��L�(o�j��	�,ǲ��2��[�Z��;��J�)��4�`��@����V���P�C���*/�dX��8|���2����9n ��<��k' *�;p�O���O����    ��;�!p�>m�U&�����'䵶ʶ�q\��ݺ��,[&Ӧ�[ݧ������@�������*�ܩ�'�T�ƍ
<O6e�I})����}}�O���(�y����v��$������=��   ��"p� �Շ�}���6�kה^���T�nfF���J���uv�47s|��9'E�Vwke׬QahHA�$��@] p�2!p��V~O�yD���j��8f[{Nlk�	�|����d�� �����lm��[�z�߳g��;t�;�   P5�,�{�!p_"s�ܷn5~W����0�{*|�t|\���r���֮��8A0I�mtCٖ�7��c[��<w (w �gs�ڛ>�95l٢ ���	߮���&عSJ%��y�T&c䂀��"�Xt�#��b�W�z"�Y   �� p� �Շ�}	#c��ʕ��k��J.^�{*|�tdD���R��[�V���5�ܲ�]��c�;�G� eB� w�Z�׫������*��ɋ"�(���{:�����M���7 ��KyPU�Q��ÿ����?�=
   �P�� �Շ�=�����ׯ7��@�X[�"W�$Qr��wߕmi���$��ǲ��Y�l�������r�Ӽ~�	� P&� � v�
��S��>��u��ރMW<��a���=+73��8@����v��U'޵������?�{   �n�X��C��c$cd�-3�ݻe�@���ld�p�TR��{JN��mo�]��cuä�Lfڭ�����l-P���L��3� Pa�5<���x@Ak��7��V��l
;v(�rE�իy������{
 w!��������o��=�
  ��D�`Aܫ�{β���==&ؼY���r��yO���&'=�txX���2��C�+&IdK%�0�ii��a���v�kk�C����2� P&� ����5<���T��U`��ګ��`pP��A�ٳ,0A�`k;Pݖ-KJ��߿��~�Rޣ    w�����W�
0�ͽ���vɶ�d�ܹ�U���qEG��MN����XB�qN&����i*��C�ࠊ[��46*���ü���D� eB� c��TT�O�q�.�����	�k�񺻍�۫��))��X<�da;[ہ�e<υ�>�;��g�   �� �����Wcd$�uu�`hH����+W�
��9��.):|X�T���-y��IS�0�-��bQ^o�
�v��꒒D�k\�P���L�@2F~O��=���W��%?�eJ%�4�{:,"��j��A%~�S:Q���Ԅ����j�3���y�   �+w B�^}�+�12��
&ض��]]�ϟ�؀\��D�𰢣Ge
y]]��L?�Э[ݓDv�J�[���}�lS��Ԕ��L�S���@���cv�
��Q�SO��u���ٙ�l[;�)M04$��(�x1�q��`k;P3�m�����?��   @9�y  @�qR��y7���^7����a�qpSS���w<���;�f"w�-EY�n��bQ�]�TسG�Ȉ�'�<)7;���     �S,*ذA�֭�;;eK%�RI*��y���g�]�f��m9nr@5�<9�v�&���3M7������(   @Y������������#���߸������m�|\�̌��P�ȶ�ɶ�r����8ζ�G�̲e�ׯWq�.�k�HI���5n��6�@���@=0F~O���߯�'�P��W�1ٶ�8�{:T��i�-[��;'7=��8��X�mm�!�@Mp��i���?��k_� �Y   �r!p� �Շ��
���n�/7�]�d�Ur�!h�pׯ+:vL����V��ij�xC]3i*�مIf�J�7��}�lK���},9w (w 5�koWÞ=j|�)�mS��,of&����t�����oWz�ҫW��l�H���v��8k�>����7���,   @9�X��C�^E����x}}&ظQ�Ȉ��d�S��W�*z�m��Qy]]2w�{&IdK%�RI�}y��*l߮������J''��0�1�w (w 5��*l٢�GU�}�)X�Bލ��&��G�!�7��lC��3gX\����v�&%���0��/�   (7w B�^}ܫ�12�ȴ��`�.y+V(��(��p���Q��K33�e|��pN&�egg��w�����T��ٙ���	)Ms@�"p�2!pP<O��jx�!5>��
k��7&{Y�=��񺻍�v��S�8���bL����9�M�?����    ���   ��4���l��J/����!��T�8V��(:rD�޽���CR�H�(��n����)� ��鑿n�\)>}Z�ɓ�Ν#v    ���ѡ`�V�6��~v��ky�����/|����_(�p!�q 6�5̵�ϚةW_�{   `Q������������#���_��7*�tI�����J%�Ê��$yk�H�r<7�4��,*0F��C��-*n�.��*�JJy�Plp�2a�;�*c[ZTرC�O=��ݻUhm�W*ɖJ2�X�Eb�E��9nȅ���@sMM�;p�s}��?���,   �b!p� �Շ��##��l�]�d��?	�VՈc%g�(:vL�P��z�d�� ���q��L�[�F��A6l�mhP:5%W*�=&�*E� eB��
�BA�T<p@�(������q��x��`�x+W*9s�s�X:�da��yO`�X����u�׿���G   �;�!p�>�5�c���m��!��i�##yO��C�￯��	��f��vI��na����,<�"��fy��*)��	�Q� p�2!pP����ե�}���T���y���2Q$9����S�����6)9wNnz:�qP�<O����Ը���fݟ���   Xl� �����ט��M�`�͛��۫��%.�T73���	%�/��*�r%�(p&Me�0���T��U����CC�;:$InbB�� >�; �	�;�
㵵��g��zJ��
ZZ���dO�"*�ij2��ە^����ռ�A-�6��N�Լx۶3�{����    ��;�!p�>�5�F�n[[Ma�n��F%��<�ʸ������s�dW��mm�X>�I�R)��%��v�6�04$��MJS���l�p[� P&� *�ilTqpP�?��}��X!/eJ%΍�R��	e<O���@y#����yO`)tuM�{���w�Ey�   ,?�  ��s�J֚`�~�7���S��y��JΝ��7�!���{L^_�;�I�ˢ�R)�NU,�nܨ`˖��g�(:uJѹslv   �a�E�7mR�f�l����Jy�,�)<����k��_����T��Y+���˖%�}����Hg   ���X6�W6��	cdL08h��.%.ȕJyO�r��S:<,��]���c�4���q������vu)ؼY�;�\)9�tb��h@�c�; �	�,%�S00��}����T��U�����L�=p�lk�	�|����d���#[ہz.}���i�����=
   ���,�{�!p�#�H�Ȯ\i
{��X�����*���+:|8�;:݁;`���"��ٟ�ݷn�]�L
C�lG��; �	�;��f���x@MO<��u*44܌�9υa�E��)%�����A50F��%����%�<���?���#�Q   ���;` B�^}��1�����3�m۔^��t|<�p��qEG��]�"��!��ı܁���Q$S,���Va�66o�mn�+��y�+P/��L�,k�]����j���R�ƍ
�J2QDԎ�e����b��ӧ�4�{"T*k���pz�7�=��}���   ��;�!p�>�u�cdM�c��+�m�Q�Gu}    IDAT�d��訢Ç��Ʋ���2iz3v�c��F��^UܲE��I.�݁G� eB��\�6��ۧ�'�PÖ-
���vC�:b;;��a���g�fg���)��{ 9H׭����7�=   �?�  ��p�\�n�;Բe��xC��_��8��Pi��w?�`h�~X����X �2ׯ�Jr����f��Sq�^�k��:���)%##l   �23A ��O��
��e$�RI���]��4��o��g�U|�d�� o�H�'��v�~uv�Lm՛o�=	   �6�X6�W6�CR�{����La�6��)���yO����˗��6݁{`�D�T���ɶ�76���Qa�6�l��|��J���@�� ʄ� �44��~������'T\�^Ac����0dS;p+�7��lC��3g���N9ϓ</���%�Ԕ�~������(�Y   �<�� �:��B��6����+8s��~��J?�(��p7�$����*ر�zHf�
�z w���LJ�6���I�]�TعSnbBѩS�N�R|�2�   �3�e��[�`�y]]�I"S*�LN�=PL��l{���������{,k��@}�}>���n��?x%�Q   ���.��������?�F�n[[Ma�n��F%.H	KM���F��ޒg�;p�L�Ȇ�����kת�m�����+VHi���ubw���� ʄ� >��ޮ�m*>��zHAw�|ߗ75��T�y'`A�&ضM�����y���d���K��=	������o���?�Wy�   Tw B�^}�񉌑�5ޚ5&سG�c%�.lV+甎�d���lG�LS�>pL�Ȅ���l�y�(o�6oVî]�W���V��$7	�� ʄ��c�ut��}��xB��)��/�NO�����&��Pɇ�=��<��s� �^�g�[�>�sy�   T
?�  @���2������)r��=�dx8�p��St™�H��m���ò�Vq��G&�d�H��|_�X��n������JΟWt���3g�J���   ��3�/��G��u�֭�mhȶ��J2ccy��$7;�О������,n����?���ߟ�   @%!p  r�H��vu��_�u�8����+���{4ܭ4U����q�+8 �z5�;P&�e�Xvjj>v76�߰A�q���eE�N)���SSy�    w���{z�(X�^&nF�33y��,75���@ѡCr7n�G0&������k�i���z㍼G   *
�;  �猑1��[��߸х�����Kq��h�[�)>yR���+غ5������L�bwMMI���X���-o�Z5<򈒑�g�(:{V��h��   �g�--
֭��n���ket�V��2ׯ�=P����+����c���^c����	���q�o�ý_��d޳    ���  |��$ke��P�}�+����'���9E?���'���=$������DvzZ���6�
�:;�uu���r׮)V|���s�4�{b    �$ymm�����[�F&M�M퓓2D���scc������|A�q�'Y�� *�+����_�ڱ�g   *�;  �-g�d�L[�i����=�f���~�Qޣ�^�mt?yR^O�+>����	݁2���>=-Y+W((miQa��o��P��ΞUt����L�#   �#���uu)��a�lK�ǲa(s��-�Dґ������9�j�����=�Je��c��?������(   @�"p  �j.t���M�o���R饗�J��G�=J��5��3���D��[����ʛ�����Ţ����[��GUr��|잎��=1   �d������'S(d7熡�ؘ�\�#u#�|م�����8�j�1��v�iV �,����Y��o��y�   T2w  pG��2�	��?8�^Rx���j�|�z�
?��-[$Bw`q8'���0���/W,��v�|Pɕ+�ΞU|��˗y�   p׼�v���׭��ٙ�dʖJ2SS�ԡ��9����3g��F����w]����y�   T:w  pǜ�=Z����g���^Rt�Dޣ��˗5��.�ޮ�:�v�pEXL&�e�X����<�BA��M���퓛�Q<<���YE������=2   �
f|_�ڵ����['�l��$ٖ��	�$�{D�.%|�J���dx8�Q���e���3���?�{��y�   Tw  pW�������Wp��+=���˗�e���j��ge_~Y�p�Ν�����$��̌43#Y+W((-�oެ`�&5�����,v?{Vɕ+<�   �lk���>����֮����f�RIfl��@~\|���_Wr�R޳`1X��� pҮ��e=�Eo���(   @U p  w�#c�����/���	�^xA�ky��2H��5�����+*��+��-
���RHS��Yy���#��@i�(o�yk֨����NM):wN�ٳ�/\�ü�   �<O��5�Q�mk����"��Y� �J=���7����=����ۇ �)��M���@ߗ�<��,   @� p  ��I�1�1�ߺU�ƍ.<xP�k�ɕJy��2pׯ����
_yE�޽���Ls3�;�T��	Cy7"��rA �Ԥ`�v�8V|��s��?���՜�   PN��Y~���>y��2�Bvcl�LL��q�#(�\���
�������b0&��F,@CCj���k��=
   PM� @�8k�B�|P���.|�e�o�%�iޣ�\������*����ˬ\��`��8�╙�l�{� �{{����8���uE��+>^��07   ��Z��W���S00 �jU��q,�2SS�cw0P	���.��>���Z�y��o X ��.~���m�׾��y�   Tw  Pv�Z���?�9{����8��X(�8V���
��q�+>��lw7�;��dJ%�Н��
2��*�mwO%�����_������   �@��IAO���~�}}2R��D���$[ځ
���\x��Ç%���E��.9c�y�+����/�Y   �jD�  �1r�ȶ����^��3����JFF����'�<)���|P�ƍ�D��d~����������԰w�ҙ�,t�pA�ٳJyl:   �����]+��W^gg��q,�2ccli*Pz�r����qn �e�fq{�s �Z���?���3_�{   �Z� �E匑���n�i���r�*����k��e�k��g�^�:�V�Bw O���2�7oV�i���J�\Qt����\�(��9   `�x�V����>��%ߗ�4���T2�|��Jo���ܹ�g�b2F��$Nm����G�}�g�   �f�  `I�ݍ�u���]x���^��^�6$�/k�/�R��U��>��%�>W��
0��}f�c��MG����*��+E��K�+V2:��H   ����==
z{���ɴ��9'ǲ����$�s��9?��o(�ɔ���@��6\x��y�   T;w  ����R�`
>�`�n���·��q�5&��sϩ���*�����{�mn�{, sn��nuc���������+���Y�.d���<}   �,�'��k�����萬�I�lK��[ځj�.:rD�����u�� �(]�v��i�F��zޣ    U����D��ż� P��2������)عӕ��=ŧN�=���̨��+�}�u�mS���� *��vw)��{#x7
6mR�q�L�*��V|�b��=�tj*��  ��#��]~OO���-��Y��2SS2Q��� ~�E�+<xPnv6�q�Ȝ�I��=��V�*ŏ<���?�GN�   e��� ����Ԙ������yς;��_�ZZx�GesN�9%�î��JΟ�{"���ہd����U��>y9O��X+�2FrNJS���Y��ᇊ/^�ü�nˏ�)����{e���� �f[[��7�v�ؘ�ۈ��#��T���E�������I�5�([��</�Q Ԑt��8<pࡍ���   �� ��/}�m�/�5.4�=>�;�������)9s��>��ґ���B���<��vv��w��;$�U�Z�BAiHA��\�Ji�dtT���ٖ���	�Q1��L�Q�Lc����,h��]~�0�c�(��P� �F.y�}�*>s&�Y���<O܂���ң���o~��=
   PKܕ�_��F�w���r���,�t�F&�]|�J������G�=�]�>�,[����
v�ihXҹ �;���v�BA��7�i*%����l����/_��$�qQ���L�Q'L�(͚lK�ڵ2��12I"�ٖ�8�{L w+�\t������=�a;��.|��������=
   Pkܵ����;�y�\��s+�;���6���Q�^zInj*�p�>-p�c�ECC
��]�bI�P~�{�Y+㜌srQ�mw���,x��X2� P&�Q�PȂ��nyk��ko�<OJ�,f���nnr҅�):|Xnv6�q����;83	 w�Z��?��������{   ��n�=9��/������ffl޳���Q��7G�R��kr�R�ca��$p�g��͛Uؿ_^O�b�`�Y{3x����ǃ��_����e9�`b��@���F� ���%��[~O�����A{���~�Z�^���7�Tt�O��d�	�,c�<�ȟ�����ӼG   j��ܳS��_�υ�~��
C^S*�;j�IS��Y���%BȪ�������
��Q�}�e����}_.�G�;���;�dt�f�><�M(w (wT)������Y#��G~w�����q,{cK;A;PS\r��C���>�w�0&;�`��`q�������o?��   @-#xP����}�������C��Zc������p�W_Ut�hvA�n�9��Y�={��#��\�� ������c��sri��76��/�y�5w (wT	S(d�׬���-��s>h7q,C�Ԯ0t�ѣ
�zK�իyO�%�</;�  �,:����y�   �:�G es������;.UwԪ��=u��/+z�=.LW�{�����m�Tؿ_v��r�� *�1�9ke�w�^������-���d��J�@���B��F�]]Y̾f���v��d�D�ڣ��@sW���;���ꍵY� K ٴ�b�����{   �<(�S���/�x�a.UwԼ�c��n����=��D������߯`p��L@�2&��^(d?z^�&6M����%##�/]�6����T��; �	�;*�mn����uu�vv��}�x#f'h�KΜQt�����������K������/t����   ��ݙ�������[�w�#e��Sr�+����˗��X��}�mmU�w��]�d���"��s�,xwq�mw�t)��/_���w (w�Ķ����΂��n���匑!h�+�;�·�Rz�j��`�Y+y�x���Ҟ��e�?޿��_�{   �^<(;��oyg�����ו�, pG�1Y�����Uz�%�ccy�-n�>�
�oWa�^َ�E�����/���7=�4�sN�ؘ����tb"祝w (w,ϓ�ёmh�꒷f�LS��s2Ir3h��'��ҫW����cǤR������I��9����:��/�=   PO,��_�Rc���S������^�$�B�W^!t��R���߯`�6�G��ڛ�}?� ���Pra�����\��dtT�ŋr�R�Sc��@��c�bQ^G�|��wwK��}��f�(�I��G�甜=���a�?����r���놵r�.��E Ȥmma�Ou���|2�Y   �zÙ  ������
����ϟo�{�zF��z6�ŗ�=K��1--
v�Pa�>�e�r� @�n��r��}}HS�-���J>�h>xOFG���� P&�(�|�͘}���6c�$ɂ�8�	C��+����
T::���O�u�9�#l����y�����   �G� ����җ�6~��?�/6�=K�"p2sݣ�GUz���ɼG�+y��<O��-
�퓷vm�� � �� P�vPc~r����JFF�/_f�{�#p�2!p��og_�Z^W���.������e�(���GP!�+W����c�>�}�{�#lP\KKb}������C޳    ��3 ���ۛ��?bGG�y�R�܁�3i*�)���=p���z��={��
y��X�mw����Ƕ�KR:=�my�e�;�{� p�2!pǧ�Vފ����uv�����̶��i��=��(�ޛ��4U|���=��Op p�Q�� *ECC�<��������{   ��q� ��8��/�[������?i.Z��_~Y����Ǫi���1Ţ�m�Tؿ_��=�q Tc���F����nywN���|𞌌(��#)I��A� eB��[��fy7��5k淳�$�B��� n�]���w���҉�;��D�^S�TW(���'���_��W�   �w�) �d���o?f���	/�Y�	�;��L�Jq�ÇUz�5����G�I���3F��
vaC%O
 O�����cѻ�TF�K%W�(���}l�3�b��@���-YȾz��իe��d[Z��4I��}.fg;;�O��ӧ����>����A���8�w�O��?���;�Y    �Xb����_�������{�zA����R���B�EPс�-LK��;TػWf9���`m��=�<O��7��e_W$�8V26�tl�M�9"p�2!p���[�b~3��萷z���e���b�8�{ w���*>qB���JGG����{U3F�<��8[�nX���G�<��3�Kޣ    �p� ��;�����,���Wl��k� pf.tR���r��y�T�%p�g���>��g�;�q�'ݲ�}>zOS���]�*�v-��~#zOFG��8��k�; �	�{�]���)���V�$��c)��� (�tI��Ê�}W.���{�W)6��T�*=p�����~3�Q    �� �8�������_E�C���X���н|�.p��mkS�{���!��Ƽ�Pm�.��|���bw�>���݌�GG�\�R� ���@��W7k�\)��#���mo�bv�nne'fp�\����q�o��td����ܫ
�T2c�>��_���_}>�Q    |g ���?�g�6x��/�8�h�wo>tC�����^�+���*Us�>��l٢`�y==yO�����A�m{�q��'�wI����+W�\����%��J���
�@��Wk�Z�mf_�*����!���vǒ�p�ґ�s����{� lP���������y�   �'qF@�N��~����4i��(5���ws����u�o(z�-B�����v�*CC
v�b�;���������y�٭�/�0Tr�j����U�7>wlZ�D� P&��
���d�ڲ;;�����4���� �Ǌ�_���JΞ]�f�+���ۚ:��{�����/�9    �g ������7���$r_�@���F��_����{��Pk���mS�k���k�@�m�nL�ܺ�=M����o{�����!p�2!pϝij�6�wtd��;:dZ[etㆸ���Ɔv X,ɥK��Q|���/� p�PllPE������~[�s    �d�a PN��/����˿B�^~���0i*E���Q����_�{��V����lG���;���Vw ���,x�%zw�f��-ѻ$���ن��իJ����I$� P&�K�Zy+W�����.��]��%���F�n�$�ړ$��7;���w9�td$�9D�^Q�T�e˅ޗ_��{    ��3 *��_���^{�g������X\&M�$qѱc
_}U��D�#U�z��y��ѧ�    IDAT�M���!�z�ڼ'P����~��ݘ�M�\�~k�>=�dl,��>�_�"E���; �	���0Ţ��+�uvʶ�eQ{{�LHi*3��}n;;�� ,���%E�g������&p��d7]��Y? 5 ٴ�R���L�y�iw   T8�8 �(�闾Sx�v\�+w`i�4����Ǐ���J�^�{��RW��-��V��;eZZ�@r����s��o����ѻsN��D���g��ؘ��q������@������+W�[�Jv�*y���V�ʞ 5��}.f�� r⦧��#G�^���8C��3�v U*Y�������^��Ӝ#   � g T�3��/xo���!r/w`i݈]|�J/��tt4�*B��󬕿a���;�o��Vw ��5|w�/��	7�7iz��JJ''��}l�f�>>.W*��'Xw (�;�y�V��]�B^[���6�U�d�/�1&���2Irs+; T��9����'OJI��D�E���v Ṷ_�Qq;   PU8�"����38xp?�\�w�@>�B����Uz�%/�=R��>p��iiQ04�`�Nٕ+� n��nD�s�R�.I��������U�׮)W:5�ǟ��@���\Ⱦre��\y3d���F�$��(��s] *���Tt�X���ڵ���L�K�Z9k9��j��֍������   Յ3 *�������������+9sƕ^zIɅy����0F^__�o�"A���ͅ�l|w�fh?!|wQ�d||>xO�ǳ���5�(Z�?�; �I����緱��즭�fȞ�R���q��=I���JǊ�_ѱc�O����-�%bmvt�s �=�׭�'n   ����v������V^���;P�C��a��F���:B���L�(�&;v������`�͍�7>dm�1����w��TR:1�m}�>��Pr���$�2*�; �I��X�6�߈��U��˖�8���5��=Id☍� �N::��w=*7=��8w��}����������{��O��=   ����  >��#��8��q�ȑ�y� ���m���5�==J.\p��+~�}�ȕJ���wޑ]�\�ࠂݻeW��{4 �di��~Q��w����s[���wcd�56�����?��T���|�����1�8^�? ��Y+��2��ݶ�ʶ��[�J&n~}�5d�{j �'nvV�
�zK��H��R��!Ioﵦ��u��   @�b5$���~ڞ���O�ǎ��{�j�w�B9'�ґ�����ǫ�Q����`����CC
6o�|�MP����wy�܍�H�_��/����J&&�^��}���׮}f��w (�j��n�����Z[����5��W��iiɾ椩Lߌؓ��ߓ�CI���=��ԩ�z�c�{�i�= Ԋ���Z���}_��d޳    �{tF ���ַ�s��?��~�Þ�g�6�@���?��f�$yOUv�����V��!y��y� �b.x��)�����������I��o����SS�Ð� ʡ�wϻ�/_.�bE�/_.��"cL�ߺ�=�k*���I/_Vt옢wߕ���{�EA�^&7n8�Z�������t�+�y�   ���������}�}��w򞥚��ä��Ԕ��~[���r����L����
��l�.�Ғ�8 �4�6
�m~�6�2hm0ވ�o��=Me�_51��MN�t||��tz�0 ���X�]�,�[[���F�n��onb����f� u�MO+z�]Eǎ)�{�EG�~�ɢv�v 5���   @m�3PU��O۳/�x��uy�R-܁�2h(]t��Jo�!7Y��b	���������!�&�B!�  �܌߭�X?���:Z���<H�tb¥���]�����.��pnb¹��]29�j��* pW��߿�/[���˗���\���i��=I�� I���;��ԩ�|"�'!p�s�8C�F���ז=�غ�_��x޳    (�b �:���_<��w�z݈8\|��Jo��������/.S(�߼Y�������� �ʶ�;�y�</5֦�6u����l뻑s���<�qΥ��J''oF�nn���t��q������ڏ�7"���3MMٓ7n����g�����{�~眪��n����bSX$!��l�2f��xñ�`g�Or'y�ܞ之����:�Ƀs�b�%��g�	BHn!��[��$��ݵ��?NUwkC-����ޯ穧���:���|�Saxҧr  �p�>7mRa�&��^��8A��,lP�3�������   @ma5@U��}������;n߮�ڵ*����p9��Y��/V��K�M��z H4k���Yy���[šw+ϳ��"�y�'ɖ�:�:Jڨ���c���{O��Ax{�X���ciP�N�#��QިQ2�G�/7��-�hy� ������l`H�Ç�P�[o)z�}��8G�}</��+V� Ըpڴ�ŋ�/~��g   PY�j �Z����`�ƹ�gI2�@m0R0$����kUش�j!���&OV��K���b��f�� @u�<k=O��#���&�G������||9_�����zz�y� I�l֘�&y��F�G3z�W=��=Z��I^c��Jo���� p�lO���7���[
�y��8�B��Cx����� �vڴc�/�G�   �M� T5���u���֠����ipjO��]���m��7TذA�Pp=և"���)�=[���*X�@&�v= �c$߷2���x^Tn�����d�5F���O�g4ah��^EǎY��_���V��}���5�Q ���Lc�1٬1������Ƿ�@���T�(d�Y��&��Fy���d��d2�$OQdly
��vz&��7� *�PPa�67mRq׮�MC8	�3�� �b��noٲ��~���Q    rF ��mm�:V�����\ϒD܁��t�鱅u�_�V����X�D�=9L:�`�_���%: ����M��<�ʘr||����0��5���nz{m��km_��zz��k{{m��'���}}����ԊL��MM2٬Q6kLs��� {c�Q6k�lV^S�1�t 4Ɩ��xc��3�E�`�߀ERq� #%��ޭ�[o��u�l.�z��#�^b������DӦk������N׳    >�x �	����x�ŭ�ƍ4����;P��$E�T(�ʿ���#G\�u��d�Y�)�h��3�W�$�}k�Q��_��x^d���Zc�a��DQ���k���R.�����0|o�J���#�g����fM)�.����dLc��Y���7�������S
�{6�ʷ���0�h $ڿ_���Ra�&��n��T���lP��iӺ�/�������   ��b�@Ͱ��^��/o6l��}�@}1�Jah�[�*�f���d�pO>o��8�~���Lq= �L�A�R����qصt�1&ɫ?/�C�CY*���S��g��7×�﹜�������`|.gm>?�t �L:-�Ԧn�Y�55ɜ�uCCjoh�1F��z|_�Z���ˡuE�ܼ^�-�!�� P%�>Pq�f�zK�{��j�m���d=�U6 u+�1�H�d���?|��,    �+  j�mm�:^ziK��6��,IA��?F�;���ʯ]�b{{���	��ś8Q��/V�h��q�\� ���	>�z�5�P|����x^dJ���i�/3�Z��)*ߕ�٨tm���`|>](���|�@{<�����a�8���e��kl�J_��ֽ�k��e��NjXhZ76���q�QƟ�`�hZ��b��UؼY�͛������ZQww�� ����pp���?�p��Y    �VB ����u�^�!x��K\ϒ܁:g��������u*l� [(�����Z���q���E2�ͮ� ��8��R;����Ǥ�`�)�1�A�r0^�qX�,֡LY���!�BA6����@0>�����@`��,�WU���ˤR�!u�� ��`���3�54H٬J�������z�>�%��a]��d��� ��ӣ��o����
��!�^a�p��/y��1 ��h޼�3?��٦����   �'W Ԭ�[o]�����~�;�2ER.gmmʿ���#GF�gp��'�,�-R�p�LC��  	U�[cd��K!���r@�?_˗�O)oN�-�EX�P�[�K���
kˡ��>k��ds����^��+���
ih0~:-e2�d2R:m���L�(���� e2*�M�uj7��Zc��_�Zc����
��7�GQ�� �ӳ}}*nݪ���*vt�7�����YI IRq��wf�|s�im��   �:�����~��/�^}�[�'�	��H�	�(�ŭ[��u�����%�^c|_AK���.R�`aw ���/��cl�A>��wJ�gM�Քt����Sf���4(4�}���vx��'�rqS|.g߶�\��*o�m��m��xCCܞR&#�J�L9�2AS�RF��g2��:�6^&clx&�*�Y�;��)]�����4� ����Tܾ]ŷ�Vq�N)]�Tj2�N� N.Z�>���溞   ��� �y�w������zmr'��TJ��ZE��6�v�
�6[����
�̉����v $Z9��,_���j�� ��/=^~��Ue)D�r��V�ད���e��d�y�P�|^��s����V�|�-r9�(R����!�H���s���j�]����<OJ�=E���ϓR)c�LƗ$�N�A ���1ƤR�L��$y���1��{^X����oL:-�N�!v�7����5�
�[k��  $^���Ν*lڤp�N񦶑WSwϋ�� ��/�t[���/t=    w8o�.����N���g��ca	�8#ke�����_�6n)�� �^� �/\7�g2�'    ��E��ݻUظQ�m���p7�>�n����o> �$��7g��^�z    n�3P7v�u�㩕+�h�,�N��P)npC[ܼY�5k<X��M��v    T�bQ��v�oWq�Vٞ���j���m��i�W^���_�b��9    ��

������af�ʯ�b�n���c�d��ە��o�칟7$�^�L*%�\�-�?w�L:�z$     NV(��s��[���cM�	Uuwϋ�Y��3F�%������(    ��� ug��?��V����$�N��y�V�Z�Çm~�:6l�-���p
e�f�y�\x�Lc��     ��PP��Cŷ�Vq�6B�U�j�7� >�1*.[���g����Q    $9# uiח�Ԛz��?V>_��A� *�D����B[�򯽦�ȑ!�^�8%ϓ?}���.Rj�"��&�    ���S�ޮ���*n�*�ϻ	g!�wc�P;+a 04�����O�<���]�    YX]P�v~��z��?55r'��Ҍ�R��-ʯ[�pϞ3��8#c�_pAv_�Pf�(�    j����[���k�T,�	�(�w�� p֌����������{]�    yXeP�v~�k�������^��,Å�;��`$�Z�ZE��o���_���;Ζ7i�R*��by�ǻ    P�lo��;vġ��;�0t=* Qwϓ|?!� @�}^w�_�^��ף    H&rF ���{��{���u���z��@��H0Q$��i����):p��	��|�S�(��"ț8��8    ����TܶM�m���+E��Pa���H�'��lo �T����{s������(    ��� H��կ~�a���׳Tw #ɔZ�ý{ma�Z�m��;*�;V���
�ϗ?kVܔ    �k���*����۷+ܿ?��9�,g�r��U. 8w���������z    ��
 �l��ז4�Y��:�v=K%p���2��vw��ƍʯ[g�#��B�1٬�y���ܹ2�څ    N'���NjߺUkueD��ġv�` 篡!ҍ7�?������(    ���# �����e^|q���g�� \2R�Q�Qd�[�����
;:hRCřTJ~KKx_�@����H    �J*T��C�۶��r�'�##p7F�}Y���"lssX���{�>���g   PX���|��)��/o�w��z�J � )�����R��M�7��d4���ɟ>]���
.�P���'    ��ӣ�Ν*n٢�]R��z$$���=O����[@��Ə�篹����U�g   P=<�)�l����l�>��,狀;��8nCE�����7+�n��\��:�M��`�ȟ2%na    $Rt�۶��u���N>'�x���v 6��ɽ�%W�y䑷]�   ���R ����{S��n����,׳�� ���R�{�٩�ڵ*l�,��H��:b��̛�`�<�--2��    �����={Tܾ]�;���뉐p�{����Fx &ьG�/�h�~��z    Շ �����x����U���;��8�(�d�Ua��7l�=zt$�B=�3f(hiQp��Əw=    ��۫��#�o�&�˹	U���� �&\���Y7�<Ǵ��]�   �:x�!���Ϭ�x�S��K�@RyCd�E
;:�_�^�m�huǈ�ƎU0�����Ϛ%q�    *&:x0�o߮p߾��?p�)�N[; ��pѢ��/�4��    ��8 0Dw��f��&�\�rV�H���Y+Y+{�
mm*l��ǔcĘlV�����w���z$    �.���}�Tܾ]�-[��6T̐��ġv�� #���ju˿����G   P�<�Y���/������X���'w Iq^�A�UܲE�P��h���}�3g*�;W�ܹ�&Nt=    $R��7��ܩ���R��z$Ԡ3�ik���y��-�٬���Nף    ��� �Y���/�Q���D}}U�%� )*�!*��������ʯ[����J|g`ȼѣ�ϛ�`��--2��    ��(R�w��;v��c���]O�:pʀ;m� ���}����9wŊ{]�   �vx�s�q�=_�_|�ou���z�3!� )*�!*����N֯W�hu���<�ӧ+�?_~K��)Sh�   P��c*��7���%�˹	u渀;m� �V:m�o�O�~��?v=
   ���j ��-_��'�������)׳|� �bX7DQD�;�45)�3�?�n\�    �PP�o����
��vv�����l 8c���~s�O~�g   P{<�y���o_شr�:��w]�r:�$ňl�NluߴI6�������Ϙ�`�\s�ț4�F9    U!z�=w�R�k��{�HŢ둀8���R�� ��=�^�������,    j�
 8O;x`J�z�f��}��YN��;����-�,k�V�͛UX���98g�Ϛ���E��y2�F�	    $I6�W�{��۷+ܹSё#�G$I֘8�~��	��C���9-_~ìGy��,    j�G ��m�ߟImذ5ؼy��YND�@R8�juϿ���۷��8�7v���--��̑�d\�   �^X�p�~���*��+ܳG
C�S1c�v�;ݯ � ���ӻ{/^���G���   @m#� b[[��k֬�׭��䬯p�I��ׯW��g]��,̜�x�&O>��    �K��5h����u=p��P��_'g �H��rh�u�-��C]�g   P�� @�0����+�o�����WoHR� P�����E2Q$��H�bQ�]�TܵK9I��Q��Y
ZZ̝+3z��	   T�۫��#���+�"����ġ�ӷ�  ����>��E����z    ��J@ �w��xjժ߲Ţ��,� �"	�|[���{n�k��@�yc�����--2�G   �4���}���������d��P��}z��`����W����u=
   ��B�; �����R�W���q�    IDAT�!x����^�g  ���[�}�?�(JD,��R�~�
��K�'�d�3fė9sd2�#   iQ������q�}�^�H�*�˖�a�a� ���}^w�c-+V|��,    ��G 0�v�k_0+W>f��]�@�;��H���)���t�jP���g̐��   Ԣ��k оk�l.�z$��#[nk�l `�54D����9?���\�   �>%!g 5m�7�qU�WV�\�|� �"	�!��huG2���3����Y�&O>׏|   �Xt���={vt���!{�둀��8�><�G	��0�c��믿�Gy��,    ��~ 0����_���������ߵk��y  g�����}Y��6�Wq�w�PN��f�Ϛ%��8�>i�w    ��Ç�ޭp�nw���v=0d�M����M�ړ��߸f�#�lt=   ��F� F��?���k�wʄ�淃��9,�@v�"�(�ށ����*n٢�-q�=��7m����--�L!|    8uu)ܻ7��ڥ�\��c�� ��f��}o����=�P��Y    � ����o>x��G*9����f�� �K(�֦�瞫�7��5�����M���   ����ܩ���#g��r�4 @���^�u���_�z    (�� FX�3�|l�]w�Mvժ��X$	 �lp���q�{��
8+6�S�ޮ��]�d�iyӧx   * �ꊏ���U�{7�vT7ϋ���0 ���h���f?��-�G   �����z��;���M�^�/���[�#[
��Z)%kivGձ����L&�_p���3�O�*�Rn�   �(�����{�ā�={d�s=p^�1��� @mI�l���|��O~��(    p"� ������;�ws�������b{ ��)(mڣH6�d,����ds9w�Pqǎ�ϓ?yrz�1C���2٬�!   
����a�}��@{_�멀�F� j�ml�����'����Y    �T(� Ƕ�We֬Yi��o��?����f�� �K(�֦��s7@�Aw��1�ر��3�M��z$   ��lO��wމ�{�*�씊E�ca��߰���G
V �<D���|�ͳyd��Y    �th ����_����`��j����-S\� F����V�"�(r=PQW���.6n�$��f�Ӧɿ��--�L��   @���
��U��]�}��˨-���� �Bt�GK�^6��w��    >w H�y����������7�7�\l8Q ��Ԉf}��;j���Vq�6�m�$�tZ���-�\ ��:�   $�><�ξ{��#G\OT���@;�v �;т�f�|�<�ښw=    �	+W �0�>���W�����F���>����= 環!ʷ����\�qz��Q/��7aB��~��O�7a�
   ��ݭ�w�ۧ�wuv�
������P;1 p6�Qx�����/��    ��w H�9+V|q�����������<��  F��f�(���|�j���Tt�
6H�L&#oҤ���3d
  ���
�{O�޽�:;�߯��\O;k��y����� ��o�u�=9{Ŋ/�    �w H���?�����7�W��G����y  ��լ�v����FͲ��½{���a���ZާM��   C����w�UTnh?p@
C�c#�j�7Н«( �SQ����C�O~�]�    g�5- H�m��?/�r���}���=F�w������sI�������s��8?4����tZ����N�7uj|=q��   ����8���3~��=�ǎ�Q�
��8E ��	�pɒ[[{�W�g   �sA�; $؂�Ƕ����֦��mN¡  ������	��N�|���wI��Y��i�O�?}���Se2�S  `؄�����n�%:x0~#0Pg�0� �h���{/���>���,    p��J@�h�����^��lO��� )��!���S!��;V���-��ԩR���  �J):|Xag�����z�~�B��d�3����� �^z����?��9    �|q� �D�3�|���~����^���瓐 $�1���gwKawYށ:uu)��6n����'ާL�7q���n  @�ZE����}w ̞ϻ�pϘ8��� ��	k�����+V|��(    P	������'�g�׿��{��a�� �d�Nz[�݁X���w����>}_���q؝�w  �e������W�w�lo�뱀� � 8��94�]��f>��_��    *�` �B����"o��׼}����kG�w������sI�������s��p��;pfA �$yӦɟ2E�ԩ4�  ����Kс��w�%���5F���3aa J�ĉ}vٲO�z䑕�g   �J�� �P�~��>���=��ϛͦM3� $\���J�݁�)����w�hz/�ާN��ާL�?q��J��   y�PѡC
P�|��)�˹�H.cd	� �Q4o��Q�\�h�Cu��    *�L$ T��;����f�gL��q�$E6Du��~:�{I�&��	H<ϓ7z��I����ԩ�M�i:��   ���+:|X���q+{g����e�3�f����^�[@}3F��/ok��/�    �� P�f?���{����}���7�gE  gǘ�R:�n�h����E���.E]]*n���ih�7q���S���ԩ�&L��c   U���):x0�wv*ܿ_���|p� *&������<��}�G   ��D� j��'����޻*��+�ÇӮ� T��	w+ŭ�4�Cf���ݫp����L&3��>i��ɓ�M�(��  $L������+z�=����vw���J�� �fG�
��˿5��'~�z    n��F�{�៿���?���ڼ]�ƕ��"�D ��t"ޖ��Q�x(���\�л$����}�DyS���V��t  0�lwwd?xPQg���:$[(��j�� ��N�z,�U��{�6׳    �H � 5ƶ�z������ˍ��F�V��;�M��6�SI�������s�Ǩ~�JQD��4ߗ7~��	��{c�H&	[Q  Pml_����8�������q=P3l9��1�H�� ��͛�?{��N���9�z    )��@��y�]��W����E� P��\r	�} �$aD�}v��ih�7y��I�����	�&M��f]�  ��XTt����ST���'{�Pi֘8�N��%� ��x�UϷ<��'\�    #��7 �a�����^~�Auw���^�X7�,���I��pf�������k���f�M�4��^�75�  ��+:|XѡCq+��C�����cq â?����GA�E 5Ϧ�6���?k����}׳    �I� �ў{�Yf׮���ٙ��`�Le�C�f� QI��paQ4xw=PGL&#oܸ��}�e�& ���OQWWb?x0�]
��7�#[�=��(8B 5-?>�/_��^��#ϸ�    \��6 ԁ=��{�pÆ�A[�I�F�V��;�M��~ ��I����C�vwC�$���d���'L�o�'o�8)\� @]�G�(,��jf�==�Gꎕ�14���YQK���E�/|��}�g    �X��:�����"X��N�FA��M7)��R� FD66���8�N�Hϓ7fLx|�0A����t  T�B!�wu��Rt��l.�z:��3��N���pP{<O�UW����7�    ���: �3{����]�W�7s��/I�ŋ�p�M��38 �W62����nm|@��L&ny/7��[�Ǐ�R)�� �a8`���r�pb?z��t J�$c�l��Պ ���!�>��<��?�cף    @R$!g a;�����WW���,I��j�������a���*E� �44�;Vf�Xyc�����'�ɸ �aa��<��˗R#;�P$WK;��ZA�@͈&N싮��������Y     I��3 8����3�-[��ׯ�X��5J�;�7u*� �"	�U�vw�j�����}�Ō�\� �酡�#Guuɖ��V��.�Xt=!��0f ��W�"	 Ԅh޼����fѸ��r=    $�z P�������Uw�X4
e?�I�]��@�%a�B���E�@û�Y �3�������c�ķǌ�7j�� �ag{z� ���n��=J;P�hi�+�T5��6�t�?�����p=    $� ��}�+�Ȭ^��IJ/^���n�5���$lP��ke�H6��@����Q�d��e����)��i� �Q*:zt��}p����es9��c�vZ��w U�67�����|��?w=    $+~  IҾXX\��5ϞQ��Ϙ��;��W ��$lL��(k�(��V�vw���tz��}̘��}��ѣ�-���zD �H(}���#Gd��.5�����@�)�ii�wl�T�pڴnٲf����]�    IG� �o���gR�6�:hk[ k���wʛ:����	�:A�;P��@^��}p�;V^s��ƌ�R)6 �p���?�n����_�v�^�ҎSc' ��XI�e�m�u����֢�y    �� 8I��?�Cժ�+�7
eo�I����� p^��!�^���ox��@ݲ��de�LS��r���Q����Ms�dHO��)=*{�hܼ^jb�Ʈ"���Yc�vZ�qz�T�.[����~��g   �j�	[ �)����^��С�$�.�D�O}J���w 8'I�xpG�ݽ?��.�܇�44�����r�{�_�7N�d��k�D�}}ǵ���nE�ݲǎŁ��m�� ��v�=v$ ��3�PX��w�>���g   �j�J! ��~������f���$�de�Cf�X� �Z6�qke���]gp
��Ȍ-oԨ��}�(��F���MM2�FIA��]  ��\�FG�*:z���n٣Ge��[׻��F�����
 ���v�'^�H�h���ë��j�_�U��Y    �q� pF���R��v��Ec�i5|��
.d�$a�A��v7��5g8�Ce2��f����B�^S�LSS�XS�Lccv� �I�`�ѣ�zzd{z��z�v���>v,�
�$K�2�s`���v�Ҏ��E;��2F��/ok��/�    ��� �!���/�^zժ��=�KRz�b5�t�����I�Ƃ�;Ί�2Q$E����ܹ����!�l6�g�q��1����J_+�f��d����m)�����+���w CV
�[��>�P�l&��\��[�z��p=    T;V C����V��::�H�?u�����̘1�O �Q6�q^��?���TE��l�L6�ˁ�lv _�44�ߖ�'aw`�r9k{zd{{Oy�ʏ�������:w �c��vv�s=j_m��	vʔ^��+���G�z    ���  ����u������7�*�d�Yeo�U��9�S |�$l$��b��/�л�y |�����Nx?U�44H��J���y���닃�\����B�'�����=�~.�̖�쥶v`���=�d	-jO]tѥ�~���,    P+Xq �����I�Y�]����e�.U�dٷ 8�$l�c��[γIC��<�L&����4(���d��3�����$ ��C�6���x����@}�� {9��ñ=�D���-�ۖ��o��    j+� �s��w��pժ�:;��̜��g?+56�p�$l�cĔ�D���w�JAw�T�?�TJ&���oh�L�T������A�����8�0�*�6�|^*e��8x^(ķ�y�tm��8�^(�
���\|�P��pꇕd��oi����I±= ���ɽ����͹?�ѿ��    j� ��b|�iϳ���{�9�V��Q��n�?{6� �I�F��;�!�8E��6�L�л	�8���}��僠��^��!zϓ|?�?&<�y�mI&��`*%y��(��%Ɇ����?Tn4���E���_z\�|��
������ ��h������;P۬4���y��>�� ����K.ٞ���ߘ���=��   �Z�� @Et|����7��y�<e�/W��d�e_@R2<	�#��[��#��;*jP ��_
���Sih8�q���'�JCh"��\�k�W
�����F����
RynT'�@m����j�>�p¦�6��GZV��׳    @��| �b�}�_y埼����̛�쭷J�� �8�$���*5�Zg�aA� *��;P�hhG�����&N�+.]z����_]�    ��L @�\�����t�����[�1*�ءc�<���w9�  ���<��eS)� ����M    Α5F�������JI�O� ��-X�oԧ>5�p;    � �a����^}����j��F�����Pǒ���U�ځK%�T��2hp�ɘ�Ͳ��Q�8�02�i.Y��짟���(    PoX� �9O>���-�|�N�֣bQ}��o�{��|��  ��r8���T*ny�}Y�#b   Գ�k�}�v  �_4qb߱��v��    �i ����{���6n|�߰�Y+o�heo�M���L��4��fE���w ǡ� *�w��rC;ov8�0����Z���q=��z    �W�� FĎ����ի�7��y�<e�/W��ke�u#	Ov�Q$Y;z�w ���Ȳ�@��'����H�m�dɣ��   �{|N% `D�{��o�o���Ѵi=�"�V�RϓOJ==��  ��<O�}� �M��kϋ2    �*�[��?�WH�O� ������wn   �d`U 0�:��ݦ�u��6n�P��d���r���s�'5.	Or܁�r���R%��	'��2hp*Ș�����Pql�����7͟�x����Q׳     b�� �h�����Y���x2F�+�T�G?*�y움��'7w�CD������{��@�p�� ����0���L��� *�f26\�쑖+~��,    �㱊
 pf������ֽ���5N��)S���v�q��?5(	Ol��Y(���ZKv Ս�; Tw`h�4d���8o�ԩ=�W�y������,    ����
 pʶ�zo��o��_����1��27ܠԕW��jL��܁sc�8�^nw/��w ���i7�������3�y
/��m���/1��y��     N��V @"���W�I�Y����$�.Tç?-��쫀��'3w��hyG� � �A�(P�[�	��pl���ѣ���W�Q˓O>�z    ��c� ���{����-��6͖$o�eo�M���쯀��'2w`D�����ޑ ��2��Ycd��� �8�p֢��Å+��r���v=    ��X� $N�]w�(X��m.���Y�\�뮓���PŒ�&�8`��M��A]"� �A���;av �8�0t�-.Y�Ӗ���mף     ��s=   '���S_�喛�i�zEʭZ��'��zz8q @�1F�<)�TJ6��Yϓ5�T   �0&>&����4���Y}?>~%� @ճS���?���n   ���
-  ���&�}�jݺ+E2����r��9s�U(	O\܁��n����hp�ʠ���J��ׁZ��=�e�Qt�%[g�x�妵5�z    ��c �x����?�^y�߫�ۗ1J/Y���|D��؏U$	OX�@��?�n	��<p�� ��ja	���c{ ��U�.��9?���\�    8w�� �B�}�͵6���m�l$y'*{��&Of_T�$<Y	���JqȽv/�I/�    IDAT�]��@� *��;ɘ8�N��'�8����px�UW����jw=    ���� �*����W_���r��@�k�U�kd�e�$\��܁D�;���; Tw�d���� ��c{ �K�l�������3��    P��  8-+V�v�'>�);}�1�ʽ�����ǲ|�I  �Q�������T|	Yϓ5��  @�1&>����.��R))$ߧ�  �L�-�t�g	�   @ma P�lk���������
C�LF��~T��/g�$T��4�u�Z)�Z�]σC�; T���Fvk�i ΄c{ �1
/�dkj��+�?�p��q     ��:1 �����W��z�տ0��%)�p�n�Yjh`$L�����v��2�ۨ9��2��|Xi �N;��ñ=P�lccT���<����z    ��` P��~����7o�%ke�����g�ϙ�~H�$<!	��rȝ���A� *��;��0;�aƱ=P�¹s�3K�^;�����z    ��aU P3���ς5k��zz|��嗫����}�w@$�H��y��N�p�� �������r���% ���@���ղeO�\�⋮g    ?V� 5�o~�Q�����Ν�%ɛ0A��n�7y2�<��$<		��$+ɜ*�n�Z$w ��u��;� �ñ=Pg3?�-�̜'�X�z    ��` P�v�q��S���i
F������\{�,�>��$<��1��[ߝ!� �A��>�b�_@�plԋt�������gw�    0�<�  0���?����O�f�M;�(Rn�*{�	ٮ.N~  ��g��y��KA R*%��/�y�1   ���I</>F	�TJ
����8V  �ةS����o'�    ���i @M���ޞ7�x�[��*�I����ǔ��r���K�w �uB�h{�(��2hp�>V�1��Vv �n�5���-\~����^�ܴ�]�    p��l @]�}�=w��_�[��$s�*���H������'w UǖrQ����d9�w ���v�;�b j��@��&䢥K�9��Gw=    �-V� uc���gR;v��[�Ta(�Ԥ�?-�\���H���;��Rnz�V����"� �A�=��wh4��o�5�z���.k�}��KLkk��<     �X� ԝ�_��7��^��С�$�.T��7K��a��'w u�|����c��2��+�s�Fv �ı=PS���������?t=     9X ԥ��~����mU�~�劢�����ϟϾ&IxrpP��4�N� *��{��C���`�8�j�1
/��}��W^9�\�    HV� um�o�ֿ֮���H���)	O*� p����{�	�@ep?��`8plT9;zt!\��OZ~���z    @2�� �{��{�������Z�܁a��'w 8����VvP�ݖ� w ��`L��91��� '��*e%���?o�U�{��y     ��*;  %�_����~�tw�m�@�%�D� �����������; TF��K!vSnc/�-Xc�: ���@���aqɒ�w������    �|�� 0��o}kfj����ޚC�;PYIxp�v�����p�ʨـ�i�5���Z��=Pe�y��kɒ�g}��;\�    ��� p
;���S���s�(m�@�$��C� fp�|����1"� �P��rӺ\/]J� @u�����1�K��p�SO��z ��ٹ����N����$ے�y�dɒeK�m�1	�vf�vnJ�,P�܄I�i�;y��z�f�ܧ�3�tڛ���%�@I�L�i�df�4��$���"/1�"�����1a���H�����2����~�}? ������O�������{�[پ���������;�(���{��K���0�7ph���2\�v����a�ww?Ѽlٻg�y羬�   0��~ x?��_�<�ȯ�N��Dx�;�]y��1p�^��|����12���)��ꧯ_�{ �n9������Z���=�+Yg  `�r  o�?������kOs��/?,� ��i��+~�Mi��=�?q=�x��J��<J���;<n`��_���Y�  `tsJ  o��~������AOs��.?$� ����ݓ4}ipi�����'��$"R�u .r&�4�B�z��n��W�U�Y   �& �[t賟�\ڹ���lY����oR~@�
�!�$"ҋF��@������Ș�9�&I����V�Z=�_x&�<   �N �m:�я~2ٸ���O�""����|����?E~0�
��`.z*�K���t/4���5�i�D�Ҙ��_/�7._8 xM�4�@:mڹt͚ϵ�{�d�  ���a ��>��ɱm��Զo�K��H�����k��t�{,�J~(�
+���G�?���F����q�S�_c����!������Pl�1d()���˖m�\��dp�|�y   �F @�v��ˏ<�;������h���H&Nt������;@a���EO�y��^�c`��iOW�����Ju��  ����O�~vd��Oο�Yg  `ls �>�`����YiӦ�$�V��n]4�]�{.������
?���>�>)��^�����;�zOT�������5*B0�)�p�U�i}���1��+oH���  ���0 ���>vSy˖�G�L��(Ϛ��{_�f�rߥ���`�PX0�P鏟��'ƿ�(�H����c�W���όa��&�5%.����3��ܰ�Yg  �8F �%r����J7�?Ξ-E��+���T�)�<\�� �e �?ʿ�q�ϱ�+��{��{œ�)����������d������Ϲ�ޒ<T{ �ͭ.��VK�W��o�񍛲�  @�8� �K��g?�(y�o���Q�2%�o�1���N.zw��2�)�$""M_~��?^�����E��z�O�/����I�����Ͻ�яG��[���O�o%#�J�= Ŧ�%62oީ��E?3�����u   ��a \?�����q�'�ӧˑ$Q]�8���>��ٽ�����n�PX0�ڛ�I�O�'�O�o����P�(6.�tܸz�f͗ۿ��۲�  @�9� ����g>3��m�_U�o�4�dh��ڨ���Sy���
� �q�P�(6�-I��`���%K��y����   # �2��G>�l��[���n���twG�7F���̘������` '��b��)S��W��7<�/��   ?�0 2��������[��##IR�FmݺhZ�6R�gƨ<\�� �e �8y�� �~�P���K�~�㪫�K�g   .�0 2t�����eˆ�ѣ#"�s�ĸ�n�d�t�hƜ<\�� �e �8y�� �~��H[ۙtŊun��ͬ�   �kq 9p�������ͿgΔ�\���k�iݺHK%�jƌ<\�� �e �8y�� �~oWK���ʕ��������   ��q 9��m��L9t�[�]�:"M�4eJ4�pC���w�fL�Ål�PX0 ���j@�����I��G�.}��?���Y�  �7�0 rf�-��Jm���,=�TSDDe��h~�{#imu�fT��l�PX0 ���j@�����ӧ���bův���e�   �,� �CG?��q���v����%.$I��+���u�"M�oF�<\�� �e �8y�� �~oF��l����������   �[�0 r���>vMeǎ�KNK"�<cF4�xc���qg���Ek�PX0 ���j@����ꝝϜ_���l���Yg  ���a ����*o�|{r�t9�$��G�{�1n�{9�F.Vw��2�h�<T{ �M���"mmIW������d�Y   ��p ����}n����Uݽ{~Z�G��M��Gm��H���p���@���Pl�=�Z������ҥ���/<�u   x�F �(s��[?\ݶ��Kǎ�FD���"�o�1JW\�N���5p(,���C����{�H}֬�+V�J��~)�,   �(# `JKG}��ң�����K�$Q[�4���j���\�Åi�PX0 ���j@���iss�������o�ݬ�   @�9� �Q���n�r�з*�wwD�Ʉ	�|�Q�4M��ɕ<\�� �e �8y�� �~O�%I�,8~���g�{����   ���0 ƀC��zGi���.?�ĸ��ʼy�|㍑L��^On��b4p(,���C����{
�>k֋���i��N�Y   �Rr cD:8X:��W6o���ٳ�(���|y4�����{>���Eh�PX0 ���j@���Oss�����}�7�qS�Q   �rp c��;���{��ʻvu$i�ɓ�������O��p��@���Pl�=�Q*E���x�Zu]����   ���0 ƨ#��'���m�'�EDT::���"�6���L���3p(,���C����{
a���L}��;���_�:   \n# `KK�}�����;Ξ-E���ˣ�]V� .�<\p� �e �8y�� �~Ϙ�����,[���?��[��   Yq p���]�l��g�{ۣ^���%�֯�ڲe���>�e������` '��b����r9�00���d�{�}��d�   ��0 
��m��by��?(=:1"�|��|�Q�=['����Ef�PX0 ���j@����9#mmg��+om��?�:   �� (�#7���ɦM�&�OW"I��xq4_w]����L..w��2�h�<T{ �M�g̨���XqO�׾����   @�8� ��J��&m��畭[����V�ښ5�t�U��J:�������` '��b�����tx``�s��q�ݧ��   y�0 
���_[ڽ�����3#"JS�D���G��KO���pA��@���Pl�=�Z������{����ݬ�   @^9�  ""���>��J�>��KO?�Q���n�d�4}���Åd�PX0 ���j@����J�)燗/���>�O��   y�0 xپO��|��7�{��ܹR��Q[�<�����jUo���d�PX0 ���j@����*iSS:�t�_v\y��$����   ��� �q�������,����z$--Ѵ~}Ԗ-�4M�ޖ<\8� �e �8y�� �~��P*E�������Yp�۳�   ��� �:t��6o����Q��h��(͞�C���1p(,���C����{r������ޏw��׳�   ��� ��Ї�]�i�/'�>[�$���@4�������iy�X�
� �q�P�(6��ܪO�z��t����?�լ�   �h�0 xS�~�s�����S�Ǯ��gKI��+��n]D��S���p���@���Pl�=���W^��w�Z�����p�y   `�s �%;︣g��}ZٹsA��$��֨]}uԖ.�T��u���0p(,���C����{r#)���E���[�躙_���Y�  ���a ��~��Iv츻t���Ҵi����Dy�|��ה�����` '��b���\ig�3I�/̻瞿�:   �5# �w��/���Uٲ�ג��j���ttD�{�Ɍz�������` '��b���T}֬G�.�����Yg  ���a �������m��-o����̙r�JQ[�$���&b�x}���G�4p(,���C����{2QomNW�x��k_�%�,   0�9�  ��g>3��gϟ��n].$I��5k�i��H�e����p��@���Pl�=�W����o�0w��3��t�q   �F  w��x�ȶm_)803�4J��Q���-[i����7����` '��b��,�R)��wu���{�ٝu   (� �%3�K�tk�c�JCCS""�W\��]�y�t��Ûn�PX0 ���j@���\r#mmg�K��1��_�J�Y   ��F  ���|��)o����SO5EDT::����#�>])�<��� �e �8y�� �~�%S�:�|,[�{�>����   @�9�  .����G����[6Μ)G����hz׻"ƍ�I
 o��;@a� 4N�= Ŧ��pik�H:0��y+W�B288�u   (:� �e��y��\ڲ���ܹ$ij��ڵѴfM���n2����5p(,���C����{&��ґE���jk�qٽ�>�u   �%# �L�����Ν���s�IJ�'G���Q��4Mu�1(o��;@a� 4N�= Ŧ��%�r:��;4nѢ�ͼ��}Y�   ^�a ���;�!�o�P޷ov�i��M���룲p��2���5p(,���C����{޾R)���?���}h�=��e�q   ���0 ȅc���;~�t�XkDDyΜh~׻�4o��2F��4p(,���C����{޲4"��杪/^���_��W��   �>� @����/��l�X��gk���h��(͜���ryx�
� �q�P�(6���d�����E������u   ��q �N:8Xڶ���-7'�NU"I���M�^ɤI��(��7����` '��b��yS�S���/Y�;z�W��   �5# ��z�S�j9{��ד�[�O^x��r���k"Ə�cF�<�a� �e �8y�� �~�몷�ח,�fǊ7'���Y�   �:� @���gf�����Ҷm+��瓤V�ڊQ�ꪈZM�%��F��@���Pl�=�)7�����+��;3��t�y   ���a 0j}�]�}Wv����$7.jk�DӚ5��JzM���2p(,���C����{^�VK�-�~n��]�Gt<�8   �;�0 uv�r�ږ�������z=J'Fmݺ�-]�~�[yxc�
� �q�P�(6����H��t��wh�����g[�y   ��q �Z�n�������~i��+"M�4mZ4�_��u��Ûb�PX0 ���j@����FD��������ڰ�[Y�   �a 0�������s�o��o��(Ϟ��~w����ur$o��;@a� 4N�= Ŧ�TiGǳ�E�~���{��u   ��q ��?��]ڹ��QY� �֯��̙:O��M0p(,���C������7��H_߯w���e�   ��F  c��?�';w~��{GG4]w��{������@���Pl�}��g�z��dɿ���W~#�,   ���0 ��>���l�zG驧�"I������Ën�PX0 ���j@���P�5�Ŵ��7;x�_f�   ��F  c��|�?T�n�x<�tS$IT{{��k"�:U����b��@���Pl��V�6�\�lٝ<�٬�    �q B:8Xھ�K[�|�t�d�����ɔ):�e������` '��b��Ǡ��i�b`�K�=��Yg   ��0 (����C<�G�-[nNN��D�վ�h���H&O֍.�<��� �e �8y�� �~?��Ӧ��E����÷d�   �� @!=���O8�gσ�;nJN�.�<t_�>�I�t�K /��;@a� 4N�= Ŧߏ��S�%��   ��a Ph����#�<���ץ/�P�r9j�t�5���J������` '��b��G�tʔ��%K���k_3l   ~*�  ��ݴ���[ߓ��B9*�����7P^Dw��2�h�<T{ �M��҉/����+nN���   �� �����-G6mz��c�M����V��%�t�U���P^<w���І!    IDAT2�h�<T{ �M�E҉��/�˦����}�]/d�   F  ��tpp��ƍ���c�5ə3�V�ڊQ[�6��I�z����@���Pl��h��:R�����U�~><�u   `tq �:��ԧZ^<z�Ҏ7&�OW�����Z�U�"��u�� /��;@a� 4N�= Ŧ��X:q��ŋ��2c��g�}���    ��� �7��O}������l��3�s�U�Z-�K�D�UWE��S�	yx��
� �q�P�(6�>��I�./Z�������}�]/d�   �F  �/�w����ԩJT*Q����hiѭ^G^w��2�h�<T{ �M�ϑ�������+nN���   �#  ކ��;�G����+m���ɩS�(����M��E2e�������@���Pl�}ԧM;�,Z�м��%�,   ���0 ���'>1���?���yS�ԩ��C����d�T]�"yx1�
� �q�P�(6�>C������~���f�   �F  4@�����_��+[�ޚ<�TS$IT���i��(͜�sE>���;@a� 4N�= Ŧ�g`���L�x�o��W�Ϭ�    c�� �;|�Ϳ������㏏y�n]������+߼�;@a� 4N�= Ŧ�_&iD���Τ��������F�y   ��p p���Ї�E�޽�)921"���M�\�ٳ����M��@���Pl��%�FD}޼SI�?i���?�:   P<#  .�C������������H�(ϝMk�F���P],߬�;@a� 4N�= Ŧ�_*�R��۟���G��oC�q   ��r p���%{������3�^y�^��4M�|/��7h�PX0 ���j@����V*E}��'�}}��s�=��:   �� ����m�������Wݿn:2���ڢiݺ�,X0���y���
� �q�P�(6��Q������ឞ�ߵa÷��   �#  2r�c���o�]������pR�2%j+WFm��HK�1������@���Pl��;U��#������[��瑬�    ��� �����{�CC��w�Z��=[J&L����Q[�:�V3}-߈�;@a� 4N�= Ŧ߿M���##>6������:�u   ���a @Nl��'�O;q���Ν�%�=WIj��.YMW^��2�{[�w��2�h�<T{ �M���ɓ/��}�eƌ�ϸ���Y�   x##  r&�۲�K�k����Oע\�j__4]uU$S�������� �e �8y�� �~�&էM;�,Z�м��%�,    o�� �;|�Ϳ�����'N�D�D��;���*Jmm����!��;@a� 4N�= Ŧ߿�4"�mmgbѢ����2�<    o�� �Q��G>�b���MM�4�s�F�ڵQ��4MGE��CHw��2�h�<T{ �M�I���tu�0z{?�~�=�u   �w�a �(r�[n�8�ۥ�g��HR�1#jk�D��?Ҝw�<�3p(,���C��������ZZ���w���#6lؔu   �Fp 0
��k����Ҿ}]q�|R�4)j�WGu�҈J%�/��
� �q�P�(6�>"��u����7͝����/>�u   �Fr 0��ԧ�mHvﾦ��s�dܸ�-]�ի#Ə�U��Cw��2�h�<T{ ����>�2���������녬�    \
#  ƀ��;�C�������,?�ĸ�Z��%Q[�:�I�r�������
=�h�<T{ �����>k֋IO���=��-Yg   ��F  �1>��\=t��(M�4�Jww�V��rGG��/�����
9��D�P�(����R)������v���e   �rq 0F���_�<�ۥ���pR�5+j�VEu��H����<Ow��*� ���C����~����ឞC���Oum���    \n#  Ƹ�xo����]�V�/�PNZZ��lY�V��hj�l}0������� ���C����n�om^�౑���w�uב��    d�a @A���-G�l���k��M�~�)�բ�hQ�V��dڴK��P<�
k�` .�<T{ �mL��4"�Y�^Lzz�>wٲۓ���3   d�a @��~��w�m���[#I����ի���i�^�����i�PXcj ��<T{ �mL���\NG��N�̟����w߆��    �� �;|�-�[����,���.$�3��bE���#-���P<�
kL` r"��b�����>�`����Y�aæ��    ��  �_����۷�Sڽ����*Ʉ	Q������7�3�x���� �K�= �6*�}:e�����eƌ�ϸ���Y�   �3�  �,}����C}��o�/��k�J%�FӕWF2}�;�y(�� �5*0 9��j@���~_*�Ȝ9�����k���_�:   �h�0 ��t�[n>t�_T��##Iy��hZ�6*�ݑ��[�y(�� �5z0 ���j@��ߧ�ZZ��J���t���:   �h�0 ��u�;��RyϞ�ə3�ҴiQ[�:j�����o�O�x�V�0 �H�= Ŗ�~�N�|!���ދӧx�����    �V#  xS�v[sr��K{�|����㓦����EmժH�M{�^���i�PX�� �By�� [��}�Y/&==_��l�����p֙    F;�  �e��z�৓��鑦Qio��eQ]�0ҟ�1�P<�
+W�Q.��b�G��V�zW����_���/%�8    c��  ޶wܱ���З�{��NΜ)��L��%Q[�,���]3������1��P�(�L�}:q��Hw��������{ �,    c��  ޱ��;�G����|�t�xk��Q]�0j�WGi��$"������'��b����T��9sN%]]_m�O^��   P0#  h����*ǎ�F�o_Wr�|R�⊨.[���$)�3�f�PX� ��������--#���;����Ԃ���}]   ��s �%��ۮhy��/%{��Pz��Z2aBR�ڊQjm�$��;@a�4��S k��ߧ�Κ�b���[�Y�>2���^��_   ����  .�����|f�޽�zT����re�;:.k!5p(,w���w� d����VK���C����;���/��    �ͩd  ����������L{��X��1��b���4uj�V���%�T�Y�   �`�����,����'߾��{��:    �  \FOO�~�5��[+��y7��_�E���w��h�KOu�>=�    �e�JZ��xr����u}���6v��:    1p �K������:;����X�eK�n��n�JGGT�-�ʂ��JYG   `�H[[�G��vU���������}/�H    �w  2u��5N\sMT��:V8s7m���ϑ�Ձ��-]�ɓ��	   �hT*�Ȝ9�������t288�u$    ^��;  �0\*�zz�==�y�d�o��l��?�AT��_z�{O���   ���q��iO����ٿ�y��=6o�x衬c   �&� �;�'O���}oT��>V��s6n��o|�S�   ��$�3g�X���քi�n�q�ݧ��   �[g� @n](��{}}}}��쳱xӦh}�1Ou   �jm���Y�;�3����}{։    x� O�����h��ڸr׮���Q�Tw   �b*�����t̟����?f�   �1p `T9W��w�.�X�4�O���-[�e˖8���G��+��lYT/����   �5�I##��;Ks�������H<�H֑    h0�  F�#�'Ǒk���kb�ѣ1o��h�����w�����re��O�:&    �@�Z�����oժ���v��?����:    ���;  �^Z.Ǧ�����3Ϝ�e۶Ŕ-[�-�x�;    ������Ԋ��%K�j5�8    \&�  �)O��ķ׭�dݺX|�xt?�h����5�}��Q�:5�x    ���V�{zb��W�ޙ3��   @� �҈�1gN�3'&�tS�ؾ=�o�嬃   �
i�����qb������K��#   �!w  Ƽ��Z��ʕ+WƢ�0<�h�߻7��糎   PX�	���%�uŊ8>qb�q    �	w  
e��ٱk�������]�⊭[�z�xD�f   `�+��lgg]�<6wuE�i�    ���;  ��b��dIĒ%�v�Ll�S�n��ɓYG   sF�O�g��%K��㳎   @�� Px'ZZ�ĺu��Ţ'�{˖��{w$��e   `Ԫ�g-�+V�дiY�   `�0p ���jk�]mm����Ɗ���m�֨ER�g    ���8��GW��M���R։    e� �5��T�{}}}}�v�Ll�S�n��ɓYG   ȕ4Ibx��xf��xdɒ8S�f	   �Q��  �����8�n]�UWŒ�0�o���������   dfx��850ۖ.��[[��   �a�  oV�Ķ9sbۜ9�4<���۷G���##Y�   ���Z-^��CK�ƶ����    0� ��p�R���F����s�bٮ]1}�֨>�xD�f   �q��87wn<�til���R։    �� �:���Y�<b��s�T,޹3�l���'��   �L��ģ�̄	Y�   � � ���O��׭����?~<��m��{�Dr�\��    �P}8�xq�^�<M��u    
��  .�$�s�Ǝ�s������#Gb�c�E��g�   �eiSS���c˗Ǧ���R)�H    ��;  \b#�Rl��M��1���X�sgL߶-�'ND�i��   �"���Ů�8��[�Ϗ�r9�D    �  pY����;˗G,_3^|1�n��w��O�   �V���΍�/�����j։    �a�  �Ѹq��֬�X�&�:}�wǔ;��e   +�$.̜�,]���㹦��   ��2p �8>iR_�6b����я�w��hݹ3J�=�u4   `�I�$�gΌ��Ŷ��xr�#   ��f�  9s`ƌ8p��^���}۶hٹ3��?�u4    �F&O�3}}�cٲ82yr�q    �m1p �;0cF���H��.����;c=��=�u4    �'�龾ؽdI�:5�8    ��� �(��J���=���G��c���1k��h>t(���   \F#&��}}�wɒ�?kV�q    ��� `��P.��zz"zz�yx8�8m;wF��;   �Y�q��Ş�840��̉(���    ���;  �bg+���F�^���Ŝmۢ��Acw   �����������������r֑    ��3p �1�|���ccww4ǲ��m�Ncw   E�&����ű}��H=�   ��1p �1�\�?����5v  ��������1�xql�;7¨   �3p �1��   ���/tu�4joo�:    䆁;  ��c����Xz��Kc�C�"9w.�x   0��L��{{c���qh����    @.� @A��T�====Q��c�cѱsg�߷/J/��u<   F&O�3}}�{ɒ84uj�q     �� �)�b[{{lko��o���y���޵+&��ɩSY�  �Q#M��O�g,��K��Д)YG   �Q��  x�4"�Μ{gΌ�����я�gϞhٻ7*O=��YG  �\I�$�gΌ��Ŏŋ���֬#   ��e�  ��3fā3"��&�?�l�������SOEb�  @Q��q~��xf�����OM��u"    � �7�Д)qh������̙X�kWLٳ'�'ND��Y�  �K�����Ϗ'.���Ϗk��#   ��c�  �-'ZZ�Ě5k�����c���1s��w�`$��e   ���/tuŉ���2o^��YG   �1��  xǞ���{}}}}Q��c�cѾ{w�߿?ʧOg   ޴4I�>mZ�Y� ���ǁ�ӳ�    �b�  4�H����c[{{�M7E��~�{�F�}Q}�Ɉ4�:"   �R���΍������7~�Ғu"    (,w  ��:0cF�1#b������ѷo_Lݽ;����:   �67�َ��Qoo<��/T�YG    ��  ����0!�X�<b��x�\�������HΝ�:   c��ԩq��;/\���"J��#    �b�  d⹦�����#��#��'��ν{�e��(?�tD�f  ��.I��̙q��'�-Z��N�:    �� �̥�r�jk{��y�^s�{.��������##YG  `��77����xj��ؾ`A�ln�:    ��  �s|��8�zu���1~d$=W��������Y�   G�$���i�|GG���s�FZ*e    x�� �\{�\�M����7��'OFϞ=1y߾��8I��uD   .���)�͝���b{oo���%�H    @��  �ʑɓ��ڵk�Ƥs�b`߾��o_49�ٳY�  �RH��1#NwwǑ���5k���   �e�  �Z����""���'���}����!Ow  �<�    ���  ҈�;sf�93b��h�p!����{�D���Q~���#  �z�$F�M��;:�hool�;�S�   ��� �1�L���#��#"�����>x0&��MG�D��d�  ���9�͙�������8�ܜu$     c�  @!�<9��\�re4_�K�YĸC����sY�  (�$�3gƙ��8�`A�5+�S�   ���  �s�Z�Gzz"zz""���g�{���|�PԎ���  �#�&�َ�x��+vvvƩ���#    9f�  ޑ)S�Ț5k�D�^��'��yF�CQ}�񈑑�#  ����8?gN��ꊽ��q|Ҥ�#    ���;  �EFJ�������"֯�q.����c���1ah(�O?��Y�  ȏJ%.̚��Ϗ�]]�k֬�R)�T    �(e�  �:^�VcSggDggDD�x�������{��<�<���I�~'E��-[��6�3�2���v���ޯ�(�A�fQ��b�U̬: �`Ќ���lY2%^D�&�<�v<U�q"�<�>�,��C�whs����Ǚ�w/����  x�*���߸��w�ɏ�]K�応    �ç�   _���t�?y��$���qn}�q�?�8�$�ޘ  �x���\no���o��[�r211�I    �kJ�  ��������N��=潝�l}�I�|�i����p8�   _[}�J.��s��[�護�7;;�I    �B�  ��������v�q{;I21���lݻ��O>I{wW�  �n�2X_��[o���o����I�1�Y    �H�  ��6��pk+nm%��nf��|��O�v�^�ܿ����I]�{&  �&�t������yx�F~���A�9�U     w  ���i�����w�$3�~~kg'�w�d��O�8<L%x  ��v;õ����V]���lm�/h    
$p  ���v�������$���e���'Y�w/��y|�w  ��2��L��՜lo糛7���j�Fcܳ     �Mw  �BON���^��{I��^/�>���;��쳴R�Fc^	  �h49���zί_σ��Ώ��A;    �
�  ��y��+�~����ڧ��ʃi��&��X7  �1��J��՜]����ۂv    �!p  xE<k�����a������?���x�(��ƺ  �f�,h?y��ܿ~=wWW�=	    �!p  xE����xs3?��L�y�~{w7[��e���L��
� �U���bk+G7n��͛y877�I     /��  �5�o6�9    IDAT��V>��J���4G��up��O?���N:;;i���{&  ���������<��Ν��<���*    ���  ����F�����g�O�歇�r�~�>�,�Ǐ��p�+ ��3��Jm-�ׯ���빳���fsܳ     � p  x����������$�T��wvw���Qf<��g���vǼ  ^#U���|�[[9�����f�{    @��   o��N'?��N������$���qn޿����3�����IR�c^
  ��Q����Z�]�������ƍ�LL�{    �+C�  �s�/,���B��o'I������N�<��Çi��Ƽ  �0�����fζ���ڵ|������,    �W��  ����t�o�Nn�N�4G��<<�֣G�{�0S;;i�r�;  ��Q��zi)[[y����ܸ�'���    �Z�  ���]]����/oy��vs�ϲ������t��Ru�c^
  ����`a!����nme����Y[K���2    �ך�  �����D�ϭ[ɭ[_��?}�[��g���L����q2�q%  �r������r���������v�''�=    ��#p  ��73����O�?I25��ݬ��d���t���89IU�c^
 ��f45���z�mn����ܽvM�    P�;   /�E��mm%[[_����y�ѣ�=z��G�D�  �p�v;å�t76rz�jv67swuuܳ     �%�   ���v;?��N���<��vsco��y|<ƕ  �*F�Fꥥ\lm}�������4     ~Ew   �r:1�����yn>|��3��a�i\\�q%  �6j4R/.~~3��V>�z5�VV2h6�=    �߀�  ���OOg��w�w���l��2��������$��1. ��0j�3\ZJe%竫����G���l��=    �L�  �+�xr2�?w��\��{{�w �W�hj*å�tWVrz�jv67���r�Fc��     x	�   �6N'&򣟋�;�Q�f�ѣ�=|���ݴ?N��1.  �<fﯭ�rs3��������̌{     c$p  ��k4rwu5wWW�o;I����A�ww3������4?N��y- �k���`i)ݵ��oldc#wWWs��{     ��  ���7����F~�������e���g�ѣ�<z���a�GGn{ �::�������ի9X]������q/    � p  �/ON�x{;����3���A6��2���ɽ��Ӹ��R ��Z.,�������<Y]���F�Ύ{     �0�;   �+z�F>Z_�G��ϝ������n���r�� �Ǐ�<>N�1- �fԍF���|�������Z��ϧv+;     /��   ~���ٿu+�u����Os���,��e�� �Ǐ�><� 嫪�ff�_ZJwe%O��r���{kk�h6ǽ    �7��   ^�������$7o>w���in<|����L�sx���Q2�g( �FMMe�E�~����++�����Ng��     x�	�  �%؛��������_����\?>���^�2qp���'i��
��bt�J�KK�\[���J���`m-O��qO    ��$p  �1�7��xy9//?w��r��$�g�� �����I��ǩ��1� ��lf8?���B���9_Y���J>[^���ĸ�    ��"p  ���|���O�w�}��le�� 3����}x���IR�cZ �u����b�++�\\����쭮���r��Ƹ�    �!p  �W���d�77�����Χ��l=~�����f��0����NO�^oLk���n�2ZXHq1���./y��v{��     �'p  ���E��;�빳�������ţ��e�� ���T''i��cX ���2\ZJa!���9^]���Z�ͥv;     o0�;   ��~v�{~���$�8;���a��r��0GGi�yz��cX ����hz:ù��#����./���J�--����<     |��  �lwv6����͛ϝW�Q���e��(sO�d�ɓt���>9I��4U�7�� P�Q��zn.���tr������.-���\���'    �+G�   �������|v��!~O����le��(3GG�<:J��8���4�����k��t2��K~>�/"�ӥ�,,���\�h�{"     �V�   ��v<9����ds��k��zv�����no���yv����b �j�v;��l��9Y\����<Z\LO�     /��   x��f�/,����W��>�����i��2{z����tNO�<9I��,��HU�/8 ��zb"���ggӟ�Own.�ss9Y\�Å�<���D     �_�   /�E���++���W>��tq����,e��(�GGi�q~��ӧ�`�WP�f3�+W2�r%Ù��o`_Z���L�fg����Ӊ�q�     ��;   P�~��������$����|5e�ٳ���d��4ӧ��8=M��,���4�>M��Y��h�xQ�J��2���pv6ݹ�\���bq1�ssٟ�u�:     ���   �+�n4� ����/����YV��r�ѣ�5wxخ/.Vsy��Juy�γgM<�xԍF29��+MO�77���\����da!O��?3�~�9�     �K&p   ^?�Fffr03�76��������U/������F���Z��oח��rqq����˳g���e'Ϟ��n�!<�����pj*��t����Φ�J.��sq�J���r4=��+W�Fc�k    �	�  �7�;�����������~o�3�����w�����ŵ��r�������T..ڍ��f���%�x��F#��ff����gfҟ����l�gfr6;�'����     �!�;   �����ov���/����ѻ秧�9�ᷚ�ލ���J�����fsq1��ˉ��]]^6�^O�W�]grrTw:�zj�Wu:�É��LN6&'wF�Tw:��������������h��q�     ^ow   �d�/��$�*�}��x�wq��u�;������u���������J��N�׬��f��U�x��j4�NgTON뉉A&'/���g�N�i��ebb/���a�y����h�����_��ٸg     �<�;   �\����%�_<~%����ð�����6������F5,�۝K�;S�z�U����e��v������7|#�$U�Sgb���G癘8����t:������֏������_�     x�	�   ^�?������|��?��[9;����Ż�7��j0X�z���g�����:��lW�~3�^3�~U.��_GU%�v]w:���ú�֝N/�v/��E����9�[��F��_��{�Vk���|2L~��~�q�     �q�   �ƶ����&���|m�����|�;����ht���_�zk�3�T��T���כ�`Щ��v=6���f��F5$áP�WG�Y��L:�Q�l��f�N�3���~��\֝�eZ���9����<�;�Gu����nҘ�����      �5�   �J������_[���������7�޵�h���`u��5G���p8Q��s�h��`0Q�z4j�כ�꺑~��~�Q�uU���U��*�A��~1o�WKU%�V]�Zu>�n�h�F���j��u�5H�u�V�n6{�v�4������6:��a�qTU�Q�n�j�u���������q�5     �7��   �oT���$������x~py�T��z+Y�3�p8���ѨQ�kIR�U]���p�'�Ѩ��`:I2LV�Q����[��J��������_��U���r�hTU�����W�Q�W�����R�Z_��uU��tFIR�Z�TU]WU�v{�$i��uUՍFcX�Z�$���n�j������$I�u�h4��d�v�4I��:�Z��Q�O�����v�~�l�.������{��g���_      c!p   ���/��b���o����_�����_��u����쏭f�I?��ػ��~�ʕ;��[	�     (��    �Ak��Ivǽ      ^�q           �D�          @!�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @�           A�          @� �3�v,    0��z;�#         ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��         Y�A    IDAT ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��          ��        v��I������tϮ�n7&��s�s1��v�c0���)�`�6�4���(>@���>gFZfd�Ekbq����	�cW� �1UƱ6S������'?s�v.��=����޿��|�  @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�           ���;           �`�          @+�          �
�      @'���    L��;      �	9��    �,w      �677�   ���;      �	�^���    &��      �G    0Y�      @'�R�    �d�      ��s6p   �r�      @'�R�    �d�      ]���     &��      ��    `��     ��xȱc��   ���      �q��w?6�   ��1p      :���?%�   ��1p      :c4=-�   ��1p      :#����    &��      蒧�Rrt    �a�      t�����    L��;      �)�~���    L��;      �)�w   �)e�      t��;   ��2p      :%������GFw    0~�      @�����Lt    �g�      tN)���    ���;      �E?SU��N   �)�      �E9p��3�#    /w      ��z��/E7    0^�      @W�rt     �e�      t�E+++O��    `|�     ����z/�n    `|�     �.{YUU�=   ��=      @�=z0<':   ��0p      ��e�    ���;      �u���:   ���      ]������    v��      輜�n    `��     �i���p���    v��      ��    ���      S!�|�k����    v��      ����_��    `��     ������������    쌁;      05J)�y�/��    `g�     ���s>�    ���      ��Y���?   ���      Sg4]�    ���      ���~Nt    �c�      L�+�    �w      `Z�|]�?   ���      S+����    ���      �Z��_\YY�$�   ��1p      �Y��z�>:   ��1p      ��/��gFG    pn�      ���9��    ���      ���/��    ��      3!缼���/�   �{g�      ̊=}�����    ���      3c4������;    ���     ���s~���ܑ�    ~0w      `�\���tat    ���      �5�����EG    ���     ���s��+++?�   �w3p    ��666F� 0f����������    ���    �s����� 0O>y��GG    ��     �S�y#� &���UkkkEw    �m�     ��h4r���TJ9�����   ���    pN�^�w �ً����#    0p    `677]p`��z�7�Ã�    ���    �sr��iWJ����:�   `��    pN.�0�J)��u���   �Yf�    �9����؟s~������   �Ye�    �9��}w fB)咓'O^�   0��    8��'O��  {%����p���   �Yd�    �9UUuwJi3� ��y�^����}�!    ���    ��r���QJ��ԩS�Gw    �w     ��Lt  �j8>%:   `��    �U.�0k���z׭���   ��     l�� ̜R�%�N��<�   `V�    �U� ̪juu���    ���    ���+:  ��7��[U���!    ���    ��r��Y���`put   ��3p    `KJ)�  �~�i�DG    L3w     ����}#� ��R��VVV   0��    ؒ�h��� ���z�(���   �id�    �V�� ����iGG    L#w     �$��; |�����ӣ#    ���;     [RJq� ��^�����D�    Lw     ��� �ۓ<XGG    Lw     �d4����9����Ew    Lw     �����ut �ԛ��֞   0�    ؒ3g�|#�4�� �lnn^_UՁ�   ��3p    `K���(�|=� Z����o��    �:w     �,���� �V����u���   �.3p    `;�������%�    ]e�    �v��};���]�����   �.2p    `�r�� pn����{g)%G�    t��;     [VJ1p��ya�4�EG    t��;     �a� [�����   �%�     lY��+� �!�RJ�?8:   �+�    ز�h�; l��^�}�����   �w     ��̙3�REw @��R.)��5�   ��    ز��Φ�\q�m*���i���   ��3p    `[r��  ]TJY����;    ���    �m)��yt tT/�������F�    ���;     �b� ���h��cǎ�?:   ���    خ;� ��p����J)9:   �m�    خ�  S��M�\   �6�     lK)�w �j8�4:   �M�    ؖ���Δ�(� �@�9��i���   hw     �����9�/Gw ��8��rC]׏�   hw     ������ �"O)ݴ����   �h�     l[��� ��I�~��UU�E�    D2p    `�F���; �Y�������   �H�     l�� 0���M��Zt   @w     �mcc�� &��rm�4/��    �`�    ��=z����NGw ���R޽�����   ��f�    ���KJ�O�; `�͏F�����   ���    ة/F ��{d�߿imm��!    {��    ��9��� �O�Fׯ���   ��     �H)�D7 �,(���ӧO�����[    &��    ���z��n �YQJyi]ׯ��    �4w     v��K/�RJ�dt ̊��UM��Zt   �$�    �#9�R��� 0KJ)��u���   �I1p    `�J)��n ��O)�{8>3:   `�    ر���; ���?�����   �q3p    `7� �Cz�ލǎ{ht   �8�    �c����|J�Dw ��z�ٳgo][[{`t   ���    �c�>�R�3� f�ś����رc�E�    ���;     ��G� 0�w�=�\_U�\t   �n�    �[  �����`��RJ�n   �w     v%�l� ���_   ��     �������F� @J9�W7MsYt   �N�    �+G�=UJ�bt �m���i��   ��     �Z���E7  �_.��v0k��    IDAT�4�8:   `��    ص��F7  �e_J����yVt   �v�    �k� �>��������-    [e�    �����}.�t6� �>(�|���'D�    l��;     �v���o���{t ��r�M)ݺ�����   �s1p    `,J)wD7  �����cKKKF�    �w     ��� Z��r����G����n   �7�     �E���)�� ܧ�ollܲ�����   ���    ��XXX��RʟDw  �t�h4��o|� :   �{�    06�^�� `K~������:?:   ��2p    `lJ)��n  ��y����UU�   �[�     �M���Tt �-��<~�x?:    %w     ���K/����W�; �m9t�ĉ��  �60p    `�>  l��N�8񶪪�!   ���     `�J)�E7  ;���`�#w    �     �U���� `�~e0��Rrt   0��    ����;SJ_��  v�MӬEG    ���    �I�-:  ؕW��jt   0{�    �R��; tߥ��p   �w     ��{�-�4��  v'��4�U�   ��0p    `쮼�ʯ��>� �^)�u]_�   �w     &��r[t 06����?DG    ���    ���9��  ��뚦�*:   �n�     L��ӧ?�R:� �O)�F�   �$�    0UU��9�� ���;   0I�     L҇� ��+�������   Lw     &fcc�ƔR��  &�5F�   ���    01G��rJ�� �ļ�i�߈�    ���;     �vct  09����   w     &j4��  L��;   0.�     L�E]����7�; ���#���   ���    ��C�m�o��  &��r���7�Rrt   �M�     L\)�� `������zUUޣ  �m�C    ��;}��M9绢; ��QJy����;����n   ���    �����Rʭ� ��)��t0�k}}}_t   ��     쉜�� ��;t�ԩ��:?:   �w     �ķ�����6�; �=��auu�~�!   @��    �'���ʯ��>� 콜�ύF������[   �v3p    `ϔRn�n  �<���߶�����   ���    �3����)�� �����͏�   ���    �=s���/��>� ��9���h�������   ���;     {��r}t �I���[]]}Dt   �.�     �R���ft �GG��kkk��   ���    �=u�ȑ���>� ��E���c+++��   ���    ��G  �PJ����}r8>%�   �g�    ����z�K)���  Z��9�ۚ�yZt   ��    �=w�e�}#�t[t �*+�||8>#:   �c�    @�� ��y`��#+++ώ   b�    bcc��)���; ��y@�׻��럍   ���;     !��⊿I)}(� h�AJ�4M��   `o�    ��r]t �Z�K)����   ���;     aΜ9��W�; ������>   �w     �TU��RzOt �j9���4�R)%G�    �e�    @�R��D7  �WJ9�4�۫���n   &��    �P���_H)}.� 脗�߫����   `2�    h�� ��x�`0�qyyy>:   ?w     RޕR�'� �����[�����C   ��2p     �����RJ7Gw  ������}ee���!   ���    �
���E7  �sq�������c�C   ��0p    �Μ9scJ�/�; �����h���pxqt   �{�     �BUU)��Gw  ����Ǜ�yVt   �;�     �����[RJ�� @'=��rK]�Ϗ   v��    �ָ�+N��n��  :�`J�MӼ$:   �w     Z%���� ����R�3_   l��;     �r�ԩ���2� �~�y���#�!   ���    �*UUm�7� 輜RZn�f����c   ��1p    �u677ߒREw  �WJ9�4�o?~��   ���;     �s�ȑ/�Rn��  ��+N�8qCUU�C   ��f�    @+���  L����~Ht   p��    h��/�����; ���R�'���.�   ~0w     Z)�\J)o��  �K���sss��G�    ���    ���FoK)���  ����9|ee�'�C   ��f�    @k=z�T)�]� �TzP���h]��$:   �w     Z-����R��  ��y)��6M�C   �o3p    ���8���� `j�K)on�f):   0p    �J)�F7  ӭ�rt8�������   �e�     �����SJ� L���N�8�����E�   ��2p    ��r�%���� �Lx�������   ���    �N8}��;RJ� L���Omnnޱ�����   �5�     tBUUw�R֣; ����~�G]�O�  �Yb�    @�K)� ̌G��>������   ��     t�����RJ��  fʃ���-����C   `�    �)��ՔR��  fG)�@������-   0��    ����/�?� ̜~�y���+�C   `��    �9��h9� �I9����i�ZU�\t   L#w     :gqq����g�; ��TJ�����﫪�@t   Lw     :����  ̮Rʋ��ǆ��â[   `��    �IL)}!� �i?�s�l�4��  �ia�    @'�K�y9� �y�)�|�i�gE�   �40p    ����G�'���� �̻��rK�4/�  ��3p    ��:��s^��  H),���i�WE�   @��    �i�������W�;  RJ�Rʛ�������c   ���    �Ç+�� �J)���y������   �w     :o4�VJ�k�  ��O�:��cǎ�?:   ���    ��[\\<�Rj�;  ��O�={�����GF�   @W�    0J)oL�� ���~��_�����!   ��     LW��{D���u]?7:   ���    ���; �bJ)�2�it   ���;     S�w ����9�{8�  ��2p    `��� �\�9/5MsmUU��  �{�X    `�,..�)���  ���rx0�����[   �M�    �FoJ)}5: �^2??��W_}At   ���;     Sgqq�LJ��� �s)�<{����4��[   ��    �J�O�^O)�Yt ��H)�3u]?':   ��    0���:�Rzmt �]�R��p8<   ��    �Z^x�J)�qt ���s~o]�G�C    ��;     S�СC�)���;  �!��������*o�   ��     L�����O)�At �v�R��Ͽ����-   ���    ��� �SJ���`p�p8|Xt   �w     �����GSJ�Gw  ��3r����{�����<���Tw��B% ���"�����^���"Xd!�lS��݆��H��:�s:)�ڄx�!�
F.I 	$���d���2��*�m�ꮳ�p$�tWwW�>���/x���k}�~�p8|T�   �	�     ̄�hԍ�Q� ����h�����'�  ��f�    �Lؿ��RJו�  8Kj�Z��  ��d�    ��h�Z����Kw  ���RJ���t   lw     f����G#�5�;  �AJ)]�4�k���+   [��    ���n�2"��t ���9�laa��UU=�t   l%w     f����?����  8W9�����+�8�t   lw     fή]����?/� ����ɓ�o��KJ�   �V0p    `��۷��xU� �-�Ȝ��u]c�   8W�     ̤n�{]D|�t �yPD�s0,�  �sa�    �LJ)��DD.� �E�R�n0T�C   �l�    0����sοT� `����u]_]U�\�   8S�     ̴v�}0"���  �b/]XXx����B�   8�     ̴N��)���  [-���v�}�p8|x�   �,w     f^J������  ���F�9r�1�C   `3�    �y�N�Μ��  ��666�?��t   ���;     DD�߿>"n)� �M>'��Φi^P:   N��     >e4-EĨt �6ٝs���`�C   ��    ���߿�wr�W��  �F)�t���k�=��t   �G�     �i���e9�/� ��^���������  �Og�     ����|<"^U� `<e}}���i.(   ���     ���Ǐ_,� ��"�|�����K�   @��;     |���F��(� �>��j�2�^:   �    �^�z�ߎ�kJw  쐅�h����e�C   �m�     pZ�֏F�?��  �!s)������9��1   �&w     ��N����  ;(��.o���G��U:  ��c�     �p�ر�E��;  v����ޱ�����!   �w     8���F�V�"�D� �������>|xo�   f��;     �F���p����  |����+++_U:  ��`�     �p����#��Kw  �V����i�Q:  ��g�     �PUտF�+Jw  2�s~[]�//  �t3p    �M��z7��R� �������i��9��1   L'w     8sss?�\� ����i�TU��J�   0}�    �,--�uD�X� �¾g~~�7�9�٥C   �.�     p�������?Kw  �-�>|xo�   ���;     ����ōV��҈X/� P�c���>X��J�   0�    �,t:�G���  c��ަi�Q:  ��g�     g�رc����/� 0�sο�4�+J�   0��    �,UU��s~IDl�n ��k�����*{   Ί�     �A���`J��  �"�oϞ=�����n  `��    �9Z[[�ш���  �"����ht�����n  `��    �9���_s�/��\� `�|�������ˏ.  ��0p    �-���o���/� 0f�j�n_W:  ��`�     [��ɓ?Q� `���>/�t�`0��t   ���     �����%����  c輔ҵ���*  �x3p    �-����o(� 0�RJ�򺮯��j�t   ���     ��ɓ'/���[� `L�t~~������C   ?�     ��<�/�ȥ[  ������m��ˏ(  �x1p    �m�����/� 0��n��h��+K�   0>�    `��޽{)����  c��9�[����K�   0�    `��۷���ȥ[  ���h4z[]��  �<w     �F�n�Ɯ�kKw  ����Ʀi�[�   �2p    ��׍�?. 0�R��'�~�ѣGw��  �w     �f�~�x���#b�t ������>�Y�C   �y�     �����9�å;  &ē������ὥC   �Y�     �C�?^E�o��  ���������'�  `��    ����d��~aD�Y� `B<,"��4�3K�   �3�    `---�aD��t �ٓs~k]�?T:  ��g�     ;�رcWF�M�;  &H;"�j��ʪ�l   ���     vXUU��'O�("��t �$�9�������n  `{�    @�XJ饥;  &�����o^]]���!   l=w     (���%"�P� `}�����M�|I�   ���;     �s~eD�q� �	�Ȝ��~b�   ���;     ����G��#b�t �zpD�g0\T:  ��a�     ��z�ߎ�/� 0��K)];��!   �;w     ǎ;7��  �P)�ty�4���j�t   g��     �@UU����F�?�n �T9���Ͽ}yyy�t   g��     �ā�""^^� `�=��n߸�����!   �9w     #�^��9�)� 0Ὰ�j�~�ȑǔ  ���    ��9��RJ�S� `�}��������7�  `��    `��۷����"��[  &��F�w��  `s�    `u:���_V� `
��R���`P�  ���    `L����s�GKw  L��R���뫫��+  �}3p    �1v���K#�wKw  L��.,,�����  ���    ����V���(� 0r��9??�`0xH�   >��;     ��N����Jw  L��I)ݾ�����!   ܓ�;     L�~�}J���  S�����~b�   ���;     L����}�;  �ȃ"�݃�`�t   �d�     ����F���"��[  ���RJ��W�  ��     &�����$���;  �L;��SM�\YU�-  @A�2     �0�n�M)�kJw  L���={�\?�_�  `V�    �Z[[{eD|�t ��I)=g4�X���n  �E�     0����k4-F�Z� �)�u9�[꺾�t  ��1p    �	���?�9�@� �i�RzLD�Q��J�   �w     �`�~���xm� �)�Ј�y8>�t  ��0p    �	����ʈ��t ��Z�Fo����C   f��;     L�K.��D��^���*� 0���3M�\�sN�c   ���;     L�����N)}OD��n �V9�}u]���ѣ�J�   L+w     ��n�9��;  �YJ�����n8|��g�n  �F�     0E�����  S��sss�5MsA�  �ic�     S��j�PJ�wJw  L�/�9߱�����!   ���     �L�ӹ3�����[  ���Z�[�~Z�  �ia�     S������x~Dl�n �r�kMӼ�t  �40p    �)����U� ��;�����*  0��    `�u��W��R� `����u]_SU�\�  �Ie�     S,��G�ы"�J�  ̈/,,�cyyy�t  �$2p    �)w�������O�n �9秶������K�   Lw     ������ED.� 0#���ɓ��u���C   &��;     ̈~����X.� 0C�0"޿����!   ���     fȱc�^�s���  3�A�V�݃���!   ���     fHUU�'N� "��t �9/��Ku]�H�  �qg�     3��.��V����-  3�W�u=���^  �>8�     `u:��o�Zϋ���-  3fi~~�W���_�  �qd�     3����fJ�`� ������7>|��J�   �w     �a�n�N)]]� `}���������t  �81p    �7??�����Jw  ̠����+  0.�    `�]r�%'N�8����-  3��SJ���K�   �w      .����O�n �A����h��    IDATC   J3p     ""����AD\�[  f�y)�k��yE�  ���    ��������t ��j�_�4͕9�T:  �w     �z����5�;  fU�y_�4o<z���-   ;��     �kkk����Kw  ̰����nX]]}`�  ��d�     |����{vJ�c�[  fؓ���o�/  �S�    �{u饗�����wF���-  3�q�������G�  �	�     �}ڿ��r�GĨt ���v������o(  ���    �S�������  �qj���j�晥C   ���;     pZ�n��)�kKw  ̲��rο:^R�  `��     ��Rʻv�zqD�R� `�ͥ������J�   lw     `S���ww��zvD�Q� ��"��������J�   l%w     `�:���s��[� �x�������K�   lw     �����?o�Zό��[  f]��;G��M�zp�  ��`�     ��N��RJE�F�  �kw�������G�  8W�     �Y�v�o��~�  ""��v�����G�  8�     �Y��zGRJ��;  �����������!   g��     8'kkkK)�_-� @DD<(����i�Q:  �l�     礪�QJ�{#��-  DDĞ�����KJ�   �)w     ��u:�;#�Y��-  DD�\J���`P�  8�     ����z��n��#"��t  �RJ�7MseUU6"  �Dp�      [fii�#�"���-  |R�y����/TU��t  ���     [���ݒs���ȥ[  ��������oX]]}`�  �S1p     �\�߿.�ty�  ���}��7���  �/�     ���v��="~�t  �.���SJ���G�n  �7�     ��YXXؗRzW�  ��F��-+++�/  ��     ��K.9����숸�t  ��V�u����SK�   |:w     `[UU��9�?)� �=̷Z�_�����C   ���;     ������土]� �{8/"�k���!   �     �����j���T� �{h��i�åC   �    ���t>�j��w�n ��r��������I  �b$     ���t:��9_�[  ����+~��ѣ�J�   ���     �q�~�m)�W��  �3土����W]u�|�  `��     Et�ݣ��;  �W�z�w�x�С�  f��;     PL�׻<����  ܫ�ٽ{�-��ˏ(  �w     ��.��Ҝ�[Jw  p����n��4͗�  f��;     P��������_��n �^}A����i�S�  `��     �UUu��ݻ�*� ��:?�|K]�O)  L7w     `,�۷��-� �����_�����C  ��e�     ���U��zJD�]�  ��yq�`0xY�  `:�     c���|$"��J�  p��)�����*  Lw     `��z�ߊ�ň8Q� �{�RJ��A�9��  ���;     0�z��qQDl�n �ޥ�zMӼ��ѣ�J�   ���     [�^�D�K""�n �>]������px��!  ��3p     �Z��{c����  �ҳF��o���>�t  0��    �����W#�'Kw  pJ߸��~�����  &��;     0z���9Kw  pJOX__�eyy��C  ��d�     L�^��K)]S� �S��v�}�����  &��;     01RJ��.�$"~�t  �ta�պ�i��,  Lw     `�,..n;v�qC�  N����{�����!  ��0p     &NUU�ǎ{nJ���-  ��g�ߵ�����!  �d0p     &RUU�z�ĉg��~�t  ����j�z]��-  �?w     `b<x�_v�������n ��vG�uMӼ�t  0��    ���o߾��FO����n ���9��5M�)  �/w     `�8p�/Z��S"�oJ�  pJ)��4Ms�t  0��    ����t>�j��/� ����u����lW  �{p$      S���|8����8V� ��zŞ={�XU�\�  `|�     S���0��숸�t  ��Rz��={�[]]=�t  0�    �������w�n ��RJ�Y__�ayyy�t  P��;     0�z��;#⢈8Q� ����v�}�C�\:  (��     �Z�^�)��#b�t  ��ջw��+�8�t  P��;     0պ��r��#w �I�'O���i�J�   e�     S���_�RziD�J�  pZ_�s�u8>�t  ���    ����v��DD.� ��]8�n_^:  �Y�     ����z�����  l�CSJ7���<�t  �s�    ������L)uKw  �)i�Z7��+  �w     `�t��a���Kw  �)��Rzw�4O.  l?w     `&���*"��  `S�Dį�ç�  ���;     0�z�ޫRJ˥;  8���F��ۚ�yN�  `��     3����hD\U� �Mٝs~S]�/,  lw     `���r�������-  lJ;"~��뗖  ���;     0�>5r���x]�  6����z�t  ���     �#��{��<�tm�  6%Eİi��K�   [��     �S7���^�s~K�  6'�\�u���  ��0p     �4UU������\� �M���뫪��� �	�Q     �,..n�ݻ��0r �$?4??��믿�]:  8{�      ��� `"]���}��=��t  pv�     ���������s�o)� ��]t�ر7UU��t  p��     N�K.9q�>/�� 01r�Ϟ��kUU�+�  �w     ��X\\�ػw��a� 0I�m~~�������C  ��3p     �#w ������������!  ���     l��; ��I)}�]w������[  ��3p     8F�  �'������VWWX�  85w     �3d� 0yr�߰��~�p8|P�  ��     �#w ����:���!  ��3p     8K�6rO)][� ���9��ݻ�S���n  >��;     �9X\\ܸ����� `�<>�|ˑ#GV:  �'w     �sd� 0yRJ���ظiyy��K�   ���     `� L�/m��7�Ç�  >��     `�,..n����0"�T� �M{�h4�yyy��C   w     �-UU�ɽ{�~oD��t  ����v��#G�|Q�  �u�      [lqqq���("~�t  �v�h4�yee呥C  `��     l��R�v�����*� �����Z��WVV��t  �*w     �m������(� ��]�j�n��-  ���     `}j�+�[  ش�G��{����!  0k�     v@��;�s>X� �M{hD��'w  �Y�      ;���/� L���F���� `��     �~����  l�CF�эu]Y�  ��      ;���5��K�  �)�G�MF�  ���     
��z?�s�$"F�[  ؔ�#�#G�<�t  L3w     �B����9�#�d�  6����#w  �F�      ���k�� &�C766�5U:  ���;     @a�~�����#�D�  6����敕�G� �ic�     0���䜟w�n `S�j��� `��     ��~�����s�� `R\�n�o_X:  ���;     �����h�ZO����-  �^�yoJ�}G����-  0�     �L��y_D<9">^� �M�`4�l�  ���     `�z��J)}k���K�  pz9罣����`���[  `��     ��n���)�o���,� �����Z��� ��3p     c�^����'Fğ�n ��r�{SJ79r�J�  �$2p     sKKKm��O���/� ��\����^#w  8s�      `ii�����W� �M�pcc������C  `��     L�K/��o���7E��[  ؔG�F���9��!  0)�     &����?真7�n `S�xcc㝇zp�  ��      ���߽{�����V� �M��ݻw�g8>�t  �;w     �	�o߾����#�ͥ[  ؔǏF�w,///� �qf�     0���Z߻w�E���-  l������p�UW͗ �qe�     0�7���KRJ��[  8���7�y睿ZU��J�  �82p     �p)���t.�9ץ[  ؔo�������y�C  `��     L��R��������-  l��N�8��UU͕ �qb�     0E���rJ��t  ��s~��={^_U�  |��1     ���v�ÈxaD�,� ����^0??��;  |��1     ���z��s~nD�U� �������+KG  �80p     �R�~�m)�gD�Z�  N-��ʦi���  ���     �X�۽9"��P� �S�9_Z�����  ���     �\�����������-  �֏�u}Y�  (��     `�z�?h��O����n �^=��#  �w     �������h������-  �ZJi�i�,�  ;��     `��߿�oZ�ַD�K�  pJ)����i��t  �$w     ���t>�s~rJ�]�[  8�V��皦���!  �S�     fP��?������xs�  N��s���p���!  ��     fTUU�{��(�tM�  Niw��-u]?�t  l7w     �������t^�s�K�  p�r�������<�t  l'w     ��R��~��s>X����w�_�_u�ǿ��NubW	�L�f��:��B!�$�@� �bA��P�u��Wݝ5��'��ΩN"QCX�ED.��%
�B�$0r]�Iw���@����RU�\^�������� �Nݭ�j�����D�  �(�      DDD]׋)�GĠt  w�^9�w-..�Z:  6��;      ��v���s~vD)� �z@��~ϥ�^z��!  ���     �����M)=%"�n ������;�����!  ���     ��n�����#���-  ܡ�:t菚�9�t  �w      nW]��j�Ί�/�n ��===���i�� ��`�     ��t:��n�ψ�,� �z����5M�� 0��      ܩ����mٲ�̔�GK�  p��=33sE�  8Q�      ܥ�;w~��O>+����-  ܾ��Kz���Kw  ��0p     ��رc����O���J�  p�����N�  8^�      ��io߾����ե[  �}9�^�����  p<�     8&���ku]�(缻t  �+�_����Z:  ���;      ǥ��Ŝ�K#bP� ��h眯ݷo�y�C  �X�     p��~eD<'"��n �6�Z��u�~���C  �h�     pB�������q�t  ��Ã������{P�  8�      ��n���"�1��-  �ZJ鞭V�]�_~���n ��b�     ������������-  �Ə9r�W]u�t�  �3�      ���������>*">Y� �[K)=�СCok�f�t  �w      ���ݻoh�Z�GćJ�  p�����&�J�  ��1p     `�u:���ύ�w�n �6~yyy���  ��c�     ���������'F�5�[  ���󞥥���;  ��     �a��Y�v���9�-� ������~��Jw  ��3p     `C��r]�MD쌈A�  �M+���^�wn�  �w      6EUUWD�s"�p�  n1o޷o�ϕ �w      6QUU��s>?"�U� �[�p��z�����C�  0p     `S�u���8;"�R� �[�����ޥ��{� `��     �骪�H����-  ��)�?^ZZ�V: ��e�     @u]v˖-g��>Z� �[�BJ�MM�l) �d2p     ���;w~��O>+����[  ��۶m{]�9� `��     PԎ;Vn��'E��n �_���������  `��     P\�4�WVV��R��t  �*���^����  Lw      �B�4�n�;;#bP� ���xe��b�  &��;      C���+RJGđ�-  D;���}���\�  &��;      C���1����8X� ��i�Z�����+ ��3p     `(�u��V�uN����[  �Ss�o�ꪫ�K�  0��     Z�N��[�lyDD|�t  �s�:�4͖�!  �/w      �����g>|ZD|�t  q����  `|�     0�.��s��F�;K�  L���z��|�  Ɠ�;      #��뛶o�����kJ�  �^����  �w      F����Z��ya�yo� �	׊�7���G� `��     0RRJ���&����X-� 0�No߷oߏ� `|�     0����5)�����]� `R���R���.��GJ�  0�     Y�n������WK�  L���Onٲ�M�L�n `��     0���˜�i�O�[  &UJ����W��  `��     0�>=�H)}�t �{n�׻�t  ���     ������O>���xW� �	���~�Y�#  ]�      ��;v����<1����-  *�_���]: ��d�     �Xi�f��� 缷t ����9_����t  ���     ���R�u]71��9  ��9��߿��C  -�      ����~;"��J�  L����h�fK�  F��;      c������F��K�  L�sgff�JG  0:�     {�j��*� 0ir�;{�ޯ��  `4�     0:��?�3s�]� `�ryy���  ?w      &���"�#��S  &�I���-���@�  ���;      ��뛶o�~a��wK�  L�{�������Ҷ�!  /w      &����Z]�/���1(� 0A�j���4��  �ˡ     �Ī�ꊔ�3"�;�[  &E�����ӯ(� �p2p     `�u���r�D�7K�  L��---=�t  ���     ��W���[��#SJ7�n �)�tM�����!  w      ��N������E�ߔn ��D��O- ��0p     ��ڵk�?�r�)gFĻJ�  L�S�������ʭ�C  �      �}v�ر����Ĕ�kJ�  L��n���W��  `8�     �h�f���0缷t �$H)=���wJw  P��;      ܎�R���9�jD)� 0�r�K�~����  �,w      �u]�.".��o�n s������?]: �r�     �.TU�ވ8;"�T� `����^v�e?R: �2�     �(TU��v�}Z���[  �܃N:�h� `��     �Q��������#s�(� 0�ι�^^: ��g�      �`Ϟ=�غu�c#�J�  ���---=�t  ���      �������n��s����    IDAT{K�  ���R�fyy���C  �<�      pRJ���&"^��s  �����.--m+ ��0p     �PU���9?-����-  c�gRJ�) ��0p     �T����_)� 0�.��z/- ��3p     �u��t>�n�O��,� 0�����;�t  ��      �����g>|zD|�t �:��jX\\<�t  ��      ��%�\r���ʹq�t ��w��~s�4S�C  ��      �Κ�����۟�Rze� �1t����b�  6��;      l���ٵn��҈���=  �$缳��?�t  ���      6PUUW��f#�;�[  �I��U�~���;  X_�      �����[r�gG��J�  ��Sr�oڿ��K�  �~�     `�u��v�}fD\_� `�<hmm������ ;      �$���o�ۧE�ߔn #O����S: ��a�      �h~~��9�3"��[  �E��7z����;  8q�      ��꺾iee��9�K�  ��VD����ݿt  '��      
h�f���E�Έ�� ���뚦�* ��3p     �����"�4�J�  ������Y, ��3p     �º��[rΏ�9�t ���9��^����  w      u](�|ZD�c� ��"����@�  ���;      ����O>|���`� �w����7]y�[K�  pl�     `�\r�%7����o*� 0�RJ;|��R�  ���;      ��i���v/�9�-� 0�^������  =w      B)�\�u;#b�p ��J)�jqq���;  8:�      0Ī��"��K)�o�n Q3�v���9�t  w��      �\]�oM)=:"�\� `D=tzzz_�  ;      ��N����i��-  #�%�^���  �9w      u]�ȑ#��?P� `������ݿt  w��      FȞ={��u��Ǧ��-� 0�~$���K�  p��     `�������t��s�[� `������?��Jw  p��     `��r]�MJ�yq�t �(�9�|ii���  ܖ�;      ��n�{MD\�*� 0BZ)����z?Z: �[3p     �WU�{[�֣"��[  F�}rί�9��!  �w      �N�c�������/� 0*RJ����/)� ��1p     �1�{�����N��w�n !K�~�!�#  �W�      0Fv��upee����-  #bk������SJ�  `�      c�i�ժ�^�s��t ����`pY�  �     `l�u�ύ�å[  F������#  &��;      ����^�s>?"��t ��K)�k.���+ 0��     `��u��V������t ��������rΩt ��2p     �	��t���n�)� 0��_^^���  ���      &����s�gE�;J�  ��^��KG  L"w      � u]ߴ}��#�wJ�  �����~�i���-  ���      &����ZUU;"bgDJ�  ������iJw  Lw      �PUU]�R���C�[  �Q�yW��;�t �$1p     �	��v�27�n B��x���Ҷ�!  ���      &�����G�'K�  �F�R� �Ia�      ���§[����g�[  �MJ�E�~��;  &��;      �N��SSS祔�-� 0dR��5�����t ��3p      n177ws��yV�yo� �!s�`0xM� �qg�      �JJ)�uݤ��GJ�  ��,--=�t �83p      nW�۽&�����f� �a�R��~���  ���      �Cu]���j��/� 0$�>^U: `\�      w���|��n?<��ץ[  �AJ���~�WJw  �#w      �.���1"~1"�^8 `(�/����+� 0n�     ��R��M۷oJD�v� �!p��`��  ���      8j���kUU�E�ΈX+� PRJ��^���  ���      8fUU]OK)}�t @aW,..޷t ��0p      �KUUo���#��[  
�[��~U� �qa�      �n��w�V��[  
����]\: `�      '�����v����J�  t����}KG  �:w      �������֭[וn (�n�v�wJG  �:w      `]������v�K�[  
yB��z� �Qf�      ���R��j!"vFĠt �f�9���+��g� �Qe�      ��������G�wJ�  l�=|��m  ���;      �!��zs�����f� �Mv�}��+ 0��     �S���[����-  ���j������.� 0j�     ���t>�n�ψ�O�n �D�������t ��1p      6�����Z��##⃥[  6KJi����i�;  F��;      �):��ק��Ή�7�n �$����W_}�I�C  F��;      �i���n޾}�3"�ե[  6�Ϭ��,��  �      �����]���9���K�  l����\� `�      E�u�ύ�#�[  6��-[�\Y: `�      �TU���� "�n �H9�󖖖�Q� `��      EUU�ވxLD|�t �FJ)�߿��Kw  3w      �������n��*� ������#  ���;      0���?�e˖3"�#�[  6Я///�B� �ae�      ��;w~9�|VJ�=�[  6Hk0��i�-�C  ���;      0T꺾����O���J�  l��ݶm�KJG  #w      `�4Msx�����^[� `#��~cqq�;  ���;      0�fgg�:��r�{K�  l��v��/ 0l�     ���R�u]7�3"r� ��6���[: `��      C���+"��X-� ��r������Jw  w      `$TU����S#�P� ���R�ɃΕ�  �      ���v�oo�Z�GķJ�  ��W,//ߧt �00p      FJ���@D�_)� �Nf��b� �a`�      ����>�n�O��O�n X'�����#  J3p      F����g�����-  �!��ʫ�����  %�      #k~~��G�9+">T� `����_\: �$w      `��ٳ���r�y��-  �`���ҽJG  �b�      ��;v����\J�  ���E�o��  (��      M�޾}�3s�W�n 8)��/--�l� ��     ��1;;�V���rλK�  ��vJ���  %�      c���ň���A� ����^�wa� ��f�      ����~;�tqD)� p��W^y���  ���      [�n��)��E�ͥ[  ���9���  ���      k�n��9��E���-  �*���}��ݻt �f1p      �^]��;"�,� p�fRJM� ��b�      L���>�j�Ή�K�  ���󗖖~�t �f0p      &F����v�}FD�s� �c�N)�+ ��     ��2??���"⳥[  ��c{�޹�#  6��;      0q������/FħJ�  ���il� ����      &��ݻogF��J�  �����<�t �F2p      &����9rVD|�t ���9_�4���  �(�      �D۳g�7VWWϋ��S� �(�gzz�%�#  6��;      0�v���͜�y���-  Gaϥ�^z��  ��       "꺾ijj�	��-  w��[�n�o�#  6��;      �w���ݼ���􈸮t ���9�xyy���;  ֛�;      ��i������/�9�^� �;1�s�[: `��      ����ٵ��~%"�(� pGr�����)� ���      nGJ)WU�3���K�  ܁VDx� +�       w����w��  �=9�'---�V� `��      ܅��SJ/��\� ���~�t �z1p      8
�n���xQDJ�  ��3���cJG  �w      ��TUիs�ώ���-  �/�|Y�9��  8Q�       Ǡ��k#⢈8R� ���|��{b� �e�      p���zsJ��N� ��I)�f�46a �Hs�       �n��')����; 0<�����E�#  N��;      �q�v�2��J�  |�+���R: �x�      ������D��"b�t @D<hzz��#  ���;      �	����"���8X�  "^q���v� ��a�      �����`08?"�U� �x����� �$w      �u����qvD|�t 0�RJ�W��Qd�      ������`087"n,� L��p���#  ���;      �:[XX��`08'"�V� �\9�5Mc# ��      �XXX��v�}fD|�t 0�RJ?�m�6�� #��      `����<�|nD|�t 0�^�w `�8\       6P]��s~L� |�����  8Z�       ��뿏��"⋥[ �ɓR�$�Jw  w      �MPU�'"��0r 6�C���y�#  ���;      �&1r J�9�)�  p4�      6��; PBJ�}��=�t �]1p      �dUU}bmm��a� l�V���t �]1p      (`׮]�4r 6��~���#  ;      @!F� �&KQ��  �3�       � �)��������  �#�       ��ڵ�qND|�t 0��kkk^q ���;      ���������_*� ���ү\~��?V� ���      �]�v}��j�_+� ���kkk/* p{�      �H���XJ霈��t 0�������SJw  � w      �!��v�n0�_/� ����=��֞U� ��      ������F�7J�  �)��m�Ɔ *�      �!����ќ�q�t 0�<33��  ���      `��u���`p~D��n �Oι[� ���      ������#w `#����Z: �{�      F@UU�9?9"�n ��`0�n  �w      �Q���Z��S"���- ��H)=}qq���  �       #����i�պ0����sR�����  �       #����i����X-� �������*� `�      0��~kD\k�[ ��p���駖�  0p      QUU�9"���- �XxI�   w      �VU��SJs�; ��p�����JG  ���      `�u�ݫr��; ��7~�t 0��      �@]ח����  F�E�^z�=JG  ���      `L�u�D�o��  F�)SSS�+ L.w      �1RU՞��r� `������� �d2p      3UUU�� �Ⱥ���_��� �d2p      3)�������ҵ�[ ���j�^P� �L�       c�i����w��D�u�[ �ѓs�`yy�>�; ��c�      0�fggצ����.� ��-��๥# ��c�      0����nn�ZO��?+� ����8�.� Lw      �1��tMMM=!">R� 9�����S� �,�       `nn�[SSS��?^� �V�� ��b�      0!���:΋�ϕn Fƅ������# ��a�      0Av����V�unD|�t 0����>�t 09�      &L�������"��[ ��Rz~�9��  &��;      ��v��s>?"VJ�  C��~��� �d0p      �Pu]�e��I��- �pK)=�t 0�      &X]���9?#"VK�  �+��KM��P� `��      L����(��܈�n ��o۶��� ��3p       ���SJs�; ���j�..�  �?w       ""���^�s�[� N9�s�[� o�       ܢ��&"�(� �V��~f� `��      p++++��xS� `(]\:  o�       �J�4����gGĻK�  C秖��V: _���v�������=g����"b@J���Hc��	�((iAꚲۈ���")�s~gN;��h��f�	����(%!�>!o �T�HDH-�(�
�Y���9_hл��9���z��׃O.      �G8y���d2yeDܗ� tK��w ���      ����VD\[k�lv ����D۶��; ��d�      �cj�濧��/�R��� tC)��]v��fw  ���      ��5��\k�&"�n :��  `1�      ������^�wMDlg�  ��˛��Oʎ  ��;       �d0|��z,"v�[ �t߷����� `��      p�F����Z#"��- @�� ��1p      ༌F�{j���  W��m���  ��;       �m4����dw  �.[YYyyv �X�      � ��p�� ���z7d7  ���      �RJ����7G��[ ���k677�fw  ���      �ֶ��d29��n R\���smv �8�      �(��x���,"�-� ��Rʱ� `q�      p���־���~����� `�m���� `1�      �/�������#�Lv 0S�����$; X�       ��`�R�q6� ��Z�� `1�      ������#�7�; ����m�C� ��3p      `�5M�Z��ew  3󴕕�fG  ���      ��4�#�]� �l�z�c� ��3p      �@�R����Ɉ��� ���Z��ZKv 0��      80'O�ܛL&���Og�  ��S�N=?; �o�       ��x�5�L���/e�  k:�^��  �7w       �x<��Z��� �@� ��      ���F���z7D��� �������?� �/w       ff0| "^�� ��d2yiv 0��      ���i�o��  F���� `~�      0s��p\J�'� 8/m��Pv 0��      ��RJ��ں)">�� 컧9r䧳# ��d�      @��m���������� `���k� ��d�      @�������5�֯e�  ������ `>�      �j}}����#b'� �7ϻ��;�� �w       �5M�w��#�f�  ����8� �?�       t�h4������ ��1p Λ�;       ��4͛"�=� ��xI��dG  ���      ��(��^�wSD|4� �hϸ�� �w       :e0<<�N)"��� \�g  ���      ��Y__���t���8�� \�R��; p^�      ����O�Z_�� ���Z�m�C� ��0p      ��F�ѽ�����  .�����OdG  ���      �N�F����  .؋� ��a�      @�>|����gw  ��j� �3w       :�[n���ٹ."��� ���j��pv 0�      ����_��od�  ���+++�ώ  惁;    ��)  GIDAT   scmm��_��Iv p�J)/�n  惁;       se8�EDldw  ��� �|0p      `�4M���{�; �s�¶m�� �'�`       `.mmm��ew  ��G�}nv �}�       ̥�m�u����#��- ��N�/�n  ���      ��u�m�}��r,"v�[ ��WJ1p ���;       sm8~��rkv ��j�?��  t��;       so8�="ޑ� <�g�u�]WdG  �f�      �BX]]}}��o�; ��Vk��� ���      X'O�ܻ�KNDė�[ ����  ���      X��z��R�+�|3� xT� ��2p      `���O�Zo��  ���������� ���      X8MӼ;"���  �x�� @w�      �����g�#⯳; �GxAv  �]�       ,��ǏOj��_�n ���; ��      XX��諵��#b'� �6w �1�      ��F��GK)�� ���R�n���� ���      Xx���k��� DD�%+++WgG  �d�      �R���7�R>�� D�R~<� �&w       ��`0x��r""��� ˮ���� ���      X����WG�4� �Y)��� ���      X*������� Xr?Vk-� @��      �t����Xk�@v ,��ӧO_� t��;       K�m�i��UDܟ� ���ٳWg7  �c�      �REĉ���n�e������  t��;       K�i��j�Mv ,)��G0p      `��F��E�{�; `��Z��G0p      `�M&���� X2Wmnn͎  ���      ��7��z�ޫ"b'� �H������ �[�       "��?�Z׳; `��Z���  t��;       ���h���� �eQJ1p ���;       |�~�SDܟ� ��w �{�      �wX[[�zD����� X� �w1p      ���4�}��qv ,�j��Pv ��       �(��yk)��� Xp��=zev ��       �(J)�����g� �"�L&��n  ���       �����#�DD�f� ��*��Hv ��       �8���/"ޘ� �� �6w       x���wEć�; `A�pv  ��       �ڶ��z�_���[ `єR��n  ���       ��`0��Z�k�; `��Z�m��� @7�      �9�F��R�(� L�ȑ#�gG  �`�       �a:��!"�%� I�߿2� �w       8���LD�*"v�[ `Q�Z��n  ���       �S�4���� �(j�Wf7  �`�       �̙3wFć�; `�R��n  ���       .@۶��d�x(� �U� @7�      ���_���fw ��2;  �w       �MӼ/"ޕ� s�m�^� �3p      ��4�L��gw �+Oy�S�� �3p      ��4�����#b�� �joo�� @>w       ����.��-� �U��3p �      `�lmm���� �9e� �      �~i�����_��Iv ̛R��; `�       �i4�}Dܝ� �����  ��;       �Ç�vD�Sv ���w       �w��r�N)�5��� ��j� �      �A�����9� 戁; `�       �̙3wD�ǳ; `N<mss�I� @.w       8 m۞�����- 0��?���  ��;       ��h􏥔;�; `�z���n  r�      ���ں���� �� ���      ���m{6"n���� �^����  ��;       ��p8�t���� �e���w Xr�       0#gΜySD|!� :�� ���;       �H۶߬��5� ���b� K��       fh4}����� �(w Xr�       0c{{{�F�W�; ���`��      ��mll<Mv t��; ,9w       H�4͟�R�*� :�� ���;       $����� �!�� @.w       H�4������ �Y�  r�      @��/��TD|<� :�� ���;       $:~��$"^�� �'�ZKv ���       �5Ms_D�qv t@�ԩS�fG  y�      �vwwo���;  �t:]�n  ��      @lll<Xkm�; ��`��      @G\q�o��Oew @2w Xb�       �Ǐ�L���GD�n�D� ���      �C���?\k}wv d����3p      ��9t��zDlew @�^�w$� �c�       �����R�� ��Pv  ���       :hkk�tD|&� fm:��� �<�       �Am۞-�ܚ� ����|p�%f�       5?Xk��� ��Z��; ,1w       �QD�dG ���R�� @w       ��ht)��� 0C>��3p      ����ݽ#"�� �Y����3p      �������'"ޒ� �PJ�g7  y�      `loo�.�|1� f�w Xb�       0ڶ��t:m�; ��Z�`��/)���564�    IEND�B`�PK
     E"BY$�8��  �  /   images/b96c8ad8-7845-422d-b49f-326b2968fdb8.png�PNG

   IHDR   d   �   ��   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  WIDATx��]	��y�_wϹ��^i���@� 0�q���$Ħʮ�R&�`W�Ul�T%8v�rQ�6�������# � �s��fv����������jzv{v�z�;�=}���g�Ò�!C����AH�� $`h04	�B�!C����AH�� $`h04	�B�!C����AH�� $`h04	�B�!C����AH�Bv�['��G$I�E��vo����6_T{���V�Y���'��1n���]+�L�p٬��J���ˉ��!��8��{�$�}�`�ƶO�LIʁ��;W$����}�*��>��&QȂ��N�cJȮ�����ݻE	��T�RC�/CE��aǁ�%�������>�8	c���΃b�����6�mz�MB�Ν�~��"ᰴ����Ƅ�]��&��WtG���E͞Mu�BNA���
<�A�H<�����Qo�BY�r"Ρ�������S�l�&ټ�%�}�
���%�)!��9G,���(����4���A�%�U�)^��Q����$A$��Aƛ �(���nH�'1P�A&�f���^-�w��2D��H�r��T���������R��|�_R~��s|�Æ�~�	�ļ����ޒ�����R�A�� �|�.4�0�]*�%���y�P�n	�㸫q���������:tZ^]�_	i_�F��+���mߊ]G��zW���4Ř3��]]�N&��C��#�/KȀ��]����|�����--2��$��WE1~ �����W�S�ID��$v�q�*{��\n��\�O�Nw��c�ſ��BZW�>oE��-��鑝r������7|!�%�3�$��C|�Y�$BK- �u:��}���ʕ5u�i}t���۲%�ٴ)��ޝ���{��J�a��z��j�JO��|������'�&�d0�S������r��T�RB����{����Uxժh��c#�͛3��^J����ʲT���
���b�B4�o���D�MJU���x�G��>2~���V� �=�Ւ�g����Q�����	%�Z�,�y�T���n�_���$~s%$���7�?ERv�]+6l���a���d�F��A3�Fe�V��mmV�g�n�TK
T�}��cC5���p�N�_�T$�"g���8"������|H��D"_�6��E'!{�:KlF�^K_�WS���d02��TdݺX���ned�:���}e������t�C%��K����QxLfAR\�c.^�_yesߓO&ac�**%�R���hd7I4�z_-o�!c��"��ߛ�f��fRSl�&���E5�X��3:ᄈ��餡�K*f��q�y3３��ȆV�GN=5[b�J˔)F��˚����Δ\��])����k�:�5!�'gh}�x�� �J�Z[�إ�6���C;�z#��#)�����A�{HCf�ƴ�m[.z��q��54���PH����ɼ�V�y\��$w�������?�Yiy�y+������w��.�i�5B2\2>��f�ԤT�{�vmO��s��:��뇇<1�J�zc^�duTx���ʼk7�TJg?�0[dS��C}�\�m'"{K�NB
�)���#p>���F+4��5]� #[
T�Pg��~ՋH[���:��GM�pNk��~R
/�L�.�����/{]O���L�����-Pa����+2�����N�����)/2PU��a�i3��IF)l[s�Z<�o�����|p�]���R�?���v��[$�ba$�tt��C�#�ɗq��A옾L�\Bz{��O��Ԡc�?r�Y1s�|k��
��Wӧj�4C#����P-�=�x��88?U���ӺH��*#�������%�1c̤�"Bv_|�@����0�.^�|�� �!�+"�� �r��_L��|SYŀT;��;��=�C�ǂ0<�.Ӧ���|�ub� �А����ܥRo�b���ڵ�C��*	�c���e�o���v�� �i�C|��b�~����sRKT���i�ݷ�W�̔ۡa"'�5f�0G�����Ͱ��sU�����0�L��h�1F$�~�K�a�a /�ҷ|�s�L3�bED�dĩ�!uB��aK��K{��#KH���6�U/���
.(�Qpa�%���QM�	d��g#N�C��K�8�\Y���5��Ȅ��^��87|?! ʈ�_n�u8�NЀ���-H-Fc:���bdB�o*fΊ���a.]j�v��y� U��٦7���;Ꝏ�A�۬!�%����Dx��b|<BJa��Z�4侕NB�?�qc�I$�:��l<���5g�Ȏ5���R�ީԱ��,�� ��\#�!���ν�^V���Pm-EL�W���а��e�D��.�=F��U?h?]�{@:r}�uz{�U:��xN��?B���^v�0�HiRa�݅}:��?.�ukV�z��Ji)o�2@^eQ-]t��'��Yg�.H�������o|y��Ǟ!��>Rx���8l�F���3lӤ���aOB���aU�|������ad�W�xCH�+��𵌃�Y����_h=5���f�QB�ǔ;N��5�4v����]D��&RQ�
OH��Qe�U��t��`,�E�a��*�1�u���!C����AH�0�Qe�X pR��K�s�� �:jY�?�)!����dc���I������.ێR���aY	' �R3B
O֑J5oO���1�ԙ�f����C#PA�n�D�۩�܄�Dǽ�ˠ&��%�m[�}}��l�L�Gc-������l����Pwq�[<���"!E7,A���>��DQ"�@��ߏ�#�4�f��Hd�nlJȮlv��\nJp(_	�im��ӱ4�c,I(��!f���ؓ�N�B�J�!4���t.g���(�Q*G2Bؖ��R�;��d2_%��<>d�d�*�uJ����we2��NQ�q�k�C���R2��m����kB��ТG�m2�t)ݶۑN�q�~�W�-!$���6c
\�R2z��n�d��.	)������香,%1Fd$Æ�WOduI+�%�
�:�[<o" l�'D2���]�U��a�/�T̆W��rM�XF��)Ґ�O@FF��"YW���y��7�0R$A�1P�Ok��T2
�B��"�4ா�yd4'A��e�j�� �d̂[�b�}�o�H��Օ���w2����rF��v��{�߷d�h�d�&�>M��"�L�����	D�'!J:�� �1E�\�e%X�/�w�v���}!�G?�x Cl��q�i��6��5K�����@��d�6߳��7G$߻s�ŬYR+TC�w��9M|�4��3�PSV2v�vt��D}VSZ�FSR�8��s28�c���|���?_q{�Q]E:�2�mU|�9�P�ɲ2��~)BBe:l�j�0r(�5@��
�]�#`��pJz.ǽ&��TZ�KtG�UB���dG[�,ڶM������Qԫ�"�a+>�(�Z�;)O��U�a���ǆ����ʓ��C3�����M�c�}��Bэ����aW��Ve7gU���$���<><�t4�����U*��1o�,�q���	A �J����+)��@�5*����cuuɶի�ͧ�GK�rorr@�_$�}���$����Y�>�[!�7���'� ��A��Ⱥ��{���o�|]O��M�*'�D��&(WJ��ڣ�U_uu}���Um�^��*'�Kw��':<�58�g=LE�\�r��i.��	Q�W�Ji���T^;�֟o�켣�si�0�le��u0h������C滴^�>{�2��-~\�2B�Ov�A��y3�q.-��l?�8i}睪.3�8uoe��dC���(���ž���ޫ��②�Ǵz]�#���G��p	؏?��#R0�@��T@�P��J\�S�Mw�ʮ�Ď<��:4�cX��L3e2���-w���ގ��ի��>�{�p8�P�X�,��ϗ�M��T��Z�*&�0dl惮|�)����ⱅ����}>�^B��r.����♧#�@W���;�._	���SY՜�T�K�)��hѓ5.�#�+�m�؝{d�C�3KE*z�1q�8�%��M�$ħA�#|��%������I��z����Qv��i����(NgǛ�f-�-{��-����n<V*!�F��LB�\���dj�/j&��И����TW>�Ri�J��[["���v�K$� �,+$A딻3B�+螞��9s���klG")+��wɈV�ՠ�,.o.�
��ް�ǹ���W]�-��ch�Ɛ�����������G�V���Jq�/'�}{ЂpAU��C#���b�J���q,ٺ��ˎ�D�\��kM5%ׯ��#�H��d2"P�e;���K����bc=�G�Ɂ3YK���*�=��f���ZN�:. pquWW|���C�%�[Ϙ���+��z�s%�ٳ����t4�p�iF݅�Msb�U�;;+%��=�ܔO����,/L��۶I���t��sU�Qy#��Pȩ[R�X�3ཽC�J�[;�Я��v<�z7�ľY�u��@%s�{���fx+�^pW<�^x��:����h4',���P*r9*jH~H2JSGJ���ӝ��Z} ��܆��|�9��k�tv��%�(s�\��I�84�P�W~����
A��zS��+'���1��G�tp �O=�G��r�����	�s�'���w���l�K煙�������m�h�����V��[�TQ7q��ʲޔ�4T�}��:y>�����˹gΔ�9���O��/J�C��Hd�:eΙ��}Sg2�=�P�>,���ľ���5eE����2�{fx�ᰄ.��[��|�omܲ�r�*�;==hԅ{����F��
����X˖I��gtv�F��l��O��I')�ǚ�%�0�Y���D3}$�ݻ��G��ߗxC�\H��2��@�(���Q��3�5L�ȢE^�D,�.��1�a�v.����E~/�_����cP�>��-F%����T�>{��<�H���r�H���O=��d^]�׬Q��+�$�[)��V	�8г�={$��.9�*'��$*_q�K�?���c�!���,\ۂ}����5�g�q���u�ђۼYl%���O���8�*����&x?1<!\e��s��������v�a'HK��3\2/��s��.�����Th�
��9�[I&$�%
�r�i���%w������%N2)*�P�"0^��Q�{s�k��3��]L���Q�K��S)�}�d7m�܇z��^����%�8�
H�\Ɯ���7F�ituݮc1z!����W8��ST\��4X���}Cj葙l�G�E(���*�@0��/�KIq��t:��b�a�Mr2�5w��Y�\?��4�6?��h����	�b�H�O;������3� a#��)=.��lh�^ɴ�I+Tp-0,!� �;P��ԩl����@d�)�h[4'�	���O9ER�>*YcC��h�i�db�L�0d �w�L�+(7��!X��9�]R�1��Sl�+�TI$���0\Ca��]ǵ���c'����n�y�m1F��EБ$EC%DW���45m���	Z�l��\����F�+|�;w�����$Ā��e�Q$?w�T0������W��C�*��j���q?�	_ ��>ށJ��{�
T�V��N�0�.�JT�e����R��_/�����~&�x�}��3�`�K�[H<�+�m�yr(e
�J�9��y,��<��*�X��	 !�҆ћ+\�6�;Ј��Q�3��MM����4��F�
)�5*v{[�2v_p��W�����oy����9�替�}+Z�Q]���HR~�_��������b�6z���@���'W��}Ar[a���C�?�쀻C�񩫯v��ޙݲ�0�߅��bU]a�*u�Q�`�+�ȝ*�N�������G��fF.z�U�=�_.�W]%]���Ad͚�R�>�� ����绪C��-҃���.H�Ǌj0o���	��GF�{�a��)v���}�=9��|�kσ��a��G}��8��D�ZG01jP2�cY�,��A����n@�`�^����hP�P�ּ��
�g�q�L>�������^W��s����.�t��b�7�5+г3����4��=�����9�<r��ٳ{I��d�t�׭����^���\��K"(;@�m0�+�9eL3��c����e&�e���`����|���~��s��{ͭ��w���Ҿl��B����Ά��8���k�˝��ƾ66���������@ʝW\!6*�5�TW��}p��2��N�f�$h6t�Z���#ɤX�ؒm�R��Ê7*�DEK
tϚ% �c�B9�����>��x�p*er�]w�)7�t�H�Ѣ�kU>�0�=T��t�¶�X�V&�%��+M *��-K7m���A3�Bw:���¼��$�ױ���m�ҥk�S�HAhAe��I���K�k3����t��pg#��A G�~`�<Wu�z�y�����<f���)&K�q��/���~�k�WA��z�%��u_��k]yʫ���6괋Ҹ�?/HP���n�q=��w�H�Qx^�w2�cy�������-?�Bc�	)ڄ���9����%I�dF����AH�� $`h04	�B�!C����AH�� $`h04	�B��J��w���c
��Y�yLVB�B9��!H��;!I9<Pe݋�VطW�CJ�RM��(�+��P�R�.Gp e�a��rp���,�t=ޤ�;!\��(�Tq�kA��Z�/X3���;!�O�:B��W8�Z�٦LB~+�DL��*�CR�F�3��x�R����Xa�u���NKR�G��;+�X�R����Y�����Z��?(_Fy�_�%)uMH��7��A9ՇSӞ�G�ʏ��CO��o�Z��	)���x*���1G��,@�.�`�Rki�{BJ�������Y>]�;(��H֒��'�(!���R�GQ���U�o�ˬ�|U�!�u�]5Q_����P.����עp��kě8�&�LB�R^D9W<R�|�=/NAx-?���JL(B�R�D9�7�%��_��?�&?�mO&!D	)���<�r�O���c�򃟤LHB�R:ĳ)�)����*����k�B�������iD����qʧ�3	��	MQB
�������闣�&�
�EJ&<!+����<���t��T��q��_�����&!�7���XZ~&��s��['/�{���LB
(Qa�7�ʏ�<-�5����Z�5�!JH���D7߫�|�O���*oM&k��RR��r��#����� �:���7(�P>u��;ʏ{�Ԅ��+��ʓ��{�Ԣ�V�*i���>��u~�    IEND�B`�PK
     D"BYWC�� � /   images/f1393e3f-31c1-44d6-9d33-bf195c230c11.png�PNG

   IHDR  �  o   .��   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���{���}�������̙�rw%Ҽ��Kʲ쀒)Y!G��V��T���v���j#�l�6M���6+�M�8i���S�M��rk�q�±%�q����ZǼjI.�r��ԮI�6;;s��;�������Cr����<'  4Г9>�#�W�&��[��,�     0�rη��Jwp������ȥ;��c1N)}=缓s~*��LD\J)=_�91"�_�p��v�Z `�J   ����t      ����,�g�[�Rz��{��h�'�xv�����~{�;;;���~��v'S �w         ��7����>��nw{4�˔�"�s�_�x��o�����3Ek��g�        �Q�Fķ眯|R�p8�4�~-">�R������ϟ?�_. �F��  �>O��l�x_����o�J'     L��s�Kgp��*���{8"~%���)�z�/� �3p ��ܙ'�     /��}v�ϝ����9������>��[: (�� �F2pg��    �4��e�>���E���ǿ���>Y: ��        �&uD���믍F�O�;w�M�� ��p�;  ��w��    ^��g��y��s�ğ�ɟ��C=4. �        h����>s������ܼ�c��B�  ���        �$ߚR�����/nnn�uCw �-�         4�ZJ�?����7�����?�U: �v�         4ى��O=��ÿ���� ���;         ��Rz}���F��h4���= ���        0K�+"~}ss�gϞ=�X: �:�         ̚�R:SU�oomm��t pp�         ̤��krο�6w hw         fٕ��766�^: xy�         ̼��k���_G�я�n ^��;         󢎈�9����3g�c �2p        `�|��������-�C ��3p        `ޔR���hto� ���        0��#⟌F�� �e�        �<kE���F?T: x�f        �%������~錩��vK'�Q�#��lmm-|����1 0��       �e|�s��?��?.�1UΜ9�v�t��s����F� PNU:          �D�9_���|�t �+w         �\ιt�a�������åC `�        p�RJ��IJ�S����)� ���         ^��R�̹s��T: 扁;         ����x��666�K� ��0p        ��vsUU�����[�C `�        ��{�#�<��KG �<0p        �W��o/ ���         ^YUU�ϏF���! 0��        �`n���Q: f��;         �G666�. ���         ����>�|�t �"w         �:w=���?R: f��;         \����?���� 0k�        �ꝼt���# `��        ��|�̙3˥# `��        ��,u��3�# `��        �!���F�� 0+�        ��RJק��_� f��;         \���n �Ya�         ��ϟ={��� 0�        �ڤ��>T: f��;         \���J7 �,0p        �kw����m�# ���        ��u��� ���        ���Q� ���         ��=�ϟ���k�R         8��?����# ���        �����7�n �&3p        �#�R��t 4��;         ��� ���        ���V:  ���         �Ϋ�ﾺt 4��;         �֩S�N�� ��2p        ����� �T��   ��H)]������   �ٲ����tǠ�n�N8V9��9?��/�1͗RZ(�  Me�   �R�V�u]_����y_��   ��z����ҥK�38kkk�&���}�y_��8��q�������!|�� ���  `��u�V+��v���+�v     f��O�|�O��9_�_���ݍ���	��J���n ��2p  �)S�ut:�+_/��     ���O�l��?��Ǳ����������P!np�ka�   �����nG�ۍn��vv     �Z]�������Gğ޷��cgg'r΅�K��� pH�   P@J):�N�z��v��R*�    �y��=�|e쾽������f^J�D� h*w   ��v��~?��nTUU:    �9�R��)�9���ގg�y������ �T�   p�RJWn�i���8     夔���E�׋���x�g�駟��x\:mּ�t  4��  �1��:�A���H)��    �穪*�A���ى��z*vvvJg͊7ED�W��U�Y�   p�꺎���8q�D�v     �^�Ӊ���X__�^���k����yG� h"7�  �i�Z����^�t
     J�Պ�������SOťK�J'5VJ�/D��� ��q�;   \���bii�ʭ6     �tu]_y����i��� �&2p  �CJ)���B�8q"��~�     8r�V+VVVbmm-��v霦�{ss�u�# �i�  �:�N������b��J�     ��j�۱��KKKQUfg�R��� �4�i   �U��*���cuu5Z�V�     ��~����>����|�#Y- Mb�   ��vc}}=z�^�     (���XZZ���ը�tδ�Z��Z: ���   ^��[�WVV|�*     |C��q���<������ ��+   /��n��ښ[�    �E��bii)���#�T:gZ-D��* Ma�   /a0�xU     8�^�kkk�j�J�L��������� ��   �MRJ������m3     p@�V˧��������S�; `��  �sTU���^|    �C�|����b�itr��?�5� �2�  �Z�V���G��.�     �������>)���}��G?U: ���;   DD�Ӊ����*��     G�����ʊ��7�9��h4�,� ��w�  �{�n��     p:�N����`�~r4}�t L#�   �k�n�G�    �1j��F�/Ԋ��lmm���! 0m<c   `n�z=�v     ��V�e��Bu��ӣ��J� �4�l  ����vciiɸ     &��j��ʊ�柯������5* ���  ���n���     ��m#��rΟ�F��藎���  �+�?��     PF�Ӊ�pX:c}hoo��Ν;ws� (��  ��QU�[a     `
���XXX(�1��m<�_�[: J1p  `.��bee%�.�     D���bt:����dUU�����g>�я�( �f�  �\X\\�v�]:     x���e�Ӽ���};;;�rss��/� �d�  ���v�1Jg      ߤ��X^^��R�iu*��?�F�ώF�7���I0p  `��u��˥3     ���n�]T�������������J� �q2p  `���     ����b����Ӯ�9�WU��=�����'K�q0p  `f-,,x1     biiɥ53�������wkk���ں�t �V�    8�V+Jg      �j�b0�SO=U:�)z9����p4�rJ�_�����C=4. ���   ̤�p�     h������tFӤ�xw���>}��nnn������]��� �8np  `�����t:�3     ���R����x�'J�4�ZJ���������?N)������~������ 4��;   3���     @3�z�x��cww�tJ���^?�����O�~r4�zD|.���O~�Y� ^��;   3e0DUU�3     �k����=�X�Y��FĽ9�����JJ�RJ_�9!�������ץ# ��  �RUU,,,��      �Q�Ӊv�=���#�T:�H������s�����h4z""~/��Ŕ�Wr�_J)}�����������_��z���O�䥲� �:w   f����̽�     �jaa!��������xkJ�����ߏ�������ۋ�h�dD�术\��R�{1��G"��o����җr������կ~�+=��x�?2 ��  ��PUU����     ��v�Q�u��e�гx��X��H)��/�9Gĳc�ӧO�F�?���I)�����璉~�_>�\ ���  �������    ���K'L���J'0'�A\�x�h��?�vD�."^�s��ˏ�h4�bJ�E��9��g~�g~�d$ ��  �x)��3    ��n�K'L�������~�O>���Kp���ܘs�������b4}1"�I���z��/��O��S��w   ���-    ��$F���7��Ø��RJ����ҥK�܋�1"�JJ�loo?�������C���|��'K�p||�  ������    �B&1:�t:�~F�L��0&�z�^����8z9��[���F�ѧ����Z:
���w   ��k�'   ��ħ;.--�M���|�g�u}�g��v;������"��}�,F��h4�^���I)}�_/��p�;   �V��    ��I�WVV���&���1��4GJ)��n��ZoL)�TD|i4��ٳg��t ��3A   ��    ��$�Ы���~F�L��0p�u:�bg看�́-E�G����h�[[[�-��y&  @c�Z�h�Z�3    ���>�3��n,//�9Mq�u�����J�t:7�s��K9�������g��Z:��g�  @c���    ��B_��9gڵ��8y�䱟c��7��ʥ7\�*�|_]׿����S��G|@��  �X�n�t    PXUUQU�?������&����'�x2�b��v��s����tr���Z�?�F����{��  h��R��   ��1�1�7�0�a���馛&r��;/���'"��ӧO��h4���1 �<Ϻ  h�V�)��    ������Ǎ7�x��L�����[o=�s��f^�7>p�����gϞ],���L  �FrK    pY�ә�9��~�DΙV7�tS�z�c?ǈ��R׵�o8
UJ�L]׿������1 ���;   �d�    \��t&2z��[����9�����DΙĈ�fJ)E]ץ3��TU������ϟ��;� 8w   �>    �eUUMd�Z�u�y��~�4Z[[��o�y"gM�F~�i^�9��	�"E��#�<��F�ѷ���Y�   4Ҽ��    ̤F�w�ygt�݉�5M��L��I�Y�檪2��I�'�����/666��t �   4P]�^�    �gR��N�w�u�DΚkkkq뭷N�n���_^V��;sa���ώF��y��y���'a   ��=    �7��0�۾��biii"gM�����{l'u?�U�{�x17RD��#�<�>���-���W�   4��   �o�R��8��j�;�񎉜U�m���_�����z;�Fιt��}��ۿz���ӥC 摁;   ��w    �������u�7�m��6��J񶷽mb�u�ݨ*s&^�Kp����u�����C �g�   4��   ����&:������X]]��y��R�{�7���Μ�Y4��0a7E�������C 扁;   ���k    �Ť����M�v��~��g�S'��ķ|˷L켔Rt�݉�Gs��AιȹL��������U:`^�  �8�    �K���=�ĉ�=��=�9����5��������~�k�L=#�������K����t�<��g�        ̽N��Vk�g�r�-q�=�L���r�7Ļ�����Dσ��&����R�����[K� �:w        f�����ϼ�;�����G�U�zU����'zn�ۍv�=�3i!���lmm}{��Yf�       �L��z��="��o~s�{�QU͛��|���}��}E��%ސ ��s.��tX�9������J� ̪�=�       ���R����"g�~������Q7��q�����ț��nt:���p�ND�?���?|�t�,2p       `����b7��|����~0N�:U���j�Z��w�3��w{���N���J'0ERJ�i�Z�}����[ f��;        3'�������0����ǝw�9��ؓ'O�������b�N���4JιtS&������~!"��'z�3p       `&���h�Z�ί�:�瞸�������:�����=���������E[�����4ϔ����777�t�,1p       `&��byy����]w]|��w��]���R���nǛ����Ї>4��/,,}��L��z))��l4�[�`Vx�       ���t:����ҥKE;RJ�׽.n�����?�����?��z�����x��w�uW�z�c?� 꺎���� G���x���7?���_*�t�        ̴�����ގ����)�R�׾����׾6}���������?��x��'��V�7�|s�~��q�7FUUG��>
KKKS�pN�u���w�}�|衇ƥc ���       ��VUU,--��?^:�y������;{���_��W����/x����cmm-^��W�7��N�������p�����$p�yի^���_�h�T:   �����+����Q鄩3c0��     �'����~�tƁ�����׿/^������ى�����::�N����������n�t��u�]w]�d�������c�=6�3���#�)%�>�A�VU��O|��Q:����       �\XZZ�2�vu]���j����N92+++���<h�����h4zӅ�K� 4���       0RJ�������at:��pMrΥh�ץ��Z����l       ���j�b8�Θ+�^/Jg LT���mll��t@�       0W�A,..�Θ�v;���#�T:`�:UU}*"�p��       �;��0�A錙V�u���EU�(s뻶���b�����       ������^�t�L��*��׍ہ��s�/x��~��&�       ���R�����t:�SfJJ)��ף���)p�rΥh������� Mb�       �\[]]�n�[:c&\����j�N�c�R*��5(���nll��:�i�       �kUU���Z����)��j�b}}=��v��U�
KUU�����        "���cqq�tF#]����YW�p�ot���ӥ# ���        �ٛ}��a�Ò��6N�Ӊ����*S$��1���-� �Y%        <���b���l���R,,,��_>w��J��i�%        |�^�'N��N�S:e*UU+++���T:�I�{{{gJG L;w        xu]���z���)S��nǉ'���Nh�����{���0p       �����kkkQ�u锢RJ1�ĉs�X VJ��G}��+�0��       �t��8y�d��H)�Ι�n��]w],..�N��rΥ�9�\�`��J        @S,..F�ߏ'�x"���K����b8�`0(�VUU�Z���*RJW~{9�+_������������ڻF�ѷ^�p�J� L#w        �
u]���Zloo�ŋcww�tґ��*c0���0�RJ�n���nG�ӹ2l?J9��Ǳ����۱�����Gz�k��9    IDATK9������F�        p�n7��n���ēO>97�WU���`�s���D�ߏn�{�?����jE�Պ~����q�ҥ��ޞ��{J�#�?��\�`��[�        `�t:�X[[������B�C�Պ���8u�T,..6�� NJ)�뮋�����z�~h�۱��'N�������HǄ�4��\��i�w        8�����8����駟�����Y/�����z�����n�Ü��*��~����+7��~?��~<��3��SO���^���#��KG Lw        8Bu]�`0��`�����3�ĥK�b<�N��ҕQ{��1j���s��s����v����4u��������ťK���ŋ�s.�tdr��E�_����A����	        ��n�p8��'O�ɓ'cuu5�A�Z���2��N'��a���ǩS�bee%��n���ի�:VWWcee�������q�ĉ�v��S�LJ��s���U�`ڸ�        &����:z�^DD���]��Ǳ��{{{�����߿�nG�պ�[Cv �Y������beee�ns��/�� �&�        P@��zћ������u��]�R��UUUTUu]O�h��p���tƑ����j��'���x\:�Z�����# �Isߊ        3���h�Z��t���E�׋�`p���G�׋n��v۸xI)�X^^��q�e�v;���^�Bs��3g�KG Lw         �1)�XYY�^�W:��TU����n�K�\�V��yk��ib�         3����N9v32r[� �ib�         �s.�������b�~��A]ץS%�d���         0#��a�z��WUU���DJ�t�a|����[�# ���;         �4���n��ŴZ�XZZ*�q�Gy�� ���         ���X^^.�Q\��k��?�tg��ia�         ���<շ�O���b�u]:����� ���         ���G��.�15RJ���T:㪸����        ��K'<OUU���X:c�t:��v��3,�|k��ia�         ���Ue
�b��a��Jg��јX���W5         h������ΘZu]G��+�qP�s�Ν.0�        ���A�n(/b0�N8����הn ��         �0)%��@�Պn�[:����         p`9��	��t��L ���N8��҉� ���n         �0no?�n�ۈ7�<k��         ���*:�N��H)E��-�q� ���;         \��s����v���64MC��T: `�        @�4d�=U�5�y��f�         Ґ��T��*Z�V錗�s� �        �1RJQ�u�F���{D���;         4FUU�R*��H��� 7�<��         ���O-�@3�        �U�9;{�o!�f;�f0p        ��H)�Nh,�@3�        @CT���a�4�_�         �!���c��         ��3phw           ���;         \��s� �Y�           Lw           ���;           S��          ��`�          �T0p          `*�        �U�9�N ��d�          �T0p          `*�          0�          �
�           Lw           ���;           S��          ��`�         W)�\: f��;           S��          ��`�          �T0p          `*�          0�          �
�         p�rΥ `&�          0�        ��� G��         !�T: f��;         �����        �!�� ���;           S��         !�\: f��;           S��         �� p��        �RJ� `��        �!�� ���;           S��         !�T: f�����޽��]�w��\����3'QT��Z�AEQK@�kk�{Ҷە�o[-�Z�h�Y�m�JB]�rP�V�]P! 9d�TY�D�E�Z�c23d����� x(`2�������ȃ�\�LfH2���n         ���s� �u�          h�           �w           ڂ�;           m��          ��`�         ��s.�  ���;           m��          ��`�          @[0p        �I�9�N �Y��         &)�T: fw         �$7���2p          �-�          ��          h�           �w           ڂ�;         LRιt �*�           �w         ���R� �U�        `�rΥ `V1p        �Ir�; L/w         �$7���2p        �I2p��e�         ��R*�  ���;           m��          ��`�         ��s.�  �Jw�  ���:w��]���V�[E��������!鈁�        �42p�3�e���r��<��3�iծþ�e�        �J�t  p�v�����         ����Cl>���㪈8�t       �#^ ���; t�����H骈X^�         f��; ���l<,��u��-         0�����w�����<r�|�       ��J' ��a� m*_���o$}."^V�       xb9��	 0k�@ʛ6�G��5�[         �U��.��܈���         �J� �f�l|wD�U�         Z�� ���yό�M�;       ��s.�  ���; ��ݛ�\�s|�t       ppRJ� `�0p�6��܍'�Z�ǈ�*�       7���1p�6P���E�y�;       ���w �>ݥ `�{�~��������޼F���c}cC_�C�W(       �����; Lw ���-�iv-o֚�j�jyUՖ�T-�HK"łZ����ȩ7"Q-�H��4"�"��cQDꎈ����i��_6#"��]�������>        @'0p`vɑN�a���#sw�i)Ǒ�i)Ǒ9���,"-�����X�S��z�SDʑ"=��"GD���?�����         0���_������g�H��"�ɑ��T9������zW�DD���or���)�7G�;R��jF�VOW������)��?��ۻ�}��(�y���kR��3���9��FN/�/����         �w ���[7�T���kG�Z��*�g���9=;R~v�gF���N��Oݬ��;r�t���-�J�t�ē�ˇ��c{#b���;���?˛6�-^rBN�W������`7         ����[���Z��K���9׎���"������zRwD��S����
vZc4">�>~���<]o����"⦜��C��Ĝ��F-�)r̛�s         �<� ̘��S���s��R-��~>r~~D><RD�?����me_��X��x��o��}3yPJ�#��RD|����O{���gEĒ�<       �SΆ 0]���5�k����u��q���^���^9�"�؎=�M�m,G���i�;���ݭ>�)�8���������=��}�w�        ��b��A9��.�/�}a��"E���Ñ�+���'#�Hnd�<߈Z>��?��˥C~8t�O��񣹊�#���M         ���; O����ڳ��+��S���s���d�>k��O�-��<�̋FJ����t�?���{��Ž�o+�        ��3p�1'\����{_�"�"�Z�S:���SďndO�n�S�o^~�E�X:�<k���"�7o�%��("�n        `���a+�O;��&G�����z��>�_��"��}6JQ[����T:�@,?��O����o�T]���        `f��!��x�QQ5^�#N�H�����x�R�l�>�� ��k����;K����9�+��X)]G��      ��s��R� �x� �؋��)U�~壃��l�Ȝ�9lwnƫ;��)2��s�??��?�ܕ��)"�,�        ��2p�E������^Q�.G�ڌXnf�GF"Һ��ޙ��Gq�G����3֦��E���=         Lw����>�����Hq�pʯ�\-.�D[�)�__~օ7����u�Ww�w�o�r�,�,       m %_�t0p�0?}K{T�:��iw[;O G��г.�|��t�Y]>p��͑㿖n      ����; Lw������ګ���)ֻ���t��OKḠ�����+"��-         L��;@�z���?�^�~5��!Gzu��ni�`M��s:�#��!3!�ya}��g�~4���S�        ��1ph#/�q�ӛ���H��FT�I=^���K��=��|�t�L:�mܹ{��-)�K�         05� ���v�SSo����7�U~Q���ڙ&�[���tD+4��������-         L��;@��۰��X�R���C��ȥ��er��~����h�����6���H��-       �M9�Hɥ� 0U� -r�U��[������9M��"qS;3���ꐏ��h��������3"�*�      ��c� ӣV: `VˑVn{�I+��_�x~�����H�8�t�[��7O?g�h�Vz֦���*�        ���`����GU������Hձ�{�s�ԕ?Q:�����xjt�'"�J�      ����*��f4��h4�s�f�UUE�9RJQU�c7D���V�=�Ǯ���������p����* 05� �d����}���)���l��"zJ71W��}�G~P�����������-"��t      <��s����z��F#��洽��RtwwGOOO���F___�j�i{�  0����׿��]]�����"��K'1ǥ�,�PRN�O���     h+1>>Q��#�{l��}�^���������~l�����i  ږ�;�$�޾��7D�3#�WD����.r=�ו�(�QO��t�>/     (��h���h���DUU�[�F���DJ)zzzb���1�|cw  ڊ�;�Axq��<�=�[��?̑�.���G���KG���w������wF��[      �{��f������X����9�+�111��Ï�{{{K� ��;��X��������"zf��`�r��Nh)GN�      �Σ�����DΝ�r�������8�C���ϭ�  c�����}K���9��_V�DN��������/�     0��F�۷/FGGK�L٣�����Ăb�����p:��- ���~��/�~TըޚR>#�8�t���J7��]w�Jg      0�5�ػwo����N�v�z=������E�ży�J' 0�����N���+�-7�g��K��d��t�tC;�nVwջJW      0�ctt4���g�m͍F#������//^�ݦF  �<���U�N[��(��[)�I,�l��?��@�v����زq_D,,�     ��1>>����h4J�����x�޽;.\�rH��J' 0��sS�������o�ȧ�΁i2\:���w      �AUU1<<����S��9�޽{ctt4�.]===���-�=	 ����SVߺ��~�Mi{z{D<�tL�����ވ8�t      ���h���М����4��ŋǂJ�@�1n��3p�G���f���RJǖ�"��nh')���t      ldd$���#g�;���s�ٳ'���b�ҥQ��J' 0����O�ð�Y-G��nh'9��      t�Gܣ���S����x�޽;�-[===�s�-��� Sd��J��t�#�/}�������{IoTSz[c����{��~���?�����3Sz�iQ�       :O�9cbb�tJGh6�100˖-�����9  ����b�N��k��s^S�ԟ��r^�s~�����S~���     ���l6cpp0�F锎���.]���/� @�3pf�o����7����♥{��ި�+r4�a,���u��͋�%�;      ��F#������sٞ={��l�K�@19�H��� 0�@�[ٿ�����"�K�@I)r,J�x8��N)nɲy�檪��      �3LLL���`�K�t��s�ݻ7rαh�\fn2n��3p:֪��/�H��Kb"������      D��0n�f��틔��� �w�㬺��Ϗ*�����t���i"����"r:�t      �*���o߾��j�`���)  tw�c����gֺ����ꍑ�V��ё1�Kg��_*      @{��*��l�N��r�1<<�Z-�͛W: �b����W�]�v�qD�s���JA�:2F�+r4��'J޴�w0���      ���sF��(�2������˗Gooo�  :�����#�޾nC^T�fD~wD�/��;�8<FKg�{ɡ'F��9     �	G�^/�1'�chh(��*� @�p�;ЖVl_��ڍ��rv3�g������w�����s�{      ����h����ΘS������X�|y��<  ���;�V^x��֕��*r�1"��&�Yio|%���ʛ6�洡t      ��hĞ={Jg�I���X�pa�  ڜ�;�^�������8R���1w���i��8:��s�C�K������      ���chh(rΥS����x��??�p�ݻ7&&&��hD�^�Z���������͋�K�Ʋe�bٲe�x����Oj�޽�� �1p�[��W��O|8"=/����1~!�Ɂ{�tV�      ����p4���NUU���o�w����C���>:�>��8�cb޼y�\;uCCCq�GDJs���r�>�`�܁bV^�;�7R~S��m�Hc�4���SZf׹O��W��      ��LLL���H錟�{���������m���q�]w�]w�]]]��g>3�����1��ZmZΘ���bxx8�,YR:fD��J tw��������� G��XT�f���x ]:�ej)��t      �'�{��)����?v�����wg��f���sO�s�=�hѢX�bEw�q��]~.4::,�����)0��� SW�W����j��W��ۈ���-0�=-��3���^>�tʌ۽�����Jw      �~FGG��h�Έ]�v�M7�����޻wo�t�M�cǎ8����~�n�9���c�����  �;�@K���ãY��;�w��"'����齥;f��7�=?��-�;      h?UU���pц�����W�w�qG䜋����D|�߈�N:)�<��b-166���/� 3���9 ����[�}݆��pD:�t�5S#^ѽ��3i~ڿ)"�U�     ���w�ޢc���/����ؿ��ǳk׮��g?<y��    IDAT/y�Kb����nQ�y��ŝY��3 L]�t 0{����G��_�������P�3ҾW�w�Kw̄]�n<9E���      ��f�###�ο�;b�֭m7nT�9n��غuk��SUUE�`&�� ����~9��m����߈�ח΁9/G��?����SK�L��{󑵮�TDt�n     ����7�͸��k㦛n����4�{�7.���(r��}�� �	���z��k��j��kS��K9���sD��}�}l\P:d:�w����uY�xJ�      �O�����z\u�Uq��w���ؿ\v�e����쪪btt��� о܁�iSmն�6vW�;"���9��Hqb�H\�7m�.�2��]�F�"痖n     �=���^��֭[�{��^Kϝ.cccq����� �g�L�n\��Ukn돔/����{�'��CK��X�xCW��ț6u�`��s�i�[      hO%no6�q��Wǃ>��s�[�^�+��2[zn�ٌ�����	 @�2p�d����]���T�809�M�.����Ϟ_��`���opɽ�N)�X�     ��566UU���n�!�����̙266W\qE�۷��玌���<  ڗ�;0)'\���U��/O)�.��'E�]�F�0��?8�tˁ�����c7D��X�     �����������w���3gھ}��k�i�&&&Z��  ړ�;p�Vo_��ޕ�9"֖n�N�{��7j��k{��p�Oϯ������W����{�[^RF���n     ��5��o�y=�P�|��-;��|����[Zz���hK� �=�lE�iKWm[��9��#�#n}�v7�;>t�9�\S��(�pt����3�[޴��P���l�ٽe㟤T})"�)�     @�k�@��h����h6�-;��v����{o��3p  ��8@/ھ�յ�wF�7�n�]w����K����-g�Z:&"bp�_98;R�_DD[�     h_�H�z�1<<ܲ�J���[6����h4Zr̤�s� �hc��Zӿ�{8��iU�wE��垗"]������\��ag䛭�|��һr�""��|      :W��l�8����o��%g�644��~{�^��%獍��[r  ���xB+o8��é����D3S�3R��[��ؼ����>��2Ӈ���F����8-��      �0>>޲����/��V�v�cǎ8��b���3~���Č� @{3p�����1E�ȱ�tPD-R�Z����l�f����f��eo��M�C[�rL3W��j������v     ��Z5p��~��-9�]�����׾/}�Kg������9GJn�s���1p~�˾�a����{S���n���S������r`�ƻ#b[�y{�����y�No��?�+���o�l��R�9�qJձ)ED���       �[ιe7�z뭑��{���_�z�\�2���f��z����3~��v �w�1�oX�jbb��)�sK� m�9�ҙ�����-��"��/"�DĒ�X�"�����3#����5���r      3��lFUU3~ξ}��������ӎ&&&��;+W��Y����  s��;+��������1�t�Q�R���#�      ��V����o}kN�����%�V�x О�a�{ٗ7���(r���-       0�z�%��u�]-9�]��ݻ����sZ��	3%�)�� бj��r^�m����'n1n      ���b=00���3~N����g���s4�?f�q; L��;�Q���;�J閈���-@D��x�      �D�C��?��3:A���f�%�  �~�K �u�U��[��ws��/�[`VJ19�1)��W\Ҿ��WG��8���9��̱H��Z�
      �@UU�s��s��k׮����=��h��0Sr�nq�)0p�9d�uk����>9��t��fDE����P�1�rʵ49�r΃���R�}UNCQ剔j�kQ����V=��k���'^2:��CϹ�݃�9�s~�4}�      `�k�M���w_K�iw9�����c���s�� 0w���j��WV9.I��,�-4Cq_D�?R��v�/j����}�Q�ۗW=�6U�c#"��u���;3��     ���b�w�ޘ����s:�����;<	�������j�i#�����-0��#�{#�{"�{rN��R�'r���f����)�/��҃����7��fDz�      hwU5�wY=���3~F'i�����N�s6r�)0p�YlM��yñ�E��+�SP��{"��qW-򿤪��fOϿ��K��*7S=��l9������     �'Њ����Ќ��IZ���� �2 `V2p�Y�7��i{R��R���n�T��wFNw�w�w�\}3��/��^:��CϾ`���3Gr�F�      �Z1p߿����IZ��p�; ��e��Ћ��{y��%���-�R�_O)�s�qgD׎޾�7�x�h�v����8�f�t~D�J�      �\T���;�����D�hk^�  ���f�����\��p��-��b$r��7G�����~���Y��г.�h�3����0r     ��Њ!�A�O2��'��i��0p�Yb����9|��w�'�R���RT_��ڱgd������KGu�CϺࣃ[�ɑ�>��      -�h4J'���s4���.sΑs6�#�� ��@f���ӺEߩ�*"��tsL�*j�ȩ?El�O�/��K*�5[-?��O��&�O���     �e�U��V�O�� �&�8�p/�?���F�5"�*����=q}��>"��Xs���Isɡg]���XE�����=         0�ܡ������En^9�,�¬vo��:"�]�7��K��*4�zօ��w�h��gRD_�         �.�СVm;����G���-�:͈�="}>r\����vF
���f��u��wo>��S�w�n�Rj���        ��e��&GZ�}ݟE�wGD*���#��+"�kz�Ư��W�.���v�9l����;��}g��}        ���;t�5�k��o\�ሴ�t�@����"�Kb���'oo�N       �rΑ��+`2ܡC߿a�p�_9��t,�{r���r�']��H��c       �if� �g�`�랚b������-t���[9�O�r��'_~W�       ���� 0y���^�m�񩖮��(�BG��?�r�'��         t
whc�nX{J��g#���-t��9�K�R��z�o�%o��Y:	         �`�C�Zٿ�7"�����[hk9"�)��Hm_���k�����p       �\�s��R� �H�ІV����������n�m=�S\\K�'m�z�        ~ĸ &�����m���
����kF�S�>���r�.��         �N��&6\����'>�#�R����'����Ӗ�O����1        <���[�`�ܡ���1�����[h)�����J���ܹ����=        �v �<w(������g#�_.�B[hF�s���y���K�          ���;���a9&���K�P���񑮮��Փ.�~�        &/��w �$w(���Y�t]D�b�Jʻ"j�7������%��k        �:�v �<w(`�uk�Q�]��S��BR�'��`o_߅7�x�h�        ���`�ܡ�V�����\�>r~F���zJ��wl_��ش�*       ��3n��3p�Zu����>r<�t��"����������K�pI3���I        �7����C���v�ꨪk"��-�Σ��������A          m��Z�E�ֽ���"���-��7rN�v~qť�iSe�       0w�� &��f؊֟X��:r,*�BK|?r�������K�pI3��=        �X��� &��fЊ֟X��5��s�@�x����7�O�>��t         @2p�b�>g�O�F�_�|�%{J�          t2w�/ڶ��U��ø}6kF�Gz��ݷ�z���c        h9��	 б�a���a����^ε�o;�ү�       ����J' @�2p�i���'ֺ�����R���*�u�)[��t
        ��� 0y�0M~lܾ�t�nD�����{���}�t         �le����}�����񎯞|��c          f;w����_���q����n]s�u�K          �
w���ۯ1n�UF#�_���շ����1        t��s��Jg @�1p�I2n���竨����/�n�        :�q; L��;L�q��s���;O��s�C          �2w8H�oX�*�����Y�����9_�C�C        �=r�nq�I0p������=��jW��%�[��KUڸ�U�][:         �G�J@�x��^���KG�naJr�|�������          ���p V�����消xf�� �{"���\s�M�S        ��RJ� �#��~���-���ql�� �'�wǊ�k��       0�rΥ �#�����+�.�">"V�narră����N����-          <97��8���ya�s)��[���ZT�`�         ����cM����4qI�xM�&eON��۹�O�         ����~Z�4��\9֕Na2�WS�V�f�         �q�᧬ھns��O�;8h9��`Zt��w��         ��u��v���_E�Y�;889����wo;y�J�          0ynp�Zٿ��)��/���ʟ���_�y�q;         @�s�;D���uoIU���҈��d��[�)r�          ����9o�u�R�ED*��J�P��۷�r���S        ���#%�$ 8X��i��׾4R�t��*��7�Z�o�����_�         ��U+ ���~�q9ծ�J�p@rN����)��a�       @�s{; L�ܙ�^���)��D��[8 ��߸��˯,        "�l� �`�Μs�U�]\���#��K���ʩvڎ�.�f�          fV�t ���o����lDza�ȕQ�}�N�v        :���`rܙ;6m��^�dD�Z:��)����q���dO�        8XUU�N ���]: Ze�I;ύHJw�3���c��K#��n       �Iq�; L��;sª���9�U����;��n;u띥C          h�Z� �i+����Q�����gH���D�D�v         �����Ym��u'���w$��,����yϫ�xͥ�n         ����0SV߸�s�FD_��P�H��q��M�C          (���YiE�i��*_KJ����U�z��\��t        L��s� �H��:��۰$��+#�SJ����OU���_u���!          ��Z� �N�������������I&i����w���$)��Τ-H!��6���(��c�U�\o�^��z)zy��(��b�L����X�$�z�R��ʍ�����9�����Ė�M����s~���1�>
4�WL=9�>��ֻ�8P�7o��-��cH�r���)�v          ���;=���⯦�ח��1��H��5����J�          �y��C�ޜRzS�ӟn�ǯ�����!          t&wz����ߖr�|�]N�Cw�jrtr�t        ���s� �:���lܽ5R~G��F'�)�G�����[        `M��J' @�1p��}��Ksj�/E�S��GhE�7N����!        PB��� N��;]�[><�i����n�fsJ{�쿣t        �b� ��Q: ��ޛ���7�]���-<�Ѫ���       Pw9��	 �u��NW��EN�,���H����[�=��)        P����9����ub�G��/���J�����1n       �'���0p��O�ye����;x����jd�����t          �����141�-R�'�W������ݸ��K�?_:         ��f�NW���/nD�-rl,��C��/]���n{�t	          �����7212����r��J��0��������!          �w:[�4[~?"^P:��y�����?=z�L�          z��;m�Į���o/������8~�go�c�t          �����5|p����<̟o��{&G'J�          �{�K���rb���Ç0:�q;          ��x���}↋��#��-�b�         ��3p���L��cඈ���-�b�         ��0p��L��ߍ�o.��)��          �w:��ɱ�H�-��)�7n         `-���&w�<�������o�㻍�         XK�7t�����-D�q;          ��S���>%�şE�ͥ[���?7n       �S�K'��n��N`�N1[�~�@�����n!"R:�9��1n       �Su�`<�T: ���;�T�_�����D���_9�        VP����S�����J)��tq��º�����(        ����Np��g�Κ���^��tq_��{�G���#�C  �ttۛ�     �ʨ��t�i�3 8}�������$��-�c}��Z���O���J�  ���f0     �S�ܝ� ��	����4��9.)�B<����O^s�ߗ �3a�     ��n�K'�?� ��g�Κ9���="o/�Q{)�#�o=|݁�U:  �T���     �?# ���_:�z>��G#��(�A��v�y��S�C  �lx�     ��j�N  V��Yu�&Ǯ���t�L9�=|��K�  ���Ǐ     g��nGιtFq���s� ���;���w�yN����W�������+  +��     P?�xz{�9RJ+�krf�;��`�Ϊ���m��n���J��\���th���� ���w     ��f�Y:ጬ���H�̹w ����ձo_c���8G<�tJ���C#�[:  VZ7��     ��n�����J't-��;��*�^s�OG����_942���  ���     ��s������3��twV�։ݻs�/�Q{)�|���T:  V�7�    �>��f�KgtO�=s�@w0pgEߵ�_���tK�廦����y�  =��jy#     jbqq�tBǨ���Hΐ����;+����IQU�cs閚��������� ���s�����     �0p8O�=3�@w0pge���h��qD<�tJ�����qç�~���-  ���     ���lv��۫qںC�N_�ٌ��Jg ��C�%"��tG��F���k|�t  �o�    @�[XX(�pVRJ+�k���sz;@�0p��1r���5����ʩk|�t  ��v���H     �a9����	�N#?}��=�9+C�<?R�ÈX���<9���k�Fo�p�  (a~~�t     �J�~Ƚ'�Gt���k��*��tw���|�ץF�ֈ8�tK��F���;��i�  (eqqqUN>     ʛ��+�p�V��Z>�
���sF�޼�oq�һ"��J��Y����G��Z�  (��*'�     @j6��l6Kg���:���j���Y� ����3rߓ��/+�Qs05���JG  @'�$     ������	 d�    IDAT�=zb�n�Kg p�9m�c��?X����]�_^���bu�_  ]��l���R�     `��Z�X\\,��"r^�����b�Z�U��{���\� NS� �˕����۬���i���|�U�X� �D����1P����s���5;;�֭+�     ������	]cvv6�l�R:�#-..F��,��i2pgٮ�s���n�96�n��"�ا�~���! ���>�s�?]��Ӵ[�W��C,--��Ғ�;     t�f��3�������ذa���|��s�8q�t g�Q:����74����g�n����c�F�?[:  :��\     ��%��'NDιtFG����v�]:�3`�β�_��S�H��)����C  ��5��XXX(�     �����h6��3�N�Պ������ �n�<�����3"�]�:K�yjǁw��  �n��     �NUUyZ�Y����ဈ�9�����t1w����oN)~�tG��������t  to~    @w������Jgt��s?~����ĉ�� ]���Ǵ}↋R4n����[j+�X�}�3  �����y�     ����B,..���z�v;�?^������c~~�t g���G���7�c����-5��6�Z�?��[�J�  @7��I     ��v;���Kg􌥥�Z�����8q�D� V��;�*�|��#���5�`D�����w�t  t�V�333�3     �Ǒs����eaa�Vc便%�G =���G����鍥;jl��b����gK�  @���������     �c����f�Y:�'����≷KKKq�ر����wf���oI)�j���]�\{�#�C  �W�8q"Z�V�     �k������\�UWrx=??��'������ wN���/���ȱ�tK}�>4z�OJW  @/��*�;UU�N     ���lƉ'Jg����b=z4��v��s�'N��z�:2p'""F&F���?r\R���R�����ϔ�  �^�n�{�t     �&�V�V�n��J'D�ٌ|0J���v�G����� ue�NDDLǖ�L9�*�QcS�D�u���� ����%'�     @a��ZN�9�?���]{�����ȑ#�l6K� ���KP�������U��ƾ�׈=��y�� �*�����Rlڴ�t
     �NUUq���h�ۥSjm~~>�sΉ6t�	�O��lƉ'�j�����6"��tG�-DT{>q��+  u177)�8��sK�     @m���Z��)k.��q#��ĉ1777n�ء{�ٌ���X\\,��2p��+'vC����}PJ���ǡ����t  ����lD��;     ��:��;]��>5t߰aCF___Ѧ�s,..���|,--m���z���s�4O.�Rc?ht��KG  @]���F�96m�T:     zV�ݎ�G�F��.���h��133333�nݺ�u�֭��=�KKK������QU՚\��d�^G9�����E��Sjl����~*�@�  �������*6o�ܑ��    �n�l6�رc��]fii����}}}�nݺ���������;��{UU�n���jE�Պf��V+r�+�@0p�����o��{Kw�W���X��ط�+w  � QUUlٲ%�F�     �	1==m��Շ��혟���R:��\9gv `Y�kf����9矌�}����k����n�)  �����8r�H�w�y����     p6fggcf�<検sW��M�ه X5���������;"����f΍�>qݟ�]�  ����v9r$J�     @W��*�;f� �C皸��=�Gn�7rl.�RW)����  �c�9����=2     NS�ٌ#G����b� �����ޛ�����wFN��n��_�G�  `y����ȑ#�j�J�     @Ǜ����G�F��.� ���������o�;�*G��-q��Jw   ���jő#G�sΉ�7FJ�t     t�v�Ǐ�f�Y: �!�=nxr�wG���tG�}����7�WO:�  �P�9fffbqq16m���     ���s������l�K�t<� N��{���^9~�tG��4���SW��h�  ��4��8r�Hlܸ1�9�h4��     ��f�����j9�q�<% N��{��������m�c}閚�9������!  �ʙ������8��scpp��     �FUUq�ĉXXX(� �8�����禴49.(�RW)������  �ʫ�*���cvv���     zUUU177sss�s.�ӕ�7 8=�f߾�`��Μ��)5v��5��t  ����v?~<����sΉ��=@    �ޑs>5l���t P#�=f��?�#v���_��H�c�  P�f3�;������)��Y     pFN��>??o� a��C�&w�.�����H��v~�;�K�   k��j���ǣ��/6l�6l�F�Q:     ���j���|���G��v �1p��wo���tG��Sί����}�C  ����v������l�_�>6l��֭+�     ��s���Ř�������9=-��	� �L�=`�/�.��DĆ�-u�r��Ԏ�?/�  t��s,,,���B4�Sc�����i     �\��:�v��.�S�� �|�]�ٻaq��?"?�tK]�85z�m�;  ��UUթǺ������`�_�>����    ���j�bqq1��j�� xL~���r��ɥ?���Sj�c���X:  ��V+fffbff&���bݺu���F�<     zD�9��f,..��⢓���a��ŶN�����Jw��[�w�go�c�t  Н������#"N������    X��s�Z�XZZ����h6��s.� p�ܻ����kr�/�Q[)��v|�'�����)  @�h6��l6cvv6""�FD������@����    ���c��_�f3Z��A{�9GJ�t t�.�ubϋsTo��xJ������)�  ����N=:��F�}}}��j4��     �n9稪*���v�}ꏭV�ԟ� �����l���.kG�ֈ��tK]��ߚڱ�wJw   �t��f�1�7�F#RJ��'�    Г���J'�J�;V:a՝��O}� ug��E��s�������SJ���G��/�@�  ��SUU�    X3����O��n� X>�-�ϻy�V_uK���-5����7}��;��	          V��{7ȑ�?y�G�h�[hTi�ᗎ�t        �]<m ����l���3��u�;�,G��w_���;          ���w���ݯΑ�tG���vxt��Kw          @��/�c���KRο�tK]������.�          u`�ޡ�N��W9���X_���R�c{�q�_u�R�          ��F� i���'�h�O*�RcUT7}�e��s�        ���K' @�0p�0[o߹���g�n����{Fn�D�
        ����J' @�0p� {o�ۗ�m�3"��tK���~����;Kw          @��w������tJ�}`S>���          PG���������)}O鎚��ܷ�Փ/�l�         �:2p� �w�1R���579}������!          PW�O��9�?�;j.�ȯ?���T�          ��F�:�������A��r�/w�          �;�B����ܜ�K��Y������(�          89�����OM}qG����-5��5����j�t        лrΑR*� ]�	�kl�_������g���[jn���S��?P:          �
�5��ݐ��n�W�n��9}�ݣ��[:          ��kddb�qi��qu�����s�        �RJ� �k���}��ӖwD���)���k�JW           �d��r��k�F���S�Ϥ���ƾ}U�          ���W��Į_���-�Q{)����3u�-�K�           ���}��H�#�;j/Gը�Շ���oJ�         ��s.�  ]��t@�����'Kw�R����V�          x|Np_[�����˥;����=�K�+          �'f�&w�.G�ZD��-��4���t          �<��z���=���E����rė��7�ɝ�J�           �c��B�M�]9�G��@'hF�_���[�/          ,���
�:96Z�t "֗n!"Gz��k�?X�          8=�gi���krN���t9����{�          �����჻^�RuGD�[�������?����          ��1p?C[��"R�'�w���)�?��[�J�           g��t@7�vp�U��D�`�""b&�k��(          �9��4<��UT��[��U���C׌�t
          pv����ɱ�խa��Aҏ�1>^�          8{��4|p��rN��-|U�?:�c�/��           V���2M�}{����_��S>:����         O$�\: ����:8����q{'I���7ܱX:          X9�c���7�H��}� �UN�>v���J�         ,GJ�t t���04���9��0n�(9rz�=���)          ����'G�����åS�9~�Ў�7��         89�H)Eιt
 t<���{�޾��j�ND~}��V������R�        �L�����?�w�}�K9v�n��r�������+<        �+�<� x|�q��^��ťqu��U�}�G_t�|�        �3e� �S���w�|F��g�J�����ο����T:          X}��o�k�幊;"⩥[�9���k�v�*�          ��F�R�&v]�s|8��;RJ���F��/�          ��Z܇&vO���ȱ�t�&��������           �V��9����})�����9<�|��8���+          ���_:`�\�����?��yw�ӽ���Փ�O�J�         ���s��Jg @ǫ��}�/�.I�@Dl+��cH���7|��[��N        Xi�� �<=?p�ۖR:9.)��c:Q��C#�?W:          (�Q:`5M�~uJ�.�����9�������          �����޼���s9�7�n��8�c|�t          P^�ܯ�s����-�;"�+���K)���ȁ_/�          t�F逕4tp���}�'¸�쟚��GJG           ��g�C�^�R����-<��4S�&��J�         ���s� �
��������t��H��-,C�7��;?�����)          @g��������T�W�na9�ۭ����/�.       X�����ج
� ���(p����}}�Td��.1�#n���n�ߥC       �ޑs^�k��5�I��Jg  У����M����㍥[X�f�����K�        �%���#w��[�n]��J> ��U�+'wn�o6�8"?�t˖S�7L��       �3188X:���  ��F�eɑ�N���F4>l��]RďN����t       ��:��J't���j?m zEǟ�>�/���䈑���.�ejt��JW        ��'=�I�:��;  ���Op�:9�75ڇS�H�Nۻ�5��JG        �-����زeK4=�YS�  ���<�}���c�wr���[8#��K���U�C        �V___<�)O�/}�K�S:��_���X�.  Й:['������#�ۻԧ�H7~��;K�        ���=�i�:¦M�b˖-�~w ���ܯ����ȿ�s�zyڝR��G_���yɭ�J�        ���>��155U:�8C  V[����H�t��s)�ʑ��p�H9�������!        +�K.����XXX(�R�3���	  ��Fɋ߹���q��ҏ�w��9����1���)       @���V�}}}�g=kկ����Oz�  z\�Q���ض��E���>+(�\D�����ݥS        V�7~�7ƽ��[:��g?����׷��Y�,  й�t�>|�������|SD�J�ۥXʑn:<��C�S       ��J)E�yկs�Eœ���x��V�Z��y�{ޚ\�� ��kq��;Ǯ��}s��{"�ވ�*���S���G�       ���u���	E\v�eq����  �V�����m)�-��}b{{�.��J�95:~K�       ���;����|f|��}]9rdկ�I�:� `��	�'OlO�>�^��`7n�29R|�Ԏ�*       ��RJ���tƚz�3�\p��\+%[" ��[��rb�+�r2;='�7���        �V'�GD\v�eq饗�?��?���J����kv=w  Vd�>|�������|S�ɑ����*�X����G��Z�       �Ѭ���ꫯ���?����\���۷ǹ�[: �9������~r�n�������        �e-�[�l���E�}hM�W^�����zNo  ��g}b�c��3���C#�?X:       ��\q����>���)+npp0^���E��(� @͜����ɝ�9��Y��N���G���J�        <��<�="btt4|��8v�ؚ]s�����믏M�6��u���}��2,�#��w�]1<���Fn|�+�vj�����c߾�t       �r��xt����s��ظq�^w5����ӟ��5���/u�� ��q�WN��><��ї�:"����������'G'[�C        :��͛cll,֯__:嬽�/��>���3�'���% ��=��}�����ˉ��5n�������WݲT�       �t�8%���Ϗ�;w�����_{�\u�U�m۶"�v�5u�� ����2tp��S�?Q�Nk���oޔ�_3�퀓�      ���R*rR�^7�tS�~��q���5���J)�K^���o��"�o4��N�99g#w X����+'wno��["*���ۻ7���M�N�       ]���}˖-�gϞx���_������kpp0����K�\�ؗ:�� ������Fn|<"��k,�x�3�����       @/(9$=�sb���q�UWu����.��{��G�R/%>t ݨ?�k/E~����7޷�*�       �R�FTU�9D�ш�۷��_w�uW;v�Hǣ��[����p4�b��ԍ�y X�����w�>8�}a�       ���R�S�����ū_����{��ꯢ�lk����o�����c���E;"�} xt���ۇF�)v��       �'��G|�4�+��"���gǽ����sO,--�i��_۷o�����_��>��'�C)9g� �e0p����o�w�¸       �i�0r��ذaCl߾=.�����{�3��L;vlծ�nݺ������/�.�`ծs�|�+�� �<�5�#���;��t       �Z蔁�I����m۶ضm[|�_���ۿ��}�sq�������ԧ�3���x�3����72򥮜� ��y�`Y])����7��        XK�F#��*��]tQ\t�E177��<���q�ر8z�h���D��|�_�h4b�ƍq�y��y�Ozғ�K.���?��������?�J��    IDAT ,��{��?sxd�-�;        J贓ܿ�ƍ�9�yΣ�w����l6���?���o���^J���Zs�; ,��{=�H�͇G��Z:       �����N�?��������Kg g�� ������s��=<r��C        J��S�{����	� �\�m1����;��i�       �N�h4�����a� ��0p�]39b����,       �i��6�� 8]�(�?�v��C��~�t
       @':9�v���1n���� ,O�t ++E�}��/�2n       xB��ǽ���� X������å�d�j_}�5����)        ��)㫣���Y  �t�+ɓ��0t���s`n�꿾���T:       ����,�v  �Fo�����/r�w�M���.�       ЍRJ��g�= `%���줈_84���"9�       �l5����tF�q
>  +���{�s�ht��J�        ���C휝7���  �$��4�x�����[:       �פ�"�|�<�F�Q: �c��eR���H;����-        ����)����pMg2n `5x��]������3�߸       `����)%�v8� ��f�H��������u�_*�       P''݆�_����� �����	��S׌�X��>       �BN��sε;�ى�  ��N�b.���S;��\:       ��x�)�u�� ���;��r�7�q���!        <�ɑ{J)��*\��N�V  k��+;Q�������       t�F��3c�RO��  �}�;Mʿ�ν�O��.�       ���w�8ܰ �N�_:�S"қ����!        ���R��"�9��9��d+  t
�N���J7ڱ�t
 @�H�J7�Zy����tBG���<+Z-$    :�C��UU���nz� �������V~�Ǯ;��!  ݤ��Ҿ��F^���N�(o�wa=��t    �ii4�rp�C�k��:G�� @�p�]9��Ӈ�z�Ǯ7n       ��F�񰯓��?��<��п��~]�<�,��8�����F���=r�/#���       ��g�ރ�,�����JB�0"�5\s11�/��b;�$N�6i{&mq�I�t�3N�Ȕ��	v�IhgB�L���L�C��!�`0�`Y`�΂��  ����=O�2�Ү��<������hG��y:��h��y�؋���aE�0�� �#p�z{Y6�+_��Ono�        ���b�eff�?��?���\{�E}�3��7�M �Vk��KM?%�w��+���=7ε�        ��8��cٷo��[�n}�|�����u��)��܇�&Of�����?���[�        `�� �#p��'3��nG�!         ��w ����,��i��7�QJ��          ��;p�I𯾔�W���x�M�.��          ,M�4��q{M�u��粻��           2�'�/��m��W��ӷ��        @��ZS���
 K��}Q�g����}o���K         �&q; ����쨵��=���M��         �m���Z[� �N�h=`t�WZ��w�$n        ���� plNp_�Z�e����/����[         �����Oϛ���y]{��e/{ـ��Zkfgg���s���LOO������b.�������[�����Sϴ�         ,˗/ϩ��:�kW�^�SN9e�� �����ˮ]�����~����ZV˻7\��m=          �k&&&�z��^�:��SO=��{�.�q�m	�I�Ӈ���q;          ���X�"�sN�=��LN.�Lv'���]�/������k=          `Ԭ^�:+W�̶m�r���y}����^j�O6^��wR�o=          `T�X�"�~���o}+333Ǽ~b�F��Z�oʊ�6�c��        ��j��' @���9���w퀷���jɟN֙������h=          `�9�䓳f͚�ڵ�׍s��B�~��        ��*���  M�q����$�������l= ��s��<\�K[� �o����       ��r�ʬZ�*���/y�8�/��~�� F]����        `��|��c�;�          �&'���/��݉�           RJ9�Ǘb��B�~��          `T,��}I�8���ݗ���z           ��Nl��           �j���5��D�qb;          ����݉� @��Z˵�^���z�]����5k���        t�(�/��������?�l�ʕ�mP��w�#p      }�֔RZ� �N��}M>:��G�|���c         �x���غ��pb�Nl          X��;�          `	���G�x�w'�        �d�ZSJi= ����9�ǻ�﫵|t�����          ����-��jɟ����{ו�y��         8��0�{�:t�״���Z>��_>�+?�L��          0d�<s�||����          �Ю]����c^7��݉�           c���ٱcǼ�d�.l          c����c�=�Z뼮D྿��ي���w]��'��         0rj�)��� C����s���ܹsA����������ى?pb;         |/q; ���g�޽y��333���_��}OJ�X�          0~��~�������޽;sss��X'�o��u�+�d�Oݸ�         `�=��sy��G�u�g��5k�x�����fnn.3339x��=�B�C%����g/+{?��+�0�hK         `	�����zu���<������.8�ӑ��X�{M���~��|�PY�7�+n�?�a           ���$�w��I�^�ă�Z:�Њ����m�         �����M�}�g.k=           &Z           �D�         CQkm= :O�          @'�          ��;         A)�� �<�;           � p          ��         0��� ���           t��          �N�        ��RZO ���          �	w         �Zk�	 �yw           :A�         CPJi= :O�          @'�        `j��' @�	�          ��;           � p          ��         0��� ���           t��          �N�        ��Z[O ���        ��RZO ���          �	w           :A�          @'�        `j��' @�	�          ��;           � p        �!(���  �'p          ��         0��� ���           t��         ����z t��          �N�          �	w         �Zk�	 �yw           :A�         CPJi= :O�          @'�          ��;         A��� �<�;           � p          ��           t��         ����z t��          �N�        ��Z[O ���          �	w         �RJ�	 �yw           :a��          �q777�����۷gzzz�� ���R�         0�֔RZϠ���~><�k��ٓ~�?�E M���         `���؜� p���暹k���?��O;m煃zl        �.� ��RJM�����}o~kP�        �%�           @"p          �#�         0��� ���           t��         ����z t��          �N�l=   �G��䄗k�Xr�	       ,]w  F�)?��h�h�U�2=}R�      VkMq� ��         ��SO=u�y���|�=��ӧV�Z�Л ���2'p        �!pz;Gs�)�|��;����w �6�z            $w           :B�          @'�          ��;           � p          ��           t��          �N�          �	w         �Zk�	 �yw         �RJ�	 �yw           :A�          @'�          ��;           � p          ��           t��        FL���  ���        `\�ZSJI��{�?��>��Rʋ�  �F�        C��1�w��G�_�	�/����� �Q!p `$MLd[��[�a���W���)���n=    `�^,\_hľ�u�;  ]'p `$����ʸ��Ƌ[O     `�������*�� ��;        ,�Zk���c��Bw  �@�        �`���#�lv�;  ] p       ��p$�����,����|?��L�         ��H�������|  t��        �����q r `�&[        �Qp���qt$r/����x��q�� %p       ��8��S_xD�p�o `~�        p�����χ`��� ��;        ��Z� �%��a�|� ���       ������v�9� �X&Z        ���/��� XLNp       ��O������|��q�;        cO�~�<�pt^  �#p       `�	��� �%p       `l	�_�5�~��  F��       ��$n,�-  �C�       �X`�  p<�        ��~��z�X� �Pw        Ɗ�}�D�  ,��       ��!�nC� �|M��si����U�H?�y��)O��       @w�jd=33�������dbb"˗/�ʕ+[����z �������#U?�ʤ��$�I�fw&�#5�N�l�]I�L�=%�N�=��X97ӭf       0X]����ݛ�<;w���ݻ�k׮�߿�%w�t�I9��ӳf͚�Y�&g�uV^��gbbb����ȟC�˸�����y�l=`�&����SSsN����G���7��<��$�%ٞ��IM�P�y��>Og6        ���q{�5۷oϖ-[��c�e�޽���fǎٱc�w~o���9��s�����/����{�	� p,K=p_�3�{�?��DR{9���$��lM�֔l�l��7d됷       0��N��}�ݗ-[�d߾}���333y�G��#��;���矟׿��y�+^���9�~���� О�}aV&Y�d�wN~�I�%��]I��lL�Ɣ�2���59�j,        �9�}߾}ٴiSz�^fgg~����<���y��s�Yg�MozS^��W����$w  ^��}�I�$oI�߇�s�Nesj6%ٔ����rY�
       0.������{��ƍ377�d�������~6g�}v����g͚5Mv!p ����\����Ϊ��^�$�3%_J�Ʋ.�f       ��ց��m�r�wdϞ=Mw������D���7��K/Ͳe˚m� �b�÷,��$kS�$��lO�WR���󕜔��59�v&       �hk����lܸ16lh�����lذ!�<�H~�g~&/{�˚�� �b��pVj~1�/f"��L�^�NɝIń�^.�L�        #�UX����|��ٱcG�����O?�o�1�|�;s�y�5����311���  t��vӪ$oI�թ�%��l�喺9W��si���U       �����M�k׮|��|�~ġC����>�7on��k'�à� `~��>NMreJ�L?�T��ܚ�sY���k���>       ����O���r����S�֚�o�=��������s`ɪ���`��$�K��\�嫩Y��|��6[o       h�ŉ��<�L֯_�C��ދ�k_�ZJ)��ˆz_�/���9 ��D���eIޒ�k3�j/�^�����V�}      ��Rkz�w���t�M#�q�]wejjj��m�6_� 0?���$L��L��������r�;       ��;t�P֯_����h���/d۶mC���q�w ������$�>�-Sy��r}�ʕ��ߔ       �%iء�m�ݖݻw���Vk�-�ܒ}����K�r �����$�*5�d*�j/��^�*v       8>��{o~���3�������[����vO�/K��`~���$L��L�us~��ra�Q        'b����={��/yh�k�'�ȦM��v?�;  ��������$�^�^{�@} �[�       X�a�_��3777����aÆ�߿h��  p�]��c��S���T��5�]       ��Foݺ5�>��������L����3`I� ��;/�$�N�-��õ�kj/�j=
       ��Zk���3����SO=5�{	�Y�Jq�( ̇��c9/ɇ�|��rK��ݵfY�M        �cXa�֭[����^]�q���  w�k"ɕIn�T��͹�nə�G       Ӹ�������R�k �G��� %�f6��^n���փ       ��5�htǎy�駇r�.��z�'�H+���  #A�ΉX���)����պ9�Ro�d�Q        ��e˖��z衇���~�\�T������X~4%��g[��C�ެi=       ÈF�����o~s������l۶��YNp������JrM�����u��W�       p��x�<x����n�:��8隥��5 ̏��AY��I�U�����       �����Nx�ǆr']������3h���$_���Z���       ,԰��۷o_���;��8� `|	��wf"��^��j��$       �777���~����ؾ}���!p _wZxKJn�T�[�       �a��{��I���}Fų�>�z�$/� �����%In�T6թ���,k=       ���ڵ���Nٽ{w�	0�Jq( ̇��.x}j>��l���ǉ�       @��ٳ���N� 0Hw�d]�Od*��^��z       @�<x���N�|  0Hw��uIn��|����c       ����=F���L�	0����
 ��;]�cI���rg��m��        �SJ�=��kffF��a?� `)�3
ޒ���˧j/�Z�       ����l�	��9 `P����[{��N�փ          ��%pg�L$�*5թ\[��փ          ��!pgT����3��k/�5�Z          N���Qwv��e*�֩���c          ��'pg�X���֩��SyM�1          ��	�YZj~.5���u���n=          �?�;K��$�\�Syo�)�          �&pg){ej>��|�ޗ7�          ���q���w��    IDAT=���떜�z          ���$We6Sus�M�)�          �K�θ����y�r{�em�1        �x(ř� 0w��ے|�N������z           pg�-O��9�����t�1          0��\���\{��n��[�         �q%p��;��R{�@�!        ��Rkm= F�����I>V{�|��U��          �8�Ë{W����\]��          �.���Srm�r{} ?�z        0�J)�' �H�ñ�5s����ܗ�          K���g���ޟ�Z�         ��H�����ϟ���          �@��i���rA�1          �T����5�����C          `)�É9-��j/��䕭�         �TJi= F����f.��T~��        �{j��' �H���935���\_{9��          5wX|W%��ޟo=          F����sG��C�fY�1        @;��� `d�ap&�\���R7��c          ���0xWd2����R�!        ���Z[O ��!p��8#%Y{��~='�        O)�� w���*�T^�z          t���omj�V��뭇          @�ܡ�U��������S[�         �.�C[W%�X{���          hM��]��+u*���          hI��pRj�w�������z        �xj��' ���C�\�U�R�7�        ,�RJ�	 02��=�dY�S���         'N� �7����#N�k���dE���3����[��tZj����;Y���~�A        �񩵊�`�&˺����A�eegMJ^�~��D�IrVj�MrV�s�\�䤦C�M$��L������rq�i=          i���A)�ɡ$;���Ů�5%�sN&��;o&���]��#�]�gc�/�\^���          �2�w)�I�����}���׳<�rQJ.MͥI�&�$ə�_
�Ǚȝu*W�����          ��܏�\��$��߮O�?�}*$��$?��'��!�G�cej����Ɯ��P��t�A        ���RZO ��!�^��O|���o�/Iꦜ��,��D�O��$��[�x���@~��6�j=          ����7�$�?��Z�,���ʔ\��mIV��Ȓ�Ù�7�T�W��S��          �b�h=`�)%s��l,��-��S���yW��$y��>���R󗵗kj��        :���z ������r��.7�u�Ͳ.e.��7�ܚd��>F�D�e*7�M9��          8�!+o�ֲ6וu��$�HrUJ>�d��4F�/g2w�^^�z          /�{Ce]�-�����RN���'�1ɡ��I�$�X���[         ��!p�rn��벾��{r8�H��$�d��4F˙������[         ���wP���.���e]~6%��7�lj����2ɟ�^>Vo�d�1        0�J)�' ���w\Y��em�+�rI&rY�?J���.F����zONo=          �C�>B���X���sr�M���zW��Y����sQ�)          p,�T����.Q��m�����S����Eg�P��P��ϵ          G#pq�y��˯gY^��ג��z�tZ&��9W�          /E�D��f_Y����ycJ~:��Ij�]tʲ�\[{�?����        ���U� �%p_bJI-ksKY�we"oL�Ǔn��N��$[��        㠔�z ���V.�}emޗ~^���I�m���xk�z_.n=          ������<Y��CY�W���$O��D'���|�n������=J��������f.����&����"��l\эHֈ�7�=�Yͻ'�J6�`�	5��z��B6�(�⅗�a���(�p��~�?Ԭ1*S}�����9�Ñ3��o�p���WO         @bྨ��2�?�����$�غ��V��o�d^�:          ���.�lJ�Ĕ�*ɭ��hjij>P{��֔�1          ,^�X��2���L��$w�n��32��^��       ����N��2p'��l-�sQ�����仍�h�)��ޒ�[�        �BQkm�  #���V�y�t�)۲j�Ir_�&�9&����<�u
          ���;�J98��97Syb���dK�&n�L�zc�n         ��a�ίT�}���+�yR�MI�Z71P�g:W�^^�:         �����GU�wJ7�'98��j��@����;Z�        ��*��N ��a��v+��J7'���Inh����$o����^�%�c          X���[��gsWM�$���a`^���zSV�       �QRkm�  #���)��t�I�K�$S����f*_�7g��!          ,<��J���������{�ٖk�M9�u          ��;s�t�L��$/KrG���2�/���7�C        `ؕRZ' ��0pgΔ�Z��h�f}�w%�j�ļZ����ɜ�:         �����9W�����7&9<ɗZ�0�vJͧj/��         `��3oJ7_�D�Nrz��[�0oƒ�y���C          m�̫R2]�ٔ���e��MI����{�o         �h2pg �D�[�yeJNI���=̛WgM>Roϲ�!          �w�L�fY�%ٔ���a^��-��ޜ�Z�          0Z������tszJ����=̋��-W{٧u          ����f�D�΃9$%�&�j�Ü�H����CZ�        @+���	 0R�i��-e"�$yF�[�0����˱�C          ~����5�9��6���=̩�I.�7�E�C          n���w,9'%�'��usj�t�:�״         `x�3t�D.ϲlH��usj,5�ɼ�u          �����T���nNOɋ�|�us���j/�o�)�c          .��2�Od[�'��us�?���E�2�C          ��rp��DNJrz�-�{�#5�ʚ|�ޞe�S          RRK7�����{�3/Ȗ�u�%;�         �=wFJ�f2�stJ�M2ݺ�9�1[�zKvo         @[�o*9'%'%�~��@��y$W��w�        �K���	 0R�Ye"�mY���m�80��C�1Z�        �\���N ��b��H+箬��9'�T�f�q��U���:         ��3pg䕒Z���L�$�i�ì��t�����!          ��;Fِ��4ON�׭[���$��N慭C          w��������s�L��aVvH��j/�n        3UJi�  #�����Բ>�f:�%�^�fe,��us�j         ��o �l�U����|4�Q�{������d�(9�u@k��?'�������u        0��Y�����zK��G�I�h��,Լ���<yc)�g����M��6?��       �֔RZg �����V��å�7&yE�-�{��7����+}8         `!2pg�(�����䛭[���WfM>Zo��S        �Ѹ� �c�΢R���,͡I>޺�Yya�'�uY�:         ��c�΢S�����KSsN���=���c��~3��         `n��(��Z���L�$�k�Ì��rE�%��         `��Y�ʆ\���$_n����G�w����:         ��1pg�+�|;��$��na��e<�����:         ��3p�$e�<T�95%g&�j�Ì<!�5���:        ~���: F��;��2����䇭[��=��Uu2G�       �$)��N ��b���t�7���$7�naFV����˳Z�          �w�%ʺ|#�1I>׺�yL��j//h         ��3p�_�tso���)9�u3�C���^^�:       �ū��: F��;�ec�������$���oK����˫[�          ���a;�n6%yV��Z�з�$��9�u        �O��u �w�N��k2�Ó|�u}+)9�N杭C        X\J)� `��Cʆܑ�iI�g�f��musέ5��       ��p�; ����T��q&��$غ�(yk&��Z��       0��� �1��(%ӥ����I���o����e�.KZ�        ���� �c��P&�ޔ<?���[��˳c>^oϲ�!        ,\np����,��\�N���ۭ[��Iْ��7eE�          �aN�u�!c9:�W[�з���gk/�Z�          ,v�0Gʁ�3��Sri��vd���[�{�         �����P���Y���ݭ[�ۓ�H���g��!          ���;̱R2U&�)93�t��r`�����~�C          #w�'e"��%I��n�/OH��zc6�       `��RZ' ��1p�yT&�$�|�u}yl�sU��)�C        ]���	 0r�a��n������-�eU���^��:       ���w 蟁;@9(��t����-�e�$������!        �7�@��a@�A�/K��$m�B_���Sus^�:       ���w 蟁;P�?g"�����-�eiJ>\'sj�        F����0`�d�t�۩9'�w��c<5��9�u        ��� �?wh��Ϲ���$[[���Jj��N杭C          "wh���2����u}�y[��]��Gl         搁;4V6�o�����[��2��+3�:         `�0p�!P��R�st�[[�ЗS�&��gY�         �����Dِo&96�W[�ЗdK.��<�u         ��3p�!R���$OO��-��I>W{Y�:       ��QJi�  #���L���INN��-���$Wo���!        �Zk� 9�0�J7�d"�Hr^���>S����O�        �s�; ����T)���7���-��$��7��!        ��w 蟁;��>��?$�n��v�'S���rH�        �q�; ���F@�ȟ��%Ij��v[���u2ǵ       �7�@��aD��|"����u��1���n΋[�        0xnp����)�\��g%��u�m�����9�k         0��aĔ��r��$w�na�������;Z�          3wAeCnLɱInn��v+I�^{��V��          ���%��2�o%9&�߷n�/gd2��eI�         �ac�#�tso�g'��u}95��W����:         `��È+��8KsR���n�5'��\Qo���)          ������D�m���n�/Ge:���y\�         �a`�D)��D^���-����|�Nf��!        ̭RJ� 9��Z�ys���n�/OH�յ�CZ�        0wj�� `���T��R�I�[�������       `n�� �g�TY�w'yU�m�[�n�I�:�׶       `��� �3p��tsI�'y�u�m<5�j/�h       ��� �g�\��S�9!ɏZ���J���^.�Wf�u        3�w 蟁;,e}�Lͳ��Ӻ���&k�z]��       �np����"Q���I�����-���1W�[�{�         ��f��H馗����-��)y$��^�k         0��a�)嶌��$��-��I>_o�a�C          拁;,B��ܙmyf���n�/��t��7�9�C          惁;,R��ܕG�1�Z�З�䲺9�k       ��VJi�  #������ �9)���-�e<%�ɼ�V��         ��a	�\9<[RsRJ��u})�y[&��zGvl         0܁�nɺ�,%h�B�^��sE�!{�         �-w IRJ��.���]�[��Q�����D�         ��0p�Y)��șI�k���o����9�u         �L��B)�������-�mEj>Y7���C          f����������'�n�B_�S򧵗j�       �J)�u �$�G�W*yO�W%�ֺ�����\Zoʊ�!        �Q��u �$w��*�\��%In�Bߞ��\So�ޭC        7������t�ɔ�8Ƀ�[�S�A���:�C[�          <w`���\����ߺ��홚/�^�}�       �Ţ��: F��;���D�N'�Lrw���,�_�^.��eI�         �_���KY��$yz�;[�0#�e�\^�Ϛ�!        Y)�u �$w�o��Ɍ�Ink�<=㹮ޘ�Z�          �<w`Fʁ�=��$�h���\S'sj�         ��1pf�t��L�iI�o�,K��d�Yk�Z�          ��R6�{y$�Hrm�f���m�̥�����1         ��f��Zyr~�myv�϶naƎ�X�T'��u         �x�s���sNNrY�fl��|�ސ�         'w`Δ��`��S���-�؊t���˅����c         �����Sec���W����-��iI���y|�         `�0p�\)�J7�%9�u�rDj������!        ����: F��;0/JI-ݼ)��naVvK�e���T��        ۫��: F��"0�J7�H��&�n��%��L����m         ,\���+���$�J��u��1S�z��	�C        �])�u �$w` J7�$yq��Z�0+����������c         ������ͧRrr�Z�0+%�I��7e��1         ��a�T���٘��-��S2���^Nk         ,������r��'��u��s�k/�7fu�         `��M�nz�S�|�us�ř��:�Z�          ���h��۳-�Hrc���cSsi�������:       ��RJ� Y�@S���c��&���-̉���rn��yZ�         `��͕n�Mr\�ϵna�<15W�^.��g��1         �h0p�B����9'%��us��䴌�:��Z�          ���e�<�sJ��ֺ�9u`j�����6w         ��1p�J9<[3�S��a���X��3���dNi         'w`蔒Z�yKj�IR[�0��L�_��|�ޜ=[�          ���Ze}�M��I�Z�0�jN̶�P7�u��^       ,,���	 0��
��V�ٔ��Ij�[��M�̗�9�u       �\���N ��e����'3��%��u���L����볦u         Ў�;0ʆ\�N����-̋��Ԍ��:��P��x�        ��*��N ��e����._�T�Nrk��ͪԼ;k������1        3Qkm�  #��)�ܖ��$׷na^��#��/�st�       �~�� f��9���T6&�B���љ�5��֛�o�         `~�� ��rP���9�1I���    IDAT��=̫N�S3�[{�p���r`no�����w(u�ޭ;��hi�@�
        `�#��-�����(5�j�ü[���_Z{�0��/eC��:�����:uERV�n���}k�/�uon�        ̡N� ��(�gk�巒�~�fY�7���j/�^�i4Hw����:�^�ĸ        ���y���n��$�I��u�<�In��|��2�:h�}�O^�v��]�d��-         0܁�t�$/N��u�$ɩIn���x����A���w��Kg��eI�к      �I�u��(�����s �|1p��ͧ�lLrW����%������i��,o5�8�����Ii�      �fC����y?c��R<'  �w`�)�|)����-4sH��c�U'����~��f�~�c���$uA�L      �`�ҥ��ʒ%KZ'  ���RY�o��#�\ۺ��vK�ے�R{���rZ��1���W�)���&yQ�      X���%�  擁;�`�u�'�s����-�Ò\�����{�yN�2C�3�����ޙR^Ӻ      ��vکu�P�|��+��N ��e�,h��g"'%�Ժ���"ɫ��g�&w�^>X7�z]��ʅ���ח䭭;      �d�ʕ����]��u �,w`�+%S���SsN����$���S�1���|��rZ�9{������^^�w�l       ��]wݵu�P�|��s�; ��x� �A)�snݜ{S�x��_{LjNLrb���^���s��|��Ų.�"��?z�q5���      �+Vd�v��?�:e(�^�z��0 X�<�E���E��|7���$�i���*IMrhJޒ����d�/$�j�����Pϖ�<����Ȓ�O$Y:��      Y)%��y?g�ڵ�������aWJ�����  ,`���S6���˱I>�d��=�����ӿ~b�L�^nMrCjnK���m��<�;���u������O�/      `(���I֬Y�vءu  ��;�(�n�^o�S2�O�'7uC�ƒ����'�u~����˖$w���� %��f*��I�d"�SJ������'���       � nq�{����G�^{��Rʣ�"  $w`�*��z}���\�䅭{Xp�'�'5�$I~��Ү���3pO�z@]      �����=IV�Z�իW�{���������: ����`�*�L�EI~�u       33�۾8����3�v�m��^��.x4~ ̎�;�蕒Z�yGJ^�dk�       �3�1铞��t:�wn3���q0 ��6�: `X������|,ɮ�s`�ݑdsJn*�͙.wN��j'?,��R;Y^��K���d�کOJ́I6$٫m:      ��N;����/���7Z��ҥK�nݺ��e� ���������d�LͥI�Ժ�Ȗ�\�����r�gl��L��_��X��1�<;ɉIv��L      �RJj��~�a��[n�e g��:(;��@Ϊ�� ,b� ��L�zc��t�*��Z�@cW���Oo����������9���&�5�E���;gꡗ$���c���     `>�Z�*��on���)�dɒ|��9��b� ����e]�9y$'yE��Zk��ԩ�_����~>Z}Ɵܟ�}I�w�y������L�$��
     ����$9�c�o}+SSS9���?<˖-k� �"�i 0���y8yej�I��~���5��Cw;��{���V��Ͽ���M/�NOr� �     `a��߻�K=�Ё��ڪU�r�!��<�� `��k��Z������[��|���k�o�:s��V�u��[��~֦��:sӿI)�Mrw�      �U;��뮭3�U)%O����fbd� @b��]J7J��Ino�s��^UǷ��Y�����i���>���n���&���=      �����r���g||�uʼ9�òv���0r|X f��`;���>���s�[`�L'y��=p��oxߝ�c~�Ǿ���Z�����?�'�      �+�R:,]�zu�9昁�7Hk׮�G1�3��Y(j��� `d�����=�+ǧ���-0K��Z���6�^y�G�Z��:�e�Z}֦�TjNM�H�      �y6lȁ�:cN�X�"�}�s���L�� ̎w� }*��L�$�.ɖ�=0���:����Ǫ�7}�f�yI�o�      ?o�ƍy���:cN,[�,'�tR�/_>�s�� ��f�t�$OM��-��J�r��/���)3��Y_ѩ��<Ժ     ��TJ��ɝN'�|����ܹ�dɒ�x�Y�re�  1w�Y(�|-�9<ɕ�[`;L%�+ϼ���!�����n:�7�lk�     �p��=I���s��'��M�˖-��'��=��c�g��� `x��R9 w�<'%�n�_��z��3/�x뎹���}���ݺ     ���j�~�	'��ٳ���;�%/yI�����7� 0���@٘me"�$95Ƀ�{�_+Yu�E�i]1�v;��?�%j�     �pj5��t:9���g<#cccM��'<!/}�K��.��N �$� s�tsIJ���ۭ[�gJrkƖ��u�|�^2~z��[w      0�Z���vs�)�d�wn���t:�s�1y��e˖5�p{;  ���`���|5c9:ɵ�[ I�J�u�����[�̇5�ϏK'�MR[�      0|Z����c���o�f�<�ȡ��}�ڵ�����<��On���� ��d�0ʁ�3w�i)97���T������ZģUo�tMI.i�     �pj=��G����e�g�}���X�"�w\N9唬Z��iK)���  �i�u �BU6f[�sj/�&y�]��ݷ���m�#ak�~�x휜d��-      �RJjm/٪U�r�I'����W���z�;{�w���n�;47�� ��`��n>��#�\ߺ�E�g���[G�g^��$�j�     �p�1�n���>��y��_��;,+V���s��ǳ�����O�+^�t�A��  �7�@��-���-� �i�{XX2�w����:����ؙI��O      Y?T�M�?�r��u�Qy�S���~����;��|'����2===���e�]��^{e�=�����,]�t��熁;  ���;���}�P��k/���O���8�����o�����������?>mSj�Ժ     ��3�#��']k׮�ڵk�$[�n�}�ݗ��/?����([�n�֭[���g||<K�,�ҥK�|�����u�]�r����N���Gg� ��1p������6c�pjj���4]:�nhaz�n�t��;      �԰��ޒ%K�f͚�Y��uʜ+���(�� f��: `1*rcv�S���uҵ���g7��ha�7]�~�u      �� �=�)����S�$���a�(�^Һ��Z�_�n      `x�E��9  �����2�O$9$�Z��0����Z7�4>���~      ���`u:�9  ���`�n���15�d�u��&�\���~�uGK����ۓ���      7����t̓X\�� ��y	0$���Z��m�αInk��h*ɕ����      `�3� `&��Lِ/fYM�[=%�˭�A)�R�      �_)���b� ��x�0������+��,ɽ�{�N�ܺaLM��      ��s˸ ��0pb���&yrJ�j��hغm��{�,��y      `���}�� 0[ޙ��ͷ�.�J�$��a�mY����S�a����Il�     �h1r��v  �w� #��L�n�0�Y����=���['�RR�      ��t:F�3�y `�����!��D6&9=ɖ�=���N&%�      f�M���\ 0��[ ПR2�dS��$�Krl�$f`��w�w�y+����o���Y=�R��w�yOJ�����ַ����U�<7�     0c?m�Y��x�  0�FT���ze��5ys�w$١q}x���k�c?���N�ejV�y��҉Z��I��t��ȿ��E��     0{??�6t��:�N�  (�4FX٘m��w&Y��s�{hkI��-.;�      `����_�|  0����ͭ�ȳS�$��%����h      ���w��q��}��.^	����H�vb5�"�V�Jr�Kr��qΓ���]ƾ:���L,7m����?�+�k'#�"�@r��4���ݜ9�M����c)nƮ#Y�lYR$UI�/ @�������@S6%��>����������b�Xi��[�G�R�J�2���r� _�F�~ ��)��"�[�_E3F�gJ��F���+�CC��t      �OJi ���=�F�KG ����g�;b&����]D���y�J䘈Z�]�ܶ�7E�P�      ��A){�m��Ϡ�7 @;y�	Чҭ��E��#➈X-��L~��T��t      ��Z�����  ��Q(@Kc1�_�J�="��t�oG����*��KG      `p�������  @)��tK<��OE��E�.����!-���r�x�      �^.���6z  z��;� Io���R��M�>�/-E�\:FQ���房V:      ���{7��J�6�C�t��< �
�NL����ơHq[������Z#ш��R:FQ�OM���s      �Z�����ʯk����^΃�� Z�#U��n��ӭ�3�����:ߛKG(+�ϖ�       ��Z��v�ޯ����v� �f
� .�������@D<_8-�}�b��g��C�*)�ϕ�      ��;7��֦��*�_��~�3ڡs����)�)EN�Dl�[#ǯG�|�Llܖ��qy ������7��      �q�����km��� �~����ͱ��wG=�)Z�Ll����@���J����         ��)��]�ętk�r4��"�xD�Kgb}ޒ.��{�xG��t����-�        ��Sp�5�wċ�`|$*�W�[E�F�L\��J�z���?�m         z� o(�ϧ��h�;"�3�,��7�r�����?R:G'�;�������        ��(�p��;��`�|D�`D|6lt�v�T�ܟ?��j� ����/}2<�      ���R� �� X�t0M��F�-"�E�r�L\[����ɩ�_:G;;4��)�;K�         `��ذt[<�����ވ�XD���5��?~������9�a���{{����s         �
� lZzG̤�q("n��Cq�h ^-�X3�g����JGi�3�������lD���        @k(��2�`̦��xSD| "�c�H|�_����|�P_��χU�+�OG�-��       @DDJ�t �}Qr����QK�D:?�����LD���E����S���
��O�?[:       ��9��  }A���J��W�������F�gJgd)�����V:�f�?|ǡH�+�s         �z
� tD��8���4n���'#�D�V��XD\�T"��>v��;��C�z�q@Α�����g��       �wJ)��  }a�t  KJш�?��?�_������q[�d�u�����L�ۥ��c&"�v,@�_����d����>r��h�������I��v�,         �OOmn���[�t�5��[�"ǏGĿ���ҹE����Ks���Y^���;�2�c���        ���; ]!�=�4�_�-�7r�/">K� ?Ԉ�:w����A�����ln��"�*�        ��*  ��������|~.��R�d�xD�͈�^6]�ڙR��s�~��VS��λ���K:w�߻�����s���Y         �w �֫��/�x��OE%���xOD�-������ی�7����Ǧ~��|�3\8�w'�1rgD��rĖN�        �,w zBzs,E��r��D���&"�K��#�y4���{?<=2T?��W�ϳ��p�C{V��w6s�r��        0���I�`<OD����+���������_4\�)��Zc�=w�G�}T��Rsˉ7���V��>:z�^�os��ֈ�#�:        �ޤ�@�K������^�D~2D#~,"~<"~,"n��T.aOI)�7r�wK�t���;��"�D������ӡ��=(z��ܶ]����s�w�6V�Z$��        �6w �N��8'^�D�Z�������#ǏD�m1Q0b�ڑ"~&"~�)fw�������S��K�bD^L)-��"�ֈ�="ޜ#�6��jDD�\�      �VK��= hw �^��8��+��xe�{=~0R�`D�#▰�}=�r��EJ���w�UZ�y�����+        ����@ze���������1͸-��W"�M��HqSD��Ke       �_��w hw xE:��W.���2v�������)vG�=�bo��q���+         l� \��Wb>"y���#1#Q�FLFD�pLD�H4c(Rl�����������֦       :��v hw h��Θ{�������g��ɩ��o�)         t�J�  @D���Ʈg����Y         �w ��';o�����Y       ��R* ���; t����;�(G�v�,         �i
� �eR������ E�_:         t��; t��"���G#Ǳ�Y         �S��K�y��wFđ�Y         �����y�]��J��t         h7w �Sw�'��o��         �� =bׯ~򟥔~�t         hw �!Sw~�n%w       �.)�� �o(�@����wG�_+�         ZM� zЮ�>uOD���Kg        �V*  ؘ]w}�ވ��t(e1�x�        ��          �

�           tw           ���;           ]A�         6!�T: �w         ؄�s� �7�        `lp��Qp          �+(�          ��          �

�         �A)�H)�� }C�         6!�\: �w           ���;           ]A�          ����          @WPp         ؤf�Y:@_Pp        �J)��@��9�� ��        `���Yc�;@k(�        ����Ov hw         �M�9���"
�          ����Z:@�Pp         ؄Z�V:@�Pp         ��ZG�         `�ZG�         `VVVJG �
�          �s�����1 ���;         lPJ�t
[^^��s� }C�         `����JG �+
�          t�ҥ� ���;         ���u�ZL�         6(�\:-,,�� �w�        `RJ�R*��KG �;
�         ����Z�KKK�c �w         � ��ۅJG �K
�          ��h4��ŋ�c �%w         �u�����s� }I�         �:5����/�o)�         \��g�F��,�o)�        ���JG�Ö����ŋ�c �5w         �7�s�����1 ���;         �8�|�j��1 ���;         ��X\\�����1 ��;         �kq��    IDAT��j133S:��Pp         ��f��O��F�Q:
��Pp         �9�8u�T�����0P�        `RJ�#�&k��˗/��0p�        `rΥ#�k��K�.��0��J         �^d�{�i4q�ԩXZZ*``)�         oee%N�:����� 4w         `�-,,���L4���Q ��;         0��F�={6.^�X:
 �Pp        �uJ)EJ)rΥ��A���q�̙��륣 pw         � ���T���̙3���X:
 נ�         ���{��z��������@Sp        �uJ)���uj4q��p�b;@Pp         �ΥK���ŋ������C�        `�lp�N�z=.^���󱺺Z: ��         �����t�R\�t)���K�`��        `�rζ��l6cee%VVV����q���h6��c�B
�         �N����h4�^����j�j�+��Z�V: m��         lX�шF�qe���?sίڮ��v�����sα���z=��z�;�- �E�        �WY+�_]:_]]}U�}�m h%w         P�������Z��e�� %(�        @��9G�V����X^^�Rj�9�� ���         }�^�_)��]���
�         ���f\�|�ʥV��� ��         �R*!VVVbqq1._�KKK���n�M �w         X��s�Bs�V����XXX����(����;         �S'�̵Z-���caa!��z��>
� ���         ]��l���B������r�8\w��Pp        �.���sss���9��qX�j�Z:@_Pp        �uhǦ�����K�.��lگR�l�v�R��Pp        �"r�q��Ÿp�B�j��q؄J���3r�n ��         ����ΝSl���Û>#��� 
�         �1���q���XZZ*�jIS� �        `]RJ���z�gΜ����6$��Vlp���V���        ��.^�gϞ�F�Q:
mҢ���V���        ��F�����> FFFZq��V���        ��._��O���}@���n����D�y
�         �B���q�̙�9��BG�R��9�JE� �        �eΜ9sss�c�Accc-9'�t�%�8w         ؤ�s�:u*.]�T:
6>>ޒs����k�A =n�         N�}p�h���o��o�k�A �N�         6affF�}@U*�Vܟo�! �@�         6hnn.���KǠ�-[��䜔�S-9�(�        ��j�8{�l�411ђsrΏ�� �>��         0339��1(H����        `RJ���KKK��P���X�䬔��-9�(�        �:��Ζ�@a۶mk�Qs�v�z�U��:w         �N)�X^^�����Q(���?=t�P�U��:w         X�����(l||<���ZrVJ�O[r@�Pp        �uXZZ*��&''[vV��K-;�(�        �:�����@A�j5�n�ڪ㖆���ܪ� �Ak^        h���~NJ��祔�	xE�9��f��}��V��~����^ �*
�        P��J��Sl���~��U*�wh�����RJ�s��V�G�<�(�       @��b;Q�}���
�9���m۶��P몗)�ײ� ���;        �I'K�o����SJ��A
��۟<v��ӭ<�(�       @�國��������a}�F��u��m�y)���e��w        h�n/����܊�p}VVVJG��]�v�����g[z @�Pp       �MX+��b��j��p}���KG���۷�t{{D������[y @�Pp       �j6��#���;���s�j��1谔R�޽�����V�/�       `�
��N�����J�055CC-�[�6��m� ��R:         �A)�_-��fs�o����e�fxx8���Z}��?�O���C���;        \�A,�_m����V�E�����At�7��U,RJ�j� }F�        ^�毦�ΠZZZ��p_0@�o�[�li��ONMM��V
�O�J        �n��}mk�Vo5�n����z="����P�ٳ�����9t�?. �C�        �A���]]�Ur��5��+��#��7��j��Ǿ����oZ}(@�Qp       ���X���u�RRt�o���]y�KJ��� عsgLLL��ܔұO���-?��TJ        �n�ܾ1�3��ٳgcy��}d���766�w�n�������k�� �F�        B�}�\w���/ƅ^�1���V�V����zE����_h�� �F�       ���ܾy9�h6��G����b���|��ݾ�WJ)���CCC�8�啕���q0@?Rp       `�)����^����O���m���ٳ'�l�Җ�s�;~���Ї��T#        ��f�t���s��R��n�����ܾF��?MMM���d��lff�S�:�)�       0�U�gm+~�R)�K�9Ν;.\x�ϣ�l߾=v��ݶ���?:q�D�m ���;        g��M{��N/���q���XZZz��u��_�n����k��)�������m ���;        E��slr��-..���L4l����ؿ;G\�9��� �J�       �����y6��m��z�9s&��u�?����D8p���K9�|�}��Զ }L�       ���l6KGH
�t��s\�p!Ο?�����{�۶m[�7�G�����w�'�:��)�       0z�ܾ��.\���Ũ�j����F#""FGGcxx8���crr2�m�V8��Qr���s,,,���l�j�M�C���{��{�BJ�"`��       ��f�gΜ��'O�ɓ'�ܹs���t�_?44;w����Ǜ���8p�@����1���#��J�tH���W�GoڻwoLNN�}NJ�ǎ�˶�c
�        ��n��~�����7��<�L���l��z�gϞ��g��c�=)�xӛ�7�|s�t�M1<<��ԛg�;��h4b~~>���cuu�e�*���J���틭[��}VJ�sǎ�ݶ�s
�        ��n*�6�x��'��G�������9ǋ/�/��b�-���|�;;R�
����r������B[~�����7622�������9?[�V�� ��;        }+����f��?�x<��#q�ҥ��]]]��{,�x≸���������N+---���b,..�t[��t��	�g���w�ިT*�w9��?9r�=�\0
�        �F�N��?��?����b�F|��_���z*n������ۣZ�ˣ��f�_Uj����Mw�T*q�7Ķm�:9�LOO�����;        }����������O>�d�ߩ^�Ǘ���x�g���~w�ٳ�X�f�٩��􁥥�XZZ�˗/���R��m��e˖��bxx��c�LOO�����;        ����l<��E����������>?��?��v[�8pE�9j�Z���\�,//G��,-"ܻU�Z�ݻwǎ;:=��_~���� �N�       ��Sr{��O?>�`���"�W�ш�z(fff�]�zWT�Վg�9GJ��s)�^�����.k��n-�wk�A�cǎؽ{w��������܉'����  ����j�     =�DY;"�����z����O=�T\�t)~��:FFF::;��F���/����V���'�4���9G�ٌF�����VWW��ٴ���سgO�������F�}Ǐ�\b8@�Sp  �r�=�\�     =e���w�ގ���_��W:>�N�<�����{��btt�������ԩS�	���FGGcjj*�m�V*�j�����/�
 ��*�        @+�ܹ��3}�ў-��9s�L���a�����ݲeK�K���f�t��666�����)Yn�i6��>r��� w        �Ɩ-[bxx��3�z��җ��љ�r���x��:^�ݱcGG��F��^���D���o����-�u�֒Qfr�?y���?U2� Pp       �otz��3g�������?�g�љ[�n��RGg�z���y�����x�[�7�xc�����t��l��}���x�  �`�t         h�J�����<�@4����Gy$���o}�[;2�R��֭[caa�#��S�Vcbb"�m��������j�����ϗ0(lp       �/LLLD�ҹ:̃>/^�ؼN{���ҥK������^�f�t��3<<���q�7�M7�����r�W�Ə9r���A ��        �N��}��x��g;6�����x���=�yOG捏�G�Z�ˍ��s�=odd$���b||<���cdd�t��������s�=�{� ��       @�V��e˖��Z]]��~�#�J{�g�[n����-m��R��[����|�g�F(�_��R���p���h������HT����K�yzff�'Nx�@
�        ���������?��XXX�ؼ�z���?�J�������Z�^p�T*144���Q�T�R�DJ��?�~{��#�Uh�V��������/MOO�n�  �L�       ��ש��Z-{챎��sss���O��7���Y���m���j�����k������<��˽X�T~��ѣ_)`�)�       ��:U���׾�Z�#���W���x���vess�T����Z�Z������B���X�������ÇgK@�       ��V�n�z�>p���\�p!�{馛�>k˖-
�t�^��>66[�l�r�]������?U: ߦ�       @O�����{.���;2�}���H�}||<����>֫�l���]��jl۶-&&&b˖-m��>�g�J��=z���� �j
�        ���������7���/��˗۾ztt����FtSq<�[�n�Rl�l=�rD���/�|ω'�� ���       �i���m�q���x���>��5��x�g��nk뜡���V��h��=rΑs.�abb"�o�[�nUj߸�W*�_>z���� ���       �i###m���K/E��l��n��/�������R����*UnO)Ŷm�bjj�#�u�*���J��ǎ���Y xc
�        ���R��s��ɶ���N��f��J��s�����*�~�K�Z�;v���dG���ع��?��j�8~��j�0 \�        �YCCC�Rj���^z��3z���j�9s&�����9���m=�k��s��u_U�Vc׮]�cǎ�ܷ���������o?~|�t �G�       ��522��+++q��Ŷ��
����ߨ��R��;w�Ν;�Z�njր��������#G�̕��(�       г���_�p�B�g�����wF|$۶m�ݻw{b��<�R:<22�;��sϥ�a �w        zV'�Н(t�w�f7�_���h�۷/FGG[~��hF�)�O�>}�N�8�(��Pp       �gU*��Ϙ��o��^҉�?WX�Vܧ��b׮]�Rj鹃 ��l�R�LJ�w�=�B�< ���;        =�E���ն��%�Z��3��6�f�%��ھa/E��U*�G��ӈh�J} ���;        ��W���a�5ݦ�w��SSSn�ק�1���r�4==�h(�w        zV'��
��h4��hD�Zm�`�I�R�}���֭[KG�f��RJ�^YYy�����CP��;        =�E�F������l����m+�fC+l��822����'�Y��x1��t���ZJ��x|׮]O:t�V: �A�         ^�F
�����T*mHT�R|k��b�y5�49"V#b��YL)���#�LJ�|D��9����VVV^8~���� �u)�        ��Xo�}rr2���ۦ4mQ��oF��R����x)�t2������̉'�� ��         ���l^���ܹ3�����4�V������9?Z�T�T*q�����  B�         ^��np����ݻw�9��土��?��?�G��+�	 ^��;         ��-�7s�G��=<<��Ç�, ���;         l�Ν;������҉j���>�l�0 �
�         ����������سgO��\�rD|&�t�رcQ2 ���;         l���H�߿������DD������R! ���        �5���j�7�xcT*�'�S������N�vSp        �אs���8��Ý�r)"�����:9 :I�         ^õ
�SSS1>>ީ���o������鳝
 �(�        �k�΂���h�ڵ�S㟨T*:z��W:5 J��          ݪ�l���n�!RJ�[���#���46�        �u�������v��fD|pzz��v�nd�;         ��j��v�j��?�V�?��� Sp        �7055�j�]�爸{׮]�;r��\�� @/*          �Y�Z����v��s�[��w��k ����ݼX��e ���=_�q��>��w3;w�+w�F!#2E7�҅��� F�U��T�d$2$*Hi 1	�m$�4-�IcHȘNz�Ǆ$ӝ��:Oi�J�']ϩ��y?(8u���.��         ����F��f}'"�>�L��" .���         0�������YD��R���xl� ���         ��p8���KǾ6�N�����K�E�;         |kkk�#s�������        ���n,--�L)��d2���� �@�        �VWW�楔���ի�*
 ��         ����s���K�"2p        ����b0��;��g�}��o�
�E�i�          ̛�`)�"Y9�k���SE� `���         )x���;��o�
�Eg�         �����~{�k�� `��        �Cz�^���v:�����0p        ��t��1�{{{wK@[�        �))�����1�;��{K��61p        �S��ȴ�c{{{�J@��        �)%�9�� �c�         ���Μ1�N��@ hw         8����+׮]�\�. �6�         pJU�yZw�D h#w         8����f� �F�         pJ]�g�~J�?
U��1p        �S:�Ι�?�N_-T Z��         N��zg�8.� ���         N���g��S� ���;         <�R:�����U� ���;         <0"�t������1�        �KKKgΨ��� @+�        �+++gθw�ޭU ���         "�.q����^��} ���         "��a��/GD. md�         ���v挜�g
T��2p        ����~�3礔��@ h-w         Zocc�T��; ���;         ���tb8 10J  �IDAT��9�c�  h)w         Zmss3RJ%�^�L&7K@[�        �Z�n7���K�}<"r�0 h#w         Zk{{�����9�M�  h1w         Ziii)��a��iD|�T ���;         ��R�������0�L�\2 ���        ���F���JF~�d ���;         �����.]*y���?. me�        @kt:�x�'J�~x�+�C���        h��R\�r%�.�;�N�[4 Z��        �V�|�r�ұ7G��GK�@[�        �𶷷c8��9�����x0 ���;         m}}=677���omoo��x0 ���;         k}}=vvvf�]Uջvww_�I8 �T��         01�f��s�������$ Z�w         �,��UU���� P��         ,������ܜ��z���, ��2p        `!TU�/_����Y>s\��/DD��# �V�         ̭�s���߿��zq�ʕ��z���;������# �V�         ̭�2n_]]�˗/GUU���O[[[�;�G ���        ������h�����ܝ��3������c �V�         \8+++����ι��~i2�|����2p        ��8�������{��A h+w         .�������>ϫ�;>>���| ���        �������(������s�|�����x|�\�3p        `.�z��F�������u�c�=��5�8 ���;         seii)666buu��
�"�7�*  me�        �\XYY����XZZj�ƽ��OM&��M� ��2p        �1u]���Z\�t)��n�u�s��L&j� ���;        ����~:��i�5������RJ�����0��a����q?1�L���" �f�        �&����ӣ�����sڝ�x�x<��t h;w         f�������?u]7]�Q�>�N�vxx����  �         ������1h� ��ߧ��;���" �w�        �}I)�1f������GUUMW{�r��t:ό��5� �?�         -�R���"��]���������D�ۍN���纮��}9"���������i�e ��f�  0�zꩦ+     ̭�s䜛��<��MW`1}3��3���Ϛ. <���0         ��>YU���|s�        �Ev7"~�����>:::i� ���        XT����gn6] xk��         @aw#�W���~ĸ .�        Xӈ����~������  �?w         .���_UU�����7�� <>w         .��9��㣦�  gW5]          �g#⧷��~p2����p�        ����r��������N�. �e�        ��{=��������. ̎�;         ��)��ݿ��k׮�n� 0{�         ̓����D�����_GDn� p��        h�ݔ҇s��?>>��_|�^Ӆ �f�        p�r���#�zD\�v����ۻ�t) �y�         ���)�����u]doo�VӅ ��c�        @i_��)��铓����_l� 0��        x_��/=�y9���tz������?���w .(w  �9�R:j�    ���9�pD�@�=(/�������6���$"��Rz="^��;q��w��9�|rrr�Ν;_z饗��hY `!}���X#�_    IEND�B`�PK
     D"BY��_3
  3
  /   images/1ff35573-e276-4514-8c59-6294c96ecf57.png�PNG

   IHDR   d   .   �!�^   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  	�IDATx��\klW>3���?�vR�ql7M���aBih 	�F4��hS���H�

�U���u� ��[�(!IqS�R�j�4&�;i�:[�w׻���|wv���cg/�u�I��uw����{�w�4`H�b濙%�k
�ٟn�N�W�éR6���KCCC�v�����$I��$���|�aM�<p�@ʿ�Al@2vPq�	�L��᠎�jii���2ڲe�,��,��=�}��7�~�o�.>��~��Cs���\AY�)�1::J�XL�c+���b����0E�Q\n`6�?a�Z̜	[w�\��4�
�"���(JB��|>��}\��y���y�j�̝�h��t1 ��������X��rrr�6�������i��̏2�j����ee��UUUTQQ!���A�Xyyy
�(>ȧIp�bA� Q�������w�gQdvk޴��;�oN�G9��9c�ڲ��1��Ջ�x��^E�2�� vݫ���vH*�Y3J#
��Sv�y�F���|
!HT��By,�|�{�1J��i�D��O1ױuT�y|բ��j^ՈcwH�V���RJ��@.i'Iי ��L*H��ͤ�wyh��3�PN�������v�j�**b$}�O���#� 0ہ�����TZZJK�.�lc� �������137~��	�Ht٫ju��+�Q%���3�|��a[Hz�$������Vjnna�֭[iѢE��OD�@�c������������Gn�;�>�Z*�B�QP���u��r¯�����cتjz�p���OИ]�/3_3��_�����0��3�K7!ǝ�xvb4O`η�3��"��V|ְ�y1Q9n�O4M�.]ҷ
�"�"��0�M7� 1�a�$������h�8.o6j�0m�{�<y7P���'�lo&c��Y3���#�1����9,b �:Dzd���drG6� ��O7j��41NG"#�L��Z�4>:zs���H�̤�1�!e�?�>�|��b\�)��{|k����8v�#
`�:��ac.$a1�1Ě����2_$}�`��[�P
b��LwWf!�a	��T.m&� c�
��b��(�1TU�'��nJ#YɎ@" ����I�������@�������7m!�8�m�9XFB�|�]�{�r|����5 �h���T��)�!_���b!L��_YYI۶m�ˮ�>����0�}�k���N�ec>�l�J��'_M�ҫV]UN��������~����w���"d����.^�H�+J� 4���Lit��g�-[�M�����A!�����g�v�|����vwM�I�i��)~�9��(+$g]�k&��+W��,)�U!Z� �"����療��D6`%��� 񋵩��O~�܉?z��G���X ��$)\��˺�|�k �������^��h�����C�O0	h3�w�*w�o�N��p�7�Ap��W>L���p��OJ͗Y_t�|����Q޾ig��o�7=!����?�)z ���ڵ�x �or�Oix��a���YN'k�厰�dG؋��\�ѣGi͚5�v�Zۑ�b	�+ H�����-̳�=��)�03qc�AQT�V�Y# Az{{EZ�������S���&-A���I�:YǬa��|��i��	igS�l�1�Ng��|�t�YA,�Ę���Ux�՜G�W����kMY{� v��g?G��g��lG�$��q��MI&K����l�anX�g\%�*c>�\�<��,�F�)D9����R/��]���q�6� �q���"�W��3_���K��9tn��w�F����6�m�K�u-����`��XS�JЩ���1B�G��������n%w���HԈ����{TRT�R��DR�����yqu�0�G�%^�1k�9���+�]��z��8�̿zK,�~�oJ�EXz_گ���JJ�"�d��@�ŋu�m��wۘv�iqa }|q>�t�q?q��v?�_^�����>0Ԑb���Ⳑ�]�z5����e%Is QN2�3�ļ/Fr�S�_�i YEx�~���2��,c�,� �t�b�!�!������"�z��5Q"&Ǥ��b������ҵ@΀�,��&����s�GI�X�e�(��܈��+A��X�`d���&�dd�/�L{�rB��bx����DVbĳ�R��Ф��7���Q�$eOrр񢧵1,���/��%%%�����l�̉ �P��������K�:���6���Z@�c��.
��=Â��g���O/Y��������]�Q�E�\��46�]̇������6k0'Q�}
�Y�v�+W>��Y�h�U��7���\��� ^��z�ϝ:uj!��9s&�����d�?�`]�ḣ��k��(�ǌ�Qbd����-�Ik�S�l�C��%�KX���Й��%vO�g<���شc�aM�a�}�=�
�7    IEND�B`�PK
     E"BY
�8b  8b  /   images/a7e3301e-fb46-458d-916f-a05c0bde95f4.png�PNG

   IHDR  �  �   ��O3   sBIT|d�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<    IDATx���]l��}����%R�(��(�"mY�-?(˃���S�$]Ңht�:l��u����C�m�i˴�Л]�z�a7	$C
�hs5�r��b9�]�ReZ�����"��8�BQ<�����z��s>�o��/S  �laa�G�"⹈8Px� ����N�*=Z�7�7�^(=   ��.Eę��}��� "6K ��T�  ���=�"�E�gC�     t�LD|:���^8z��J ��� xU�s���C      �ӓ9�?>z��ϖ  M� ��������K�      �!�9��>??���C  `��  <P>�R���w      찱�����=Uz  �� �I�."z��      �TUU���8Qz  �� ��ѣG�^D�.�     `�����ߔ  �"p �����8�s���w      4�_=z���G  �0� x �u��#��;      ��9/�  � p �A�"⟖     РO�����  �iw  :onn�q��     �&���Xz  �4�;  ��R�g�7      𩹹��,=  v�� �N;r��#)�ϖ�     PBUU���  �Iw  :������     Fק���*=  v� �NK)���      JJ)���  `�� 謥����;      JJ)�Å��=�w  �N� �Yu]���      Z�@���K�  �� p ��r���     �6H)���  `'� 褣G�.F��K�      h��.--�(=  �� �N�9��     �6?_z  �/�;  ��s�L�      -��  ��� �E���'K�      h�g���N�  �C� @�,,,<ӥw      ��`0���  �~� �ϔ      �R�Pz   ��;  ]���      Z�������#  `��  tʣ�>�;"�)�     ��R]�~.  �%p �Snܸ�LD���     �bw  :K� @�|��      ������  �!p �k�      wwpaa�åG  �v� ���     ��L�  �w  :c~~���8\z     @��?[z  l�� ��H)=Wz     @���9v�؁�;  �^	� �ӥ      tD������#  �^	� ��;     ��?^z  �+�;  ]ы��Rz     @�|��   �W��  `+���zO�[UUU���݆Q��������p'ccc�k׮�3    �j}}��az�ȑ#�o�����C  `�7  tB]ק�z�~����1111>>����v�~����cccQUU�z=A;���<fggKπV���?O>�d�    [���q�֭�y�f���ō7�ڵkq�ڵ�~�z\�v-rΥ�ދ�~��\D|��  �*  ]�����XLOO���t�߿?���SSS�gOg�     ;dll,���bϞ=q���;>���o��V���ƛo��.]�˗/G]��ݺ���C� @�� ���LLL���|������LLMM��.     `D���8t�P:t�����|�r\�x1.]�/^��7o\�#>Qz   ��;  ]PE�������Ǐ�������     �]�^/>�~�sׯ_�.�믿���zlll\��7B�%G  �V	� h����G��ޭ>_UU;v,�񘙙�4     �199'N��'ND]ױ�����Z���q�����,..>�ꫯ�m�� `;�  ��`08���RJq�ĉ8u�T�ݻ�     `h����������ӧOǕ+W��^�������J#��pD� ��;  ��Rz_����8p �}����      m355SSS��OƵk��ܹs���/�[o�5���9�DD�ǡ�  � �;  ��s~�n__ZZ��~������     莽{�ƩS��ԩSq���x饗��_����}��҇w� `���  `��^_8~�x|���     �6==�>�l|��}�C199��/�����=;��  0,w  Z����c�؝�v�Сx��g#���*     ��ؽ{w<��S��}.>�āv�e����x!  6g. h�7�x㉈�u���>}:z�^Ë      ����8~�x?~<^y�8s�L\�zuۯ�s���x~� �p� h�������gggcvv��9      �{��cii)���ę3gb}}��_#���� ��� �vO��sssM�      (���x�������g�Ɵ�ٟE��^^���  ;�*=   ~�������ɦw      �{��x�gⓟ�dLLL��o=y�ر�a� ��"p ��N�      �6�����?��1;;���ҿu�����  ;A� @���x�N_�r�J�S      �eϞ=�O}*�����|J��C�  �M� @k-...Dľ;}mee��5      �������x���o�q�;  �'p ��r�'��k/^����&�      �RUU�},&''����  t�� �6{��="��_lj     @��޽;������9��GDjf  l�� �6�k�~�ܹXYYij     @�;v,�����ȁ������  �!p ���q<��󱶶��     �V��*:t�gRJw?�  �	� h����������矏����     �j9���SM�  ��� �VUD<������<������-     �k0ĥK���L��Ɇ�  ���K  �;YXXX���[}��W^����|�#����5     �����o����]�I)�� @��� @+UUu�^�+��_���bmmm�      Z���_�o~�[y��� �b�Y ��꺾��="bee%���/����NO     h��^z)����G]�[y|����C��  �%p ��rΏl��޸q#��կ�ٳg���      �s�ʕ��?����7�qO'�����,  �/��  �NRJۺ�~[]���o~3Ο?�=�\LOO��4     ���_���ַ⥗^�ֱ������/��2  �w  ����._�_��W�G�~��111�/     Ш�s\�p!�����������>�S�  `�	� h�	�#������w������O�O<�w�ީ�     �����p�B���k�ꫯ����N��� ��� �:���;��q�������'O���'O��     ����f\�|9.^�.\�����x����  ��  �N��{h�����/��b|�[ߊ�z(N�<��[     ����㭷ފ���������t�R\�|9�n������YYYy��7 �{!p �u��Zl�}꺎s��Źs�b߾}q�ĉ8v�X�ݻ���     F���f\�v-�^�������o��V\�r��������c!p �u�  ��R�ox���8s�L�9s&<KKK�����R�s     ��X[[��7o�͛7�ƍq��ոv�Z\�~=�]�kkk�'���"���  �&p �����^�|��x��7�^�]�v���\������L8p �}�F    �����X__�[�n��������vȾ��7n܈����W��GJ��  �N�9  �Q��������{��^|�{ߋ����bjj*���SSS�o߾����ݻw���x���^     �����9G�9666""b0�����u]���f�����ǃ� ����3d���,�?�Qu]� h%�;  m�Tz�{��:VWWcuu�=���z���\���c����X��J_��W��ٳ�g    r;Dg�\p ���  �Qk.�o���/�hx�(��ݾ~   @+=)"r�!  �NU�  p���     ���\\\\(=  �M� @����싈��;      F�c�  ��	� h�~��z;     @��� ��� �*UU-��      0
RJ���   �&p �m\p     h�#�  ��	� h�;     @3�  ��� ��Y,=      `D/=   �M� @��     �1}�����G  �;	� h���      Fŭ[����   �$p �m\p     hH����  ���  ����̾��*�     `T���  ��� �������      0J\p �m�  �FJi��     �s��   x'�;  ��RZ*�     `ĸ� @�� h���      F̱�H�G  �mw  �d��      ����ѣӥG  �mw  Z#�t��     ��Tz   �&p �5rγ�7      ����  �6�;  m�;     @��  ��� �6�     4��룥7  �mw  Z�رc�1Uz     ��I)�� @k� h������      F�� ��� �
u])�     `D-�   �	� h�^��;     @.� �w  Z!��;     @�=����#   B� @{��     PH]׮� �
w  Z!�,p     (dssS� @+� h��ґ�      FUJI� @+� h�     
� �w  ��w     �r�  ��� ��p�     ��;  � p ���8Tz     �� �
w  �;r��LD�K�      aK�  @�� �v�-=      `�훞��*=  �  ������      0�v�ڵXz  � (.��;     @aUU	� (N� @q9g�     �[*=   �  WU��      �� @qw  ��9.�     �8Zz   � h�;     @y�  �� �6�.=      `��gKo   �;  m p     (,�t��  � �w     ��\p �8�;  mp��       bbfff_�  �6�;  E9rd2"�K�       b||�H�  �6�;  E�z���      ����gKo  `�	� (*�$p     h����  %p �4�;     @KTU%p �(�;  E�u-p     h���l�  �6�;  E����      ���  %p �4�     Z"�|��  F�� ��\p     h����  %p �����      ��;  E	� (��k�;     @{�� @Qw  �r�     �U<�裻K�  `t	� (M�     ���͛�K�  `t	� (M�     �"9���  ]w  J�     �H]�GJo  `t	� (�駟�{K�      �/�z=� (F� @1+++��     �L��w  �� PL���     ���  #p �����      -�Rr� �b�  �$p     h����  #p �����     �}\p ��;  %	�     ��w  �� PL��@�      ����H�G  0��  �R�*�     �16==���  F�� �br�w     �;Tz  �I� @1.�     �SUUӥ7  0��  �s�_z      ?*�$p ��;  ��]p     h'�;  E� (&�$p     h!� (E� @Iw     �v� P�� ���      -T׵� �"�  �ҋ���#      �Q)%�;  E� (�رc�""��     �	� (B� @�n��_z      �I� @w  ���zS�7      ��  !p �����      �%p ��;  E�     Z�PD��#  =w  ���J�     �^c333{K�  `�� ("�,p     h������  =w  �p�     ��RJw  'p ��     �M� @	w  �H)	�     �M� @��  �;     @��u-p �qw  ��     �ޡ�  =w  �H)	�     Z,�t��  F�� �R��      �]M�  ��� P��      �&p �qw  J�     ��� ��	� (E�     �b)%�;  �� PB{K�      ����  ��� и����J�      ��  ��� и��I��     �o��G�]z  �E� @�rΓ�7      ��]�vm��  F�� ��	�     �allL� @��  4N�     ���@� @��  � p     耪����  �h� �8�     ���k� h�� ��      �s� �(�;  %�     : ����  F�� ��UU%p     � � h�� ��      �R� �(�;  ��9�     �A� @��  � p     ���  0Z�  � p     �� h�� ��      �R� �(�;  %�     : 缿�  F�� ����      ��;  M� и���      �s� �(�;  �s�     �3��  �h� P��     ��'J�  `t� (A�     ����S�7  0:�  � p     �]�v	� h�� ��U1^z      [3���  ��� ШÇTz      [SU��  4F� @�RJ��7      �u9g�;  �� �(�;     @������  ��� Ш��1�;     @��� @��  4*�,p     萔�� ��� h��     �C\p �Iw  �;     @�� h�� ���)=      ��K)�/� ��!p �i�      pO��^  #p �Q)���      �'w  #p �iw     �n� ��;  ���Z�     �-w  #p �Q)%�;     @����  4F� @��      �s� ��;  M�     t�� ��� hTJI�     �-{""� �h� Ш���      �R-..�;  !p �Q)���      �7u]O��  �h� �4�=      :&�,p �w  �&p     ��;  M� �4�;     @�� h�� �F���      ������  �h� Ш���     �{\p �w  �6Qz       �&�,p �w  ��;     @�� h�� ��	�     �G� @#�  4M�     �=w  !p �iw     ���9� h�� �&��      �"p �w  3333Qz      ���*�;  �� И~�?^z      �.�,p �w  SU��     ���  4B� @c�      �%p �w  �$p     �&�;  �� И��M�;     @7	� h�� �Ƥ�&Jo      `[�  4B� @cRJ.�     t�� �F� h��     ����  �h� И����      ؖ=�  0�  4��k�;     @7�N�>=Vz  >�;  �I)�*�     ��y�W�Ko  ��'p �1w     �����w  �N� @cr�~l%     @GUU%p `��  4�w     ��J)M��  ��O� @c��     tTJ�w  �N� @c\p     �4�;  C'p �19��      ؞�` p `��  4�w     ��J)	� :�;  �I)��     �]w  �N� @cr�.�     t��  4A� @��      �%p `��  4�w     ���Z� ��	� hLJI�     �Q)%�;  C'p �1)���      �6�;  C'p �19g�     �K� ��	� h��     ��RJ�Ko  ��'p �Iw  ��ha    IDAT   �����w  �N� @��      �R�(� ��� ����Jo      `�\p `��  4&��;     @w	� :�;  M�     t�� ��� �$�;     @G���  �� �&	�     :*�,p `��  4i��       �M� ��	� h��      �%p `��  4I�     �]w  �N� @��      �%p `��  4i��       �M� ��	� hJ?|�	     �ew  ��_z��Z^^���z����ґ�����@UU�1Q����R*��-�@D��Ǜ)�A�y="�kq3���s^����N (f}}�������g      �MUUM-//���; �aUJi<�<����kWD�RJ�rν��w5"���=�9窪V#�f]�k?��r���^�wq0\��_��K�w�"��}�K_ZJ)=]����HD����"b|0DDD�9""RJ?�1�u���V?       �v9�^���Z 5��~x�c�1��v����v㻼���"���nD�\U՟���W~�W�7�yT�w�o��o���깈x6">�r��  �w�      �)�9g��Q2O�������:""���W#�ň��񍺮������_����6����Ω�ҧ"��\D�� �j���     ���ATUUz @������^UU,//�DğD���9��~��^,����[�{��{677&��3񩈘+�	 �K�d     ��s� �f#��"��RJ���|!"��s�r����������:A�~��[�����?�s��`0�k)��қ  ��v     t�`0(= �K�"�SJ�86�����R�������7~�7^/=�������9��9����l���G  ;@�     �}�� `��"�r�?���������?�9��]�v��_��_�Rz\���#"眖��2��Ku]����(�	 �A�s����}�eg]�߳ϝ	I�$Pe����ش�VQ���"(-��ը���ҁ{�3#Jr@��9�d���j��"�6`*��,|c�l�4�,�$& M($s3q^�~�G��I2/����}���]k��������^��]:      [d�; �XT9��F�s�9r�`0�����f�d3�������������L)}M�<  ��4     ���� 0vgG�����8~�����ѣ���׼����2��<��녈�ќ�9��  ��     ��w ���g)���:�+���[��:����ҡ�6S����_\U՞�h�҈�� 0K�     �Ϟ ���~�h4z�`0xw]�����sK�\M���{����)�+"��J� �E�y      ��= �Fu"�������`����~fqq��5iS]pEľ�����
�       �V��t �Y�����}0�^J銥����4)SYp_�Rzm������\  �0��      �g� ��/�9�`0��N��waa�s�C��T�{������WD��s��� �?��	     �~�Ѩt  "���l4����:�������C�KU:�������*"���v �m&�\:      [d� ��rnJ�ʺ�?9_T:̸�~����r4��/+� �S��	     �~&� lKO�9�w0�nJ駖����t��h���s���F���v �mN�     ����  lk/�9|8�"�J�٬V��������9�_���K� ��rΥ#      �E&� l{��i8~`8>�t��h]�}8^RUխ���Y  X?�<      �Ϟ @k<?����`𓥃l�\� 뵲�����9����Y  �8�     ��w �V9?"���F?�w�ރ��G+&���:��M�� �R�y      ��= �VzY�ӹy����*d=�}�}m,��qQ�,  l��N     ���� �Z�����u�����N�����ڵ�@�����  �u9��      آ�hT:  �����~0����՟��zGJ:�m9���o|����@� `z��     �~�|  ��ڵ돮��'�r2ۮ������s�Λ#�y��  0>&�     ��	�  �!���cǎ}���?�t�G�V�~���)�E�SJg `�L�      h?{>  S�))�?ۿ�w�r�mSp����>����8�t  ��w     ��3� `��WU��~����A���~��;���xL�,  L�i      �g� `*�L)�z���]:H�6(��=)�k�C  &�b'     @��� �ZUJ���`pE� %/����F�J�  4#�\:      [4�JG  `�^7�*�X�}0�.�T�? ���     �~�|  �_�y�`0(6ļH�����"���z  �c�;     @��� 03��u��x����2�te�� �,�<      ��P# �ّR�r0,5}�F��ಔҵM^ ���b'     @�;v�t  ��?��+�����6yM  �w     ���� 0sRD��.x#)��߿���;#����  �~,v     ��= ��ԩ��7����k�b/����\PU�{"b~�� `���	     �~u]��  @9�s������I_k�����]�N���I^        �<C�  f�W��ͽweee�$/2��{�9u:�_��gL�  ���N        h�g��ͽ#�&u��������dR� �]�     گ���  (,����p�<��O������-��I�        (C� �5o�9���ྲ�rAD�fD̍��  ��	�      �g� �5U��k���x�'��zU��y{J���</  �g�     ����  p\J��UU���덵�>֓���w#���<'        �=�u]:  �HJ�[�=�ܥq�sl��`����q� ��b�     @��� ��RJoX뒏�X
��]w�Y����9�� 0},v       �T�����3�����~�ȑ+"�_��\        ��T�u�  lO_}����8N���p8|fD,�!  S�w     ��Sp �TRJ{����z�-ܯ���9�GĎ� `�)�       �T���_�����-�R�}uu�?F�3�r        �Lp ��y���Wn��.�_s�5O�9_��� 0;Lp     h?w  ��u+++l��M܏;֏��7{<  �E�     ����  ����z�f�T�}���ύ���E          �N)���:����{UU�#"m�X        ���. �vHUU]�s�p�|���`��ƍ �l��	     �~�|  ؀��n�m��~�7t"��7z           fKJ�M�^on#�l��~�w�<".�P*  ���s�      l�	�  l�����d#���6�}�F @��;     �4Pp `~f#S��]p��;~0"���H  �<w     ���� �&<u׮]�a�_^W�}mz��l:  3/�T:      [�� �f�_��I?�u�o����o)  3��*     �O� �Mz�Z'���UpO)-n-        0�� ؤ��|���p�����-� `�Y�     ��}  ،�ҿ���g쥟���s�=�H  �2�      ���  �UU���-����\/["  f��N     ��P�u�  �T������)���>77���1�T        @k)� �;:�Ώ���,��S���          ��X�9���S�8���D        Z�w  �����N��)�u]�|2y           �a�쪟�����/�X           f�K����O��I�v�zaD�h$        �urΥ#  �~�u]��d����s�d�y           �a'�?�����Ή�N<           3)��=�~��G���������1�H*           fN������G����{J�I        �Nιt  �DUU/x�{�|#���<  lUJ�t        `�9� ���b��
����9���          �z�`0���xX�����l           f�N|Q=��om.           �,��-'�~��~�7tRJ��|$  fAJ�t        `�y�7��9�⡂�w��8�H$           f�y��v�3���N����          `���겟Xp��Y           �a)������g� ��H)��      ��KG  `�\|�UD�u�]w^D��bq           �UO�ꪫΏX+�>|��0R          ����;w>+b���*          �6��6b���R��e�  0�R��      �i�s. ����k�����f `�)�        ��Rzz�?LpWp          ���+++�"�+
� `�yT%        p_y�uםW���=�t        �6 `R>�UU]�O* ��R*        �ƪ�zR�Rzb�         @;�� ���u��*"�          (�UD\P:           �-���*"�Q�   L��R�        �6�s~\�+        h��s�  L����;           ��㪈xl�           ̼�V9�sK�  `���JG      `��  0A�V)��S  0�,t        g��J)�,� ���        ���*�l�;        �. 0A;���+� ��g�     `:�� `�vTq�t
  �_UU�#      0
�  L��*�t�t
  ���N     ��`� �	:Z圏�N ����	        ���*�l�;  ��     0��  0AG���j�  L?�      ӡ���  �^�W��)  �~
�      ���  ��R�b_, ��g�     `:�� `Rr�_4� �FX�        N'���*"�_�   L?w     ��`� �II)}���ϖ ����	     0��  0)9绪���t  ���N     ��`� �	��J)�Y:  ��B'     �t�� �����4� �FX�        N'�|Wu����J `�)�     L�>  L�h4��ڷo߽�w��  0�,t     �_Jɾ  ��}���[���T�(  L=�      �g� �I�9*"���H)�U�8  L;��        ���W9�O�� ������_     `[3� �	�ˈ�����Y  �v;     �Ϟ  ��s�h�Z���ѣ�DD.� ��f�     ����  0!ynn�ck�}����.	 ��f�     ����  0!���𥈵���[
� `X�        N����P�=���2Y        �60� �	���?N,��L  fAUUg�      ۚ=  &�.�Cw���w��"�`�8  L=�<      �Ϟ  ������_<Tp��z�RJ.�	 �ig�     ����  0�����g����<  ���        �I�ɉ/Vp����� ��Pp     h?{>  �[J��'�~X�}yy�/"�F 0,v     ��=  ��s������7VpO)���F# 0��:�      ��� �����:�9Y����        ���;  �s~�#�{T�}uu��#��F 03:�N�      l��� 0.)�C9�?x�������z��w  ��b'     @�j ���߻������j�k�y  �1
�      �R* �)�R:ig��-�����E��D 0S�     ��w  �!�t����?�g'm�z�C��&�
 ����     �~&� 0u]�{yy���}vʖQJ魓� ��Qp     h?{>  ��)�ꧼ�\\\�����$�  0{L�      h?w  ��o�����Mp�)��O&  ���锎      �)� 0oI)�S}x�;Δ�["���# 0sLp     h?w  ��hUUo=�N{ǹ��xWD�8�H  �$�     �O� �-�����)��3�|���  0�,v     ���F  lEJ���3�����?>�D  ̬�R�      l�=  ��楥�������Ѽf�a  �q�y      ���� ���|i]w�^x��-� `���     �~
�  lҧWWWߵ�/����K/��V��	 �Yf�     ����  �9�_��z����u�q��Ͽ#"n�l(  f��N     ����^  6*�t����������[F�_~�є�U�� ��Sp     h�N�S:  ���^�wd�_�P���O~�/�?��L  �:w     ��3� ������[6r��ZF�^z�(�t��2 ����<     ��P#  6"����/���F���g��}wD|x�� 0��     گ�锎  @{�����=h�R�/"�&� `F)�     ���  �)G�rJiÝ�Mܻ��"�77s,  ��D     �v����� `���~c�s�a����z1"����  �=      �M� �u8�Rڳك7}ǹgϞ��9�a�� 0{Lp     h7w  �$�����Ż6{���8�;�k"��[9  ��w     �vSp �>>??�VN��;��/��hJ�#��V� �l��	     �n�{  8�c�c�_~����[��\ZZ�hJ�ꭞ ����tJG      `<� ��t����Փ��O*w��qeD|b� `zY�     h7�  8�������8�X
�w�>�s�ш��8y  ��O     �v���ԍ  �.Gs�?�����8N6�;���古�^7�� 0}Lp     h7w  N������q�l�w�|SD��8�	 ��0�     ��� x�]x�+�<�X�8{�^=�~8"�0�� 0Lp     h7�=  �����.����8O:�?�ܻw�9�E�X� �~&z      ��'� ��������{�O<������SJWN��  ��O     �v�� ���v���O�������Ɯ�oM��  ��O     �v��^  "�w����4��O�3���:���['u  �ł'     @���͕�  @Y��ܹ�R��&�0ڽ{�}�N�E��I^ �v0�     ����  ̴{�~��ݻ��E&>BsaaᶈxaD�?�k ����     �n�� 0�H)}��={>=�5r���vo����Q� `{��	     �n ̤QD�����MM\���Q�۽1"~,"rS� `{��J     �v�� 0srD��Z�����v�o�9���k �}X�     h7�=  3g_��}s�l�����|]����.  �UU㷟      ����\�  4��nw�-�0Z^^����ĵ (�D     �v�� 0r΃n����.6Bsyyy9"^_��  4ς'     @�yb/ �Lؿ��.��g�۽2缯d  ���     �^UUEJ�t  &(����v���P�O*���WRJ��Kg `��     ��^ �T�)�奥���ˋ�#"���)������  09Y	     �^
�  S�X��'�����Dl��{D���ү��^��� �dX�     h/{=  S��������_)�mSp��XZZ�ú��w�� ��Y�     h�����  �;���n����AN��
�{��e�ΝGćJg `��     ګ��]� �ͻ���|ݞ={n)䑶�]��ݻ�޹s�wD��Jg `|�     ��^ �������maa�s���̶}n��ݻG������)�AD�H\�    IDATU:  [c�     ����m� ��9�s�.//�b� ��-'��hyy���ƈ�t�,  l��V     ��aF  �R�#���۽�т�{DĞ={n9v�س#���Y  �<��      �e� @k�x���g,--�T:�z��A���7"�w8^�s�>"W:  ��     �^ss�� ��"b���t��hݟU.--�+"�6"��t  6F�     ����  �������m+�G�����vo_]]}~D�:"VK� `}<�     ��� Za5"^����M���]:�f���A�^���kWVV���t������ ��yl%     @{)� l{���v�����o�ݻ��q�`0xID\O*	 �S0�     ��� ��;#�U�n���A�ajF�n����է��E���y  x4��      �e� `{I)J)��F�����1�O���E���W_�ku]_?ST� h;��      �e� `����,,,�V:̸MU�����Ż"��~���RJWD�K#"� 0���     ���; ��������vo.dR���~�������K���3s�?��� 0�����     `�)� ����~vqq��K���h---�E<XtND��9�8"� hXUU�R��s�(      l��; @���{"b����M��4e&
�ǭ��}Ɂ�Z���r�?g�� 0K����hT:      �i�  �9����iaaᓥ�4m&�:>�:p������҈xUD\T8 �L���Sp     h!� &��9��r�Yg�e���w�S�L܏[XX�RD������9�����.��F�Y�� L-�      �d�; �D��߫���C�}���ե��3"�~>8p��c�����e���ʦ �.
�      �� 0V7G�;v����Y��~2�:am���Fį��D�Kr�/N)����� �"�      �d� `KF9���RzOD���vo/h�r�yk�8"��`0��ҋr���_V6 @;Y�     h'�<  ��������rο���|O�@m�s����=�x[�׫�9�g���=�������xlр  -��x(     @�ر�t ���K������СC��zu�Pm��	k�h����s��k��꺮����礔.���"�ܢA �!�=      ��> �����9�RU�MUU}�կ~�_��r�`m�s�~?��󶈈^�W���_u�ر����RJO�������'� �L2�     ��<� �AG#�o#�o"�orΟ��O���}��{����Jd�:
��������<⳹��?��ǎ{|J�	)�'�u��qVUU��9?&"Ύ��a
�vw,"��.�9?����D�h���	?D�߯� 3�ȑ#�O*�     ���9�N<8� fI'"��:�:᧳��s�{;"b5">Q #�s(�r�联���u�ň8\U�=9���??77w����{w��;V �LSp/`��sk?  3�.xgD|�      l�[��֟���?�K�  `�U�  0s(      �����P�  L?w  ����      �qw�}�}  &N� �F�-|     �ϑ�8V:  �O� ��=P:       f� �F(� Ш��Lp     h�C�  0� hT�Y�     �eRJ&� �w  �f�     �er��x  h��;  M3�     �eRJ�Jg  `6(� Ш���;     @˘� @S� h��O     ��1� �F(� ШN�c�;     @�b @#� h��W     ��=  �� @�Lp     h�C�  0� h��      �c� �F(� Ш��	�      �c�;  �Pp �Q9g�=      ��  �Pp �Q���w     ��Qp �
�  4j~~^�     �}� h��;  �:��-~     �ϡ�  �
�  4��[o=��9      �C�  h��;  %.      �1� �F(� P�	      -�s�� @#� (�(     @��� �
�  �`     �ERJ��3  0� (���      X?w  ��� @	�J      `������  �lPp ��     Z����7� �F(� P��;     @{�{���  �Pp ��C�      �n�"�. �٠� @	&|      ����  �
�  4.�d�;     @{��  ��Pp ��     �C� ��(� P�	�      �� @c� h\]�&�     �DJ�`�  �w  J0�     �%r�&� �w  J0�     �=� h��;  %��     �K  `v(� и��	�      -�R2� ��(� P��;     @K�u�� @c� (�P�       ��	�  4I� �ƥ�Lp     hw  �� @	&�     �DJ�`�  �w  ��tLp     h���Mp �1
�  4n׮]
�      -�RRp �1
�  4��[o=�J�      ��RJKg  `v(� Pʡ�      8���Lp �1
�  �r�       ���Ç� h��;  ���     �sssKg  `v(� P�	�      �_���~���!  �
�  �b�;  ��ۻ�9ӳ������n�7Yd��,k,Y���@H��D�!eI@BBd�a�r��d�'$�x�v������~� ��C���y��kg�]��޼���.   �w��ҲG  �>�  dq�     �w�  �^�  d�     ��N�   ֋� �,��      �J.� �Tw  ���     й�� �Tw  Rx3     �����  ��;  )�q���     ����;  K%p  ED�     :�Z��� ��"p  ��     ��5� X*�;  )�q�     t."�  ,�� �.�     L���  ��;  )�      �s� �e� �b�ϲ7      �r�5�;  K%p  ��      ������  �z� �b�;     @��qt� ��� ����w     ���� �R	� H�����2f�      ��Ο?�;  K%p  �XJ��=     �:���z�= ��"p  ӝ�      ����  ��;  �>�      �d  `�� ��;     @�"B� ��	� �$p     �Tk�v�  ֏� �Lw     �N��\p `��  d�     t*"\p `��  �i�	�     ��;  K'p  MD�     :w  �N� @�;     @�Zk��7  �~�  ����      <��  d� ��w     �~�� @�;  i�      ���w  �N� @�q�      ��A� ��	� H�;     @����ogo  `�� HSk�     tjcc�w  �N� @�Ǐ�     �Ԯ^��Y�  ֏� �4��̛�      }�[J9� ��� �f{{���Ҳw      �7�  ���  d:*���     �� H!p  ���      |�� �w  �d      ��  �� ��w     ��� H!p  ��     �?w  R� �&p     �� �w  �	�     �#p  �� �T�5�;     @gZkw  R� H�      ��;  )�  �r�     �?�8
� H!p  U�U�     ЙǏ� H!p  ��      �y|�֭;�#  XOw  R��(p     �˭RJ� �z� �j6�	�     �r3{   �K� @���#�;     @_�  �� ��_���     �/w  �� Hu���ǥ���;      �w  �� �+�      �� �F� @�      �� �F� @�      �� �F� @�֚�     �w  �� Hw     �N���  �� ��;     @'�  d� ��w     �~��(p  �� �t����      �֗����do  `}	� H�Zs�     ��.]z�= ��%p  ]�U�     Ё���� ��&p  ]k�V�      Ji����  �z� ��@      ���  �z� ��;     @�  �� ����X�     Ё֚� �Tw  �-�{���;      �]D� H%p ���      ������  �z� Ћ��      ��8�.� �J� @/�      �j�w  R	� ��~�      �u���)p  �� �.��\p     �������#  Xow  z!p     ��z;  ��  t��*p     H�Z� �N� @/�      �"b/{  � �BD�go      Xs.� �N� @/\p     H�Z� �N� @/�      �"B� @:�;  ]��
�     	� �� �.\�z�v)�({     ���q/{  � �E+��&{     ������ @:�;  =��=      `]mnn
� H'p �'w     �/_�|�=  �  �d?{      ��r� �.� ��      	Zkw  � p �'w     �!p �w  z"p     ȱ�=   J� ��;     @�֚�  tA� @O��      ���� ��;  ���)     @�k�  ��;  9::�     $h�ͳ7  @)w  �"p     H0���  tA� @7�ŽR���      k�p�X��  �� �+�      Kۥ���  J� ��;     �r]�   �� ��;     �����  �sw  ��Z�     ,��  tC� @W"B�     �\.� ��;  ]�     ,�� �n� ��8�w     �庖=   >'p �+���     `��� @7�  te�     ��p�X��  �� Е�
�     �g^Ji�#  �sw  �r�ƍ���{�;      �AD̳7  ���  ��z�      �u�Z� ��;  =Zd      Xײ  ���  �h/{      ��p� ��� �Nk�w     ��� ��;  ݉�;     �r\�   O� �#�;     ��� @W�  t��&p     8{����F�  x�� ��D��     ���K)-{  <M� @wj�w     �3��  �,�;  ��q;{     ��k�meo  �g	� ������Rʭ�      +���  �,�;  ��      g("�  tG� @�Zkw     �3�Z���  �%p �Wײ      ��Z��  tG� @�j���      V��|>��  �� Х��<{     �
�*���#  �Yw  z%p     8;�f  ��� Ыk�      V�� �.	� �����     ��� �� �.-�{����;      VQk�r�  x�;  ݊�y�     �UTk�u�  x�;  �j�	�     ����� �.	� �ٵ�      +ho�N�  x�;  =��      ��~�=   ^d�=   ^b�Z+��� /t���rpp�=���ѣ2�c�    �Rk-E� @��  t��6?<<�]������׳g@��Ey��a�    ��/}��R>��  /R�  ���֮eo      X5�V� �� �n	�     N�� �n	� ������Z���      �""������  �"w  z��      �
"��Rv����do �� е����      �
��d�  ��� е��V�     �U�����  �2w  �VkuE     �<��.p �kw  ����     `DD��;  ]� е�l�MV     �S�$p�8{  ��� ��=z��'_�	     �[���������  /#p �k7nܸ�;      V�/J)-{  ��� �)pI     �-DD��^��  �"p �{�֭�      S�����  �*w  ��Z�${     ���ZK)���  �*w  �7�k"      o��Zj�>s �{w  �7�k"      o!"������;  �U�  tocc�W�=     `�"�J)c�  x�;  ݻr��^��a�     ������  pw  ��E�N�     �)�����G�;  �$�  L�V�      �)� 0%w  &�����      Smss�g�;  �$�  L�0���      0E����u;{  ��� ���yDdo      ��Z�G�  ��  L�0��     ���(�0|��  NJ� �$���Ok���w      LI����x1{  ��� ��8��ne�      ��Zk���d�  ��� 0�q�     �)�����ٹ��  NJ� �d��Q�     �)q� ��� 0%��     �$"��Z��  ^�: �ɨ�
�     N���*�w  ��P 0��엵�1{     ��Z˹s�~��  ^�� �����zW�w      LA�u�ʕ+��;  �u� ��a~��     `
�a�Q�  x]w  �惈��      еZk)��w�  x]w  &����'o�     ���w  &G �������     ��axx���w  ��R 0)����Z���      =����ҥK��w  ��� 05���Q�     �^ED��~/{  �	�;  �DD�     �.�P"���;  �M� ����Ok�(     �<�0���d�  �7�
 `���     <_D\��緲w  ��P 09���G�0<��     Л�(����  oJ� ��\�x�q����      ����R���  oJ� �$E�k�8     �ak����  oJ �$��~$p     �]�0|o>�?��  oJ �$���'_�	     @)��g'���  oC� �$]�v�r�u?{     @/�a(�n�  xw  ��E�k�H     PJ)�ֽ���f�  ��� `���     �����RJ��  oC �d�����0d�      H7��J)�;�;  �m	� ������#� {     @�Z��W����w  ��� 0e���Z=�     ��Z�a�ǋ/>��  oK	 ��E�{�0d�      H�䳒�d�  �� p `�Zk��;     ��f���Rʻ�;  �4(�  ����݋�0lg�      �Pk-�͝����[  �4� ��VJ��'_�	     �Vf�Y���g�  ��"p `���     XG�0�r{{��;  �� X��� {     �2=������o� �� p `�vvv�R��V��     ��������7�w  �iR  �*�9�Ͳ7      ,E����wׯ__do ��$p `%Dķ�a���     `f��8���d�  ��&p `%���܏����#.     ��"��f�o���}��  N�� ��Qk��l6˞     p�666Jk�w  �Y� �2���{��̥     `eED���������-  p�  ���Z�+W�    �U���qw�?��  gE� �J�����l6�u�     ����c�  �IDAT6C��/���v�  8+w  V�q��/�a��     p�Ν;�㝝����  gI� ��������s��-{     �i����Mk�OJ)��[  �,	� XE-"�l6���     �f��݈���b�i�  8kw  V����s���iq�     ���l�����{{{?��  � p `e���~kss�K)7��      ��Z��l������������{  `Yf�  �,-�*�|�TJ���X=<x��͛���:�[Jy�=  ���ZJN�Ν���͎�����f��8����儍Gk���x*��g�M�^��~ "�k��[��Q)�=��G���q)�w��a~�5#�?���Xk�=����s�  �v���R�y�L    IEND�B`�PK
     E"BY'�Y��  �  /   images/4bf63cb1-3675-4452-8ab6-1403298522d5.png�PNG

   IHDR   d      X�   	pHYs  �  ��iTS   tEXtSoftware www.inkscape.org��<  SIDATx���KA�_�&�Ҕj�PZL-1����?�7O=x��[�ދ'�{�xl=x#"�P"�ɖ�T�[b�&���ݢv��xa��o�;o�f&
I ��ё��v��F��5�M������Yj�ۧ�����ZZZ��v�����$��\�v�T�)�Q�Z���?�;r�V�B�x�1E����� &M6���������FM�0��UUu���[�;<<$��K�Z�L���B�@�LF/_7Ft�o}<YB��.��Ȉ�8��p�\�b�hY��|>D�A=�\����l!�>����=�����y�ϐ!v�[V�������ѓ�=��a��ò���;�\��)�mr.�&�277'�A,C�d�����ƉpF��F)�uI�
f�`���(_���X��N�ǐ�v�����4�q$����"�q�	T���.�[�$�F���E��:MdW���a��n��4�'�b�to���f�����<��.�1L� �=�%n ���r�F�I�wQR�V!��{�G"[��Zbh_+���Ol3$����%��;�'���������(Ϥ'�0�j�����U�99��Xf{Ƕk�Cv�8����
�����v� ;;;����W��t)�x�D�ֱLmll ��PX���ښ^����.�P̂(p$mP!��/eqqQh��!Fk�\��jX� 8.1�d�"��{�n��Il�~�&#��r���>�t�z�JE���>��-��ޞ^�n�a<I��+nDE#E������O�[V�0��T*u�pZl�k'���UV�R1�n�y0q�<��>���$���I�"�t}�4���������J�u�    IEND�B`�PK
     E"BY�}���) �) /   images/146a6d58-0553-42c9-b8c7-03425202d69a.png�PNG

   IHDR  �  A   s���   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<    IDATx���y�e�?�Ϸ���{rL�쮞�8���D@DQ��\\����Sw�׽���o�kw]�]uՠ�r� �A#�1�LWu�a�=�g}�L6��]�OU���z�B���Lz�SϷ�GTDDDDDDDd�e: ��E:Q��E :Q��E :Q��E@�t ��U�V�4�g��Ed���S���e�Q�9"�c:#=���Dd���pPD�=���f�7.ܴaÆ��KT�t��ŋ����z	�� �� Kͦ"""""�4l��U�n����j�t�N��NG���ۯ�oUճ ��-�����:�U���ܞJ���f:PR���!�����{�l8E�/"?Wիj���ر��@IN(���}�OE��ƁDDDDD45�E�|�\.o2&	X�;������ϱ,�S ^d:Ŗ�F����R���t�8cA�@���? x��,DDDDD�
�Z��/�T*�1&�X�;H�X\��_�:�Y�����(� �\��>�gԧ���^�:�w�ޏ�[ Y�q������3TT�/<ϻ�t��`AO8�qN ��sMg!""""����j�z�Ν;��u,�	V(.�/�6�������:�oU�|��6$�X�h���s������Lg!"""""U�	�u�`:HT��'L�X\��78�t"""""�#����~XU[��Dz�������� V��BDDDDD4�k\��� Qb�@�(�%���s"""""��7�iժU=��D	W��X,�DUo0�t"""""�ixز���6$
X�c�X,�V՟8�t"""�NcYl�>�;�:[Uq�u�x��>�t_��xŶm��bz���yǲ��pLg!"""�T�t]]]�P�g*�~�7&����<8��&��4�<�{��6M1�=����q�e��9���0�E��?."��yc��������ؿ��u��?��DD�H"�l6�T*e:J,} ��r��oz��^����Y�cHDR�B� g��B�3�b;ٯ����'{��~�|����0�9E�n {�KU����"rPU� v�H����"r@U�m� ���e%�aU�����y�nذ��r�ʬ����HVUs�V+e��< h6�� �eY�T5 '"Y =�:ϲ���:ODzTu>�y�Ke.F��[K�L]]]�cP��=i0������ED��\.�������P�X�������b�eq&%s���h�n&�f��h�V��n9�� �� ���N١��Dd����}���I��{Dd����Ӂ�AD��K�kYֱ�T�8U=���_4��ǉ�  ��Mf&cYr�,�&��z�Z�t��j�Ꙟ���tX�c�X,�JUoB�ض��ol3-�S-Γ�7�<����a�Z-�Q(�|�o@e����eYe [���J�2d0cb���X�bI��X�`Y�U-���(���lR�"r��t�v�y93��u�2��X�c�X,.WՇ0�J�x�T
�܄S�D��9M�6 �l�YU7��&U��/_�u������}}}��j���+,�Z��+D��
����&���m�l����	)�  U��R���ӞGgA��b�x����t�vbI'��*�*:��	U��eY� lR�͍Fc3��I��+W.h6����٪�l����f�Q�uuu!�ɘ�A	��r>FD�W.��f:G;���D�X|��^k:�	,��.�f�Z-���Ь40�
���<����e=������7�3�����_�l6���}��| '�� ,7�����m�r9>RG�Kb9��s;iԝ=��|���ZDV��b
K:��V��^���A��xTD�}�a���|���q�f�q��"��|�?AD���yw:
�FAKp9 ��������.,�1�]�G��S|�G�Z�Fp�T�k � xTU�G:�.<�5�w�I"r�����<�Nth9���l$����E��r���� ���q+W�\�l6�-�%���!��:E#e� ���~ٲe�*NQ�8�B��O�,�U=EDN�, liȲ,d�Yضm:
�P�]���u��M�h�+
�&"2�#JX�i�x|Z����=���U��t:����@�t0��X�jUO��\����� ^�Xӹ�}2��c�ii4�V;�۞���y��s��=?��%�Fc  ��X�i�x|Z,��C������Ǟ��2�(L�bq���/�3D�_U׀�t���t��N,�~��+L�z�9��O >n:GT���t���Z��f�i:
Mn+�{�#"�������7�:��ŋ�f2�5"r&��bd���p,
�c��tp9 ������t�0��GToo�1���g:K����T4�MT�U��G�+"?�˲�ڲeˀ�@DQ�z����ݻ׈ș�����5Cbض�l6˲LG���r>�G��c:D�X�#�q�?�%�9�%�ƣ���jh4�OX�<	�'������!�=I9�s2�����1��>�p,��l6�t:m:E ��!���++�J�t����G��8�Xc:G\��ӑZ���*|�7��� ���Z��T*�'L"J�R��ޱc�i��RD���5n��T*�l6���:��ө�<����aaA��B��l���q��DiL�;E>�� �����˖-��ǝ��x���t�T˲�p6�~әh�,�BWWR���(�f,�G�[�u�c:DXX�#�X,~FU?i:G��w6��Q�Vy|��T�f˲n�}�6�Nm+V�X���kU�� �O��^�t�����r����a`A� �q� �5�#��ͫ3�����ܯ����R�<��?�(���|���ܲ�׏v�t&�� ���8����[���z�OU�r���u?j:DX�#&��?ײ��M�;����U�����"ru�\�j:����x��� "��Kp���d2���2�B0�rnYR�����' �*|�G��B�^�mYW��=�{��a`A��b��AU�w�9��%=��j��p��^_��n޹s�~Ӂ��}�Y���X�u����ә�Y��\.���d&�|6{4���Xn�+"�$.��GL�X\����˲�� 8T�Z�Vh�%=�x|Z�Tu��|_UP�T�W��}�&�����ͯ�j��VU}-x�[dtuu!�ɘ�A�4�r�ｪ�^��^���ux���m:D�X�#DD�P(l��t� �R�R�l۞�$>j�<��di�Z�y�\kY���r�g|���!��w[���,k����Z�� 9Ɋ�1 �������f,�:����sEd�Q�a �џ� p @������.��j�v�}��ڵm۶��O���+Wf����e�AU��%�3u�T*���.����t˹eY�f���E�l61<<���W\׽�t����GHoo�|��`:�l���V��Z��3�,��P���xw7�6�ڲ��>h:����bG��±���wU�� �)�=�b�DUU���U��˲|��T*[;y�DDR�B�ly������M�l6�t����t˹����;��11+�]�}��AcA��B�p��|�t��rgѱ栾FY���j�Z�����*����߫T*�C�!"�dɒE]]]�|�_$"�Tu��.�������=��M#+��x�y��]���r��l��|�hY?#7d��x�3)��lvFϛ��� ?�J��EةbA��b��W����s̔m���r�~3�.^*�B6��7��P�C�Ѭ�p���Woݺ�FU��dٲe�R��R Y��KG��h��K ,���6k����eY�����<�nl��f�q����g۶�U} >$�F�(r4;3)��ڽhh('��	�r9�ȇcA��q�	�ݦs̄eY�������w&U���p,�9DT�"����6n�Ȼ	���7�^�; ��Z�e �"�@�R  K ��hixLU)"��"�p�K{oo�1��+"��� �M�M��M3���;wn[~/U�}�v�u`:D�X�#�q���1�c�Ds��	�â^����J����{=
�O�1��"�t:}ͦM���D3�z������-�"r<��c��X`�ٔ��� �GUf�������6*,�����"r!���<��ǱE�L�y�V����l���fBU?�y�gL�z�8����9�+�˵e|*�Q���QUT���3��A _O�R_�b:�N�P�UD^i:�$���Ƚ�V�����&mFD�|>�2˲ޫ�o�X��ZM'sf3:gΜ��d�Æq"�r���s�="Fw@�ݡζm���=���Z-��,���l6Q�V�j>uU �cY�������U�
���ȿ��A�� �(��}߿=��ܓ���/^<7�ɼMD.p&8۶��f��n�l
��`�ܹ'�������Q�6��u�7�$�}6�)�9��]��c�ذ�%ݼj��F#v��Ly�U���g�R���0��K�.N�� ��D�_��=������}wRV����� .��p�����B&�}��e���W<�St�r]�e�C�="���cYV�t��j�Fc�:�!�N#��iA���Ӧl��~���=b:��X,^���Z����CI*�W���۷�-�� /W��	<�LAL	��V��s�"��r��o:G�X�#��������jCw���Q�%��j�����Q���[�u����n�a�}�y���A�6$"����|߿'��q�gx�����,1�'Ix[�����}\]�}��AbA��q���t��h�N�c����k�����}T�U�6���}��r�R��t2c��ՙ�{�np��,� �#"���-q�%~��ՙ={��ID>�e��$	�c^��Ҙq��y��\�Mԩ&,�Q,_��?5�c:L=�t���P7�`IO���%�& W���5>[N �8ο����L��ݲ��������n���q� �] ڳcm�Y��l6۶MG������,s�����l��u݅�C�="XЧ.�������R�����W*���;�X,�Q��M砎��0Fw�_�l�]�ׯ��Ν��,�Ȧr��p�D05%�A��1���)Ǭ���ǂ���ñ�#�oR1W��g]����0]��<
��9�� p'��}߿�R��b[��/_�r˲>���r�����	�݋c19e'q��AЌ��y���9��Ē>3��j���E�m���{�պ�c�4E�p���q�8�9�e�q��Y]�!������G��np���� �F>��chh�ǱMC؋�F�m���5��@Dx����q\A�?jc�f��O_�����0W���C �#�J]�[��b��\U� ��EQ1�Ǫz�y��4�e˖-J�R��~Ǚ�W�m#��²,�Q"�]��l�t:�� �;m'�ˡ�j�ډ[AgA�Sݶm��?��v}H�1��$K�Ԩ*��:�O� n�O���e:ŗ�87x��D�x���e�P.���^�|�۶�T�c V��W�v>�'"����fI�����P௛��J��.�,�S}�H����h�6��۳qjXSŒ>�V��j�ʑ%�p���]�\^o:�_�X|��~�t�ɨ�v���j�[w��q�t�#�>��z˲.p��<q�J���fy�({�ض�\.��A;����,R����Y�'Ƃ&z6�����Q���(��Ȓ�L�z�S��T�_��C��8N�� zLg!����ܧ����m�Ry�t�#�������� ^n(7-G�Ner�s˲���hI�M�Hww��6dA�zD�.��H���J��9sB����Y��W� � |ݶ�˶l���0�L�B�k"��s�¯�Ȳ��6
?z������aZ�&1;q5=
G��r�\ ;�7�MT���WΏ��}b,���������i�T�qoL��@��}�X�y|�m"��z�~Ŷm��C�����J��o5��( � ܨ��7�����|���ٶ�I �'MY�%1.�P���d��dft��>j�Z�;�O��<��X�#"*�VI����:����4� �/���R����:��X�B� o:Q�����F���m۶�0h�ʕ+���� \�6%"rh5=�~m�N�'�Y��h�Zh6���snYr�ܸٱ�O�="�TЁ��� u�C�:��w��y��T�+<*�L(
�OD��t��D��z����T*�d�B�P��� ���,q���آ\�'"�m�Й�"U�����P�t��.�,�cA����1���3Z)M���d23��n4���y��SJz�Z�.k� �����F��2%V�P8ID2���M��"��f�y�֭[7d�ҥ����� ���>%]]]�d2�c*.�ܤ�V�ǰ�O�="�ZЁ��t`�(��Q��F�}�G��@�ٌM1?\&�I�XW��Ą�����r_۸qc4v(���8ί �6��Ȁ� n�,�����{L���E˲>�" <|IZMg9��tueA�zDD�����Z�u�C��Q�$|&����1���Y _��y>�wL�R�
�O��gL� 2IU���u�e]].��m��X�|y�m��}�frtuu!�������Mw*􉱠GD�:��#�S����9�w ��e2�ܴi�^�aƳbŊe�V�r �X��Lg��]� �%)�`���DY_�b��V�u)�?�g�P\�cc9��m����֯aA���Ӕe���=O�(��>��z���vR9�YU]��Q-�"�r�#�V�	 ����R)��4m�J��n�9�"�����w�P(����덷l�2��%�e�PU�k���Q�����P�N�a9��m���b�X�iZ���G��Z�ǎ׋c�j �@���y�.Ӂ�S,�,
�<�������m��qC�Ȝo�@Q������M�yޛT�4 m������8�k�r>�T*���4������+c�a�[Io48x�`��nD���:y�뺗��[1h<+V�X�8�U�z'��LD��q�ڛ�L�d2�02�ADOw��M==����y/�6 �1�#��Vӣz��r>�t:͕���ӌd2��8Zl6�P��t7; ���K�����ry��0�9�8�D��3�{G}�F�9��FUo�@u]���V����3E���G�6�e9�\*��B]�X�i�:���وrIo6��{lʪ�^��N-�ˑ~~�q��
����q��pԽ�p̝��m�j:�Um��{����p)�H�ob���V�ahh(�ް�O.�� ��q�=d,�4+c#.��:�z��j�j:��T�Uwª�n ��R��x�wU����q:�s�x�t=G�;K*��	��':�788���G�T*C��^��� |@4�j�Z2���r>����)|,�4ku�\�шDIo�Z8x�`'�� pe��x�뺗��?""�B�B�<�x1&g�G�;���@UD~h:Q��b:�D<����G|�_�.�y�fl5�������hk{��S �Y��L��z��1����\׽d۶m;L����8'
����7 �K��cǎ?�u(T���3E��Ff�}"�J�!�u_���0�'j��&<ض��Z���$�9t���S`x���L�t��144�g�""����u�s\��h:�D��|��8� ��ڪ��u���� �7��ڤ��!�������<�G�3�'JƎ}{۱�z�W6��e�6W�'�h4�V���z�O�,s��ŢE�n�<��y&����`Y�c �#c�A� ����ɧ�M��t�X�y�.�!�kÆu�u�`��sU�k ?�6a�r>�l6�rn:ζm̙3�+�{w�NY5�f�X�p����yg�q�<ә��8N�q��[�u�ސ��$��w���g�}<[�ly����>�~��<Q���_ϰ�O.��"��}~SX�)�eq�}a��F�����D����i,\�===�m{����d��)�Ji�q.�[ ok����_����z?2��x�s����f�R�����U�� b7��&Y�'���X�cA�а�O.Ȓޮg�L�J�    IDAT�?.<�7��@�q�����o��s ����o�QիD$����6RU_Uי�AdоE�%f�YU}��J��/�� $���M��86������J��4t
�eY�3g,�_j�	����֮]OM���±�;�/)�J�mW��nw�eY �7��B��1��Om`Y�ܩ�ݱ~��ĝ�y����r��"�R �2�'Jj�������r>1A6�=|*�bk�ЍݑcI�lJ�L�Qŉm�8�c�`���~�0�Lq�u���}@������˟g:��\.?  �'�EDn3�!L�r�n��Nw{�V���ј�����D�\�+���Dm��>����U�z���9sp��Nwы�:묶�9���8�sF�a{���m�?E���c������DT��� <����DI�Z���>�󉍕s��G/بm�J:?�7���������'�D�t:��;s�Ν�K�����0r��P(��h46 xO;�wN+
2������Mg 2�7�ry����n�u�7���Fps�CƎc;�1�V����aC������łNm������qWœ~|�eY�6���׈��e��������m"��q�x�Y�����x�!([�n}��9��IDn2���J�r}*�:�W�M� <s�ܱr����fkl#gN�FW�>�2�Z����>v|ZRWͧ�	ܔ��^��. �x��r�#��?��g��>����W��*$��p�8�4Y�````��[�u��>n:OT�]+������Fg�nH1��������V�,X�7�L:�~wP/v�|>r�P�����{����D�(:
��|\M��1��w�a����=K�.}!�K$wS�i�}?��KA;]��꣍����rG=ϚF�j�D����[5?���b�|��X,~.G�͊��s�X\n:oppp3�L� j�������_����� J 4���ɶmtww��� :��fY�'�Ļ��ea���?~�#V/X�f�� ^(�Ͽز��T�����i��@U�4�B�}��ڤc�����<�;#���ܬ�fĲ,�r9��`A�H`I����8������{�v��|>��8�e�e�����/��A�K�RW�c��n6 �F�d�\U_��y�<۶9�3,��lv��]S����ϛ7���$.(�J�3���b�%�e=�H�g��~���_b:k```�_��A������t�(�<���J��Ͷ�#�%⭫��%=�D��c�=��v���GU�:�_0�j��w�'V$[�׿`:OU`:Q�8�>c�� � x�tj�T*�g�c��"����-����T��r�|��y�YD��Y\�X|�eY�!���G����M�`��C��cA��u�f���@�t
_*���y�%���)�� �͚�A�s+�z�� ���~ `��/+�J�&�	}}}�ǹBUo�ۦ\�����r���sPp\���Q�9�BR�}���C��ƍk��~����K�Ӽ��9t�,~���0��z���u+c?x�����<����b���j���ţ?��,k4�1��1wJ�;+�ʐ�q��}�l� O�H��.���:EZ:���r�]����|8���L p�y�����V�Z�3�j~ �P�H�K���KL��X��1wJ*����ƍ���{���f&�(�L���&:E^*��Jz�)�/����9�κ<���03z[شi��c��8�k��z'���Rկ�\���bpp�1U}�t����\.����i:��y���S,p���R��"�Z�u?�aÆI�r���!�3X�uQ__��b��u 7(��a�n4�2��UtJ�M�{,P@*���y��|<�-���r�Sl��Q��Tuu�\�e��Ʋ�� �B�uT�z���Z�U�y�N'"�����M���9tJ���D����~������t�:O�L,�+�ms%=� >Z�T�\�T~?�_x�}��R�B�uT��ݻӪ����C)˲�{�JQ�y�# ~c:QPD�=D����j�~ �6��&��fY���bǶm��������m7��,��jᩧ����1è�hM>��c�!(0�c: Q@ڶ���B�cǎ��{t���<tt�l�t�t
	:���J:Kz�}UD�GW�f��㏿�P��Ʈ]��h4�|�D�O���o:͞�p̝�ⶁ�������,�z��Lg����r,�	ǂN�ŕ������p]wx�/�nݺ�o�>�3���={�`߾}\5��n���"��{�ry=�ͦs���m688�k % _4�� Aww7R���(2t�5˲�����r�~�E��~5�m�Z_���l��V�صkj���A�D/����6�q�� D����jF��;��GT�B L��T"�l6��1����b�%=<���j�Zr]7��z衍 �	�T����޽{��~/I D�sK�.]l:͎�r̝bMDr]�b:G'�<���t�N#"��r\9� l4�c^���&�K=ϻ`�Ν��zU��پF�^Ǯ]�0<<��{z�c����L��٩T*�(��A4S��s�=*�� ֪��Mg��e�����Sb�C,0����u���~�f�y5�}3����={�j�LEGxg�X|��4s��-��t�Y��t ���y�@�t�$��S�bA�D�٬��$��~ю7{�GX7�_�l6�k�.��&���E��3��f����Mg ����J�~�!��\׽RD���,I��7;�)qX�gD\�y�9��>��7�,kZg�㩧�B��+=S1��~�t��e˖�`��D�%"7�*7��r�|w��|!��Β$c����w.��S"�(�i9��绮{���}V�������<U�޽{y|�9.
��A3�~�����j:�t���h{��'wz��j �?�	,�9sx�p�cA�D��rH�ӦcD�& �{�w���:�*��H{�ZmW$z&KD�,�J�S��1w��F:���t���6]׽�� ��W�m�����X�)���,Wҏ� k]���� �t�* ������!�ڵ��E�	۷o���4c7b����g``��fĄ����/0h:K�ض�\.�rN XЩC�r9d2�1��Jϛ�����vU����}{��������F3�7+W�\a8����{M� �*�x{�x��p��\০���9��:FWW�݁ay�뺗�j�V�,�:t&��H{�V3��nN�����43"�1w��V�u��4}O>���l6�*��t��K�Rk�g`A����f���e:�)OxY�\��� G3w��xrxx�v��s��{M�Px��4}����).6W*�ߘA3�q��Z�\~/F�K�Ԃ@T�R)�r9�1(�XЩ�d2�N,鏶Z��\׍�Y�[�lI�޽�����3��@D��r���s�����; �5��h
8� �祟��4,�4t�H�L�l�t�v��V��x�֭�ݴ�q��f�y�^?�t����f�L����n��e���(�˷�Z��l4�%
��t']����S���/z���;v0d<�b� ��r?*
��A����)�g2n2� [�n}�� �2�Ť�kO>sNaA���N��:b�����U����"b��ό>�Q�x�D��E��ƈ�y� �e:�xD��7r�Єq]��l6�j �2�ń�ޤY`A����瀞��r��旅�g���s���U�� x9�Nr�#�C�ԩj�ͦs�GU�5��±q�ƚ�y��Mgi'۶;q�#�!t"$������_���'��;�l�. o1������bŊ��s��q̝"�iY֍�CPxTU=��K�@�t�vh�Zh6��=M:ѨT*۶Mǘ�GE�J��� ����/�,k���b:���j���4u�t�f u�9��⧃���M����寫�k�!;�W�U���,�D��Z���3���e�ٗ��[1�e<��|���Xl:�ⵎ��t��M�6�p��DG����y��e� �'�EUQ�qk�:b�����J�u7n���"b
�p%���<�/����7���c�9�m����ڶ�� <d:K��G�iR,�D������_U#�i�z��L�P������,��j�ʳ�c²,!��G�l�2`:�ߖ-[���jg��t������ڄ�:^L�f6\���g���s���{�w��Bm�G�B�T�!hr����<f:�U��t2gǎzzz� "�Lg	Ş6�XЩ���C� �7��{�� �Y�r��ѝ�_m:��%"W�l�xPU�F���?4���ڰaC�u�w��Mg	SL��MXЩ��p�h����v]7���bqU�ټ�;�w�����A��,+����[�&�d����<����N	!�נ�&,�Աbx�r����R���t����ժz/�g��Bf���9��7��&f��] �M� �Ce[�ø�{���#��%NL�8�XЩ#��CQU� 8��GLg���˟����Ǩшy���L���T���(,���j��r�k"�v$�Fb��XЩ#�l��1 /q]w�� �)
/�m�� ���B�!"�(
/7��&&"s'��Λ7�.�!(���� ^`��,a��5)�:u��ݭ|����z��2�B�p����8�Y(zD�K�R)m:M������M6l���A���]"�
 O����MuR�XЩ���C�'�j��J�����'�ϟ""w������۷�t_�\�  �7)�,���j4�r��������t���l�BƂN%FcD�f����ܹ3��\���ȍ ��B����0.�T�v��c5D$�'�P�T*�_H�Jz��Q)d,��1btw��K�,9w�ƍ�]������Dd��,s�a\��52ED��m:E�I'��/�J�X�dɵ�w�B۶MG
Ț<)D)���!.z���J��n�u#{'aٲe�R�ԭ zMg���0�+����tz�z�~G:�V b:uU���4��������7�0�J�� �m�c���ݻ�j�̆P��@*�B*Ŋ�ɸ�N!cC"�J��.U�l9��뛟N�o�\�Y(~�a\tm۶mFN� j�T*u��=���'�J�/���l��9-�cl��Wf�p�J�J�W4�Q�d�����^���� �q'�z ���B�5�a�gM���	��A塁��-�CP4�z����;D�By�T~�eY�V�cp�7%cS��l�t2�+�hqm�+<ϋt9#w��4��b��E�OL�����	����k֬���ln�+ L���+�IZI����$9_�DG�1!U���y�(�P(>���2���0��A����7�MD���3P�����j�ڻ������ڵk���>������^%q%�Z�bΜ9�� ��߄)��~�QD>�yއ�^�ǹ���A�1�a��M砧s]�) L砎��r�̯�0<<�!U�O�q��f͚W�J�u��|���'i+骊j�j:��N����������CL�X,��ӦsP"�+7��$��S[��զ3P�V�Z�cY�_����ݻ�V ���?i%��lFz�����N�����}�<��X,���� ?'("���(BD���BU`:�笳�ʖJ�sm�~XU�����0����5Z�Jzįi)��ĉ�h��|��DyC8 ���}���@��,�h�0.bl۾@r���T*�A�����/�J_ؿ���u�juő?�V�a������.��J�mۓ���{�Iƭ%�Qm����z9_�t��T*�#9�tJ����� �a:���8� /4�����	r��'/�,�<�?"r�؏�߿ܕ�F��ݻwc����h˲�p��Dl76ꞔ� �W�)Q"<t��y�j��C�J�t:�^'"+Lg�� "�søh����@������T*��f͚+lۮ��v��7��IL��&�z�P˳eYX�`,+��'�׸������h�M�l��Q/� �}���R�9��pø�}����z����43'�tR�T*}���#��U�b �G��L�L���ݻw��h��v�m�X�pa�K:G�;�$("<�~k6�}�ƍ#�p��|��M��s؆q�5����N���G}�Tz�իWg���^-"�I�Ro�$���hL�l��/X� �Lf�q�ʶ�C礇��{�8���}+�hTD�~��jo�I9-x���W+V�Xf:����N�9(�Z���c�T*=�T*]��f]�#ǣM����?��RU�޽;�ŖT*�@DB{�v��5/��_(�":ھ��v��q�t�����>�w��S��y�f�� �g:H�SU-
?�7��B��m�֭�Ј�3�8c^�V{���������������݋y��!����5&�N��`��Џz�ب{X��y\A�X��h�&۶_��S��Lfٲe�|߿�|�Y�D佽����s��)4WG�$�N���߿f͚+���VU��L�90���l�*��ۇ���Y��D2�zzzB{�vu�d�
:�Z�|�Z���-[�<i:�dD�.
��k:�(���/�ȋ���q,���G�ڵk���>�?�f��;44�V�H�}����}̙3'��;RWWzzz�w��P^���*�̙��}z&t�����Q��n6d*������t�#��8��y��}�˲Z�/����c:D�k͚5/�}�b o�	����R���?w��@_wL6����3zf>
ƦH�٬�(0��S,Ep�}���s<�{�t��(����L� :U��ҥK�Y6�)�T*C��[�9(9D�Ufy��m�ڵ���h�}߿#�v��B�����������V��!��U ��S,El��aY֛]���� S�8Ή �b:�
�t�� ��� �LD�<�9(�{{����u����QU/�W e��jahh(��02:��~hύϝ;����{�8�<\A�؉��BU��f:�T���� �]L��˗/��f=b: %Ʈ�[��i:D�X�v�J��e=== �F7|���vc���V�سgOh�?o�<?����B��R�%��S�D�CHU���o��1"b�n
��t�)�ٶ�� �i:H���#4�D��CU�̝�$*�J=�z��\��v�o��@�Zm�{�j5�޽;��= �N�RW���m n�^�]�R�R)V�$��"�J�Fۿ�y�gL���|>�� ^g:�4��P(|��<�(n@�^(��U�lo��X������{ �[D�۝�����u�޽�s�lJz�u���U�VݸnݺC{#�Z���z�. /"o;q�=9X�)6"6�~��y4b����D�/L� �&�ω�i<v���m۶�P(l�%��P������t�$9�S�[������ Xe��Z���h��}��z�)s�1��i=����|���_��;��6mڴ�P(�#"� �"o�pW��`A�X��h��Z�vA\�����s,��B|��(D/����Xg:H'�(�զsP|��u6l���w�w��e˖�|߿ز�� ���x�|<�f{����&+��D仪�����O�?��b��U�@8;Ӆ������=�������s\�5�]i-Z4/��^��}�!:��\���w�ƍ#s����
,�4;o��5k�<GU/p�Ŧ�B�e�ԼF�qh��(%�AU���l~��G����ry��8 �1�Ku��X}�Qg��h��U�5�7o�n:�T��
���|�Y�fie�V�0�1�Ө�&^��,�����t��9���s�z����G�)U����h6����m�ކ�]���l��k��{��8��'m���:EZ�F��z��y�5d�������t� ��_
�ox���t�Nb��&��MǠ��'_�����߲��U� �zs������B��®]�vڶ}����A�����8γ |$��G���S�Eh���<����S�8�kT��L� 
�1�e}�t���t �/U���Qw�'���q�TzXD֫�� ��5�V����!�1�AU5������s�~m�����~ݰE�����"+B�헻�{��SU(
 �	����Q���dP����A ���fb[�R��tr��7    IDAT�(k�ڵg�J�u�Lf��\�����cզ)oY�O�91�UU�;���-BS�4M���H�Ї�=ϋ��d"�� Ǚ�B���|�t�N��- e�9(��7��C�N=��B�T�D�&��op.���\SU�բrm6�� ~����䋺�;,"o���a��bM:ERD�r��j��s�B�3"r��DaQշ
��L��0s���x;�����R�tn�m�f��2 +ǚ6U5z��4������E���VU}#�h�7E���i`A�ȉ�ݾm��qǎ��n�8�� ���D! �d:D'QUt��͞��j8h��r��K��e===Fv?ۍ}:��j�ͦc�[�.��=�B �i��J�)bA�H�ȇHUU�R�Tb3Ɣ�� �@���M����8�kL���e��Ӵ��w���J�R��o�X��k �@9�����zBIw]��� _3lY��)bA�H�������_1"��m�ϝS��\D�=�Tu�t�U�������߿f͚+ TF7|{��LA�ڱj�4V�_䋺��W�z]���(\c���p<������l�\��ss�|�2UM�� ���8ι �g:H�j: Ň�>�yޯL�[�TZ��Q���ȳ�Z|��f$�U�� �8��j�u��U�_�x񻺺�~`u���)�l6k:
M��	m�#N;�@�Px�����D&��?�J���I��>:M��\e:CX�;�<{�x4��np�D�����+遭��ر�@*�z����a��bM��"!c7��f�U�ͧV>�wD�ϝS'�۾}���t˖-� ���V����6"h/zы�]*�.ۼys���?��cզ#�>00�EU� 6׏��I���q��7���[�|�ɝ&CLG�TJ[��] ǚ�Bd�����n�!�l����h����3N�N䬳�ʎ��j���ȆoKL�j�o7� �
�S�zA���PՏ�za���*M������|�R�<d4�4�ر�r ���A�m�����I�(�D䛦3�V�T�����+H��h35<<lz�$L="rs�%�� b����1� :ez�FD>W.��n,���7��GM� �
U�d__�|�9�ϡ�d������1'�|������ �/���s���8x��a��7��uP�6���4>t2&w��t]��M���+W�Pկ���M�������p,�4�k6mڴ�t��k�ڵg���_e������N2�+
����cզ�GDw߶m�A���`��(L��ѱ���?Tu�m��Ӧp"�j6����Y��FD�tѢE�L�H*U�;M(.��'�tR�T*}����w���&"��3�+*Z��ժ��4_Dnqgm/V�T������t��(X���c5- �ڲeK�.8��{ ���AQ�f�Y>�˲b�yI��]׽�t�����u�J�sK����Tj#ǣ�4�+����׉c����8ΉA�X�\�VU?�k�Gݣ���.w�����^H��8/U�X����ŋ�5"�Tu��iߎ�DZ��J��e===.�u �`�Y�Z�z�tS�}������*��' �4��
��Vz&tj�|��y�?�0]���� �
�� ��q�l�b�!�HU�2��"�*�Ɯz��׬Ysa�m"��ٻ�8��2���TU/� 4�{�Ӊq��BwD�Q�q���2,.q��5㨃3��':��+QY5q7�%aIW'D[ۤSu�v6�$�RU�����L:��UunU}ޯW�B���!�^���<�ۣ�:Wԩ������!P!��b�;���M�B�ZH$�F�wD`�������4���U�f:���Xko �r������/z��ȓ�3Pd�2��mq����sٲe�
�U�il{4_QU��p׮]�P�ٮE@�Z�n���S�жm�v�GXZy��,Щj?��[k�AM�y�� ��ATCڌ1��:D��:���ru��N;����늮��_�HZU/0�U�����|~AOO�9{�����!�X,vgGGG�T/�= >9�H��Y�4&�: 5�|ӿ?�\���f%55�(">���q]C�"�$����ȭռ���e˖��Z{9� $�y�6�vc̪������RU�<�w�"iI�P��������N.��O���pv��UL>�G<G<��%��SU8�6� ����������&�d,(
�QO� 7�D��^&�y�7:�S�,[�����~k� ���y)zTuEKK���t�7�=�8O�R�S��\����t�[x�-����ʒ��8��=>��s<�=`���OV�P�~1��|@D����5�� ��CP�|����_ݲw���T��X,v��J%�WG��5��/�����H-Y��YU��f��g���?kkk{�Ν;�O�"A���_�' "�u|p�kKǈ\a�N�xj�pq��;�}�� �5�Լ���S�A�ȓ`�N�-���[�wvvv��% .0O$��LTXU�[DV�����������|�������+����,Yr^__ߤ��A�3��>'"�+g�J�Tw���N�x���5���y.�ՙ��z9���N�,U�����)��2�s���SDN)�u@�����W7o޼�ԓ�ɤo��p�b�9gxx�;"�\U'=-���m�]�^�e�W��Ø>}:����X�S�
gS�EdC5�5� 1�����Y���k���)anv�N�QT0��4Ջ�����<CD.��b������5|+�1����D]�y޷E�M�:�����t����"k�& ��֎S��a�N��v�@��X,v�T�p�������]� �'Ƙ���u�:Q�f`}"�l6;0��_��'���E����XĆT%{�� ��N�'�p,�J��ʖ�����y_�wNvI&������|���ʎS���6U�˩�"�����Nn>I��흪�1�9������G�0\�u���: �ůM���K�6577�ND.���o ߃�jPD��������S��ҥK�T��rk`�'��= >:�A�-����7�1WEp�{��#��˩�zC�vr�Ijkk��H$�nCT		c̻�t�։�^�(2%�v���z1���������Ū;=���P(|k˖-���|�����r]�Q�ȿ{���\.���^#�H�s�P8@���ʎSݫ�:����}���OV"���%�sձ�:::����w�é��^NE& _:���3�<s��������k��� p��~������X#�/�u�����y�\n�d����:�L��s"����W����Nm�"��ݻw�sq��J�R��'�9���1�|�� ��Ԫ��*G�iHU�?ҋ����Ƙ�U�- fpJlI���NDV͜9��֭��Dc�gUuF��߀��ܒJ���f�wL�a�M�Rר��Wn��^=,Щl\Nm�l6{���OF[[��x<~�U���,Ч�#��۹\�9���8�y###� "����5R�� �>����C���<�{��,��}P��~/�L�*�M��@ss������ 8���ʊSݫ�:�������\�|2DD<����]g!j��R��l6�v�VYk��bc����i�-[�k�� .�P)�0�ۦ�=�dtuu%D�ոW��i��I{{�+3�̶�����7����km@��_Nu��: ��S�"ri��-�}�] �u����Xk��:C-c����`[[ۮ���wvvn���	`9��= �ljjJ���7nܸ�Z�9 �ܹ� N���T����N8�ɜ��d~�?ʜ�"\���(���ѐJ��R���}�D"1�*�BCCCeJ41"��l6��Nn>I,xI,K��:Q�RU��St�4�d�c̤�pR�9sf�i�^��7����Ed��|e�ƍ��
��� �@�������s���F&z�����pV�c��T뇑�����+�SA�+�Ţ�#�4%����̟?�Ӯn>]]]�X,vX���j�y������e���iӖ����XU]+"�655-���^�8 U�2X�W�YCCC7�$���U�� ����|>��T�����\��1���鼋�O��ݻ���u�F����Ϫ�u���$���|M�ȥ2�6�ϔ�"��X,v��?��:�A��_$"���hD��d�7 >>�ss��oR���U�3�VV��^9A�Is��LU?2�^�fx�w��~�u����}�a������7 Ak+`c�U}��E�����ʈ�� ����JD>�yފɜ�� <T�Hew��;�G�iRS>�ᵮn>�dr�1�& 1�Y�� ��!j������y
Nsn(���0��9�x�M���7mڴ�u�q|�|�!��|��\.w�D�S�b2�|�1f3"�<�]�+�?qiRNm5ƼCU�.n>YƘOx��D���mmm|�:Ac���Շj�� ��U �J��'��髣\��R�� ��uBBD֌5ꛐ0� ��
d*;vu/?�4a.����'kpj�� ��Qt4555]�:D���--ijZZZ�5�įU]���tww�H���]:��K�6��W��.Q1OU�dɒY=1��}FD6T"T9q�{�q>M��o�_͚5�jW7��ŋ����_�D�������Vs/�:1`��TӧOw��� V��׺��{]�������<�y����M"��iP��6�L^66�}j{"W���G�iBNc)�������W���~@�u"�/�}�L�!j��r�A4777қ��p!�T:����s��� X�:���}l�'�a�����J*7Nu/�T2�]�?�F'7��T*u>��]� �#��u�Z#"Ϻ�@�� k��D� �����N���������D|������y�'z����G+���8ս|X�SI\~ө����ѫ��|�N8�㬵׹�ADG��������QKD�#����	MMM�cT�0�5Ƙszzz^���}U:�κ5U��_
�l�9h\""�X�`�K&rRoo行�@䇧]���T��V�e�w���������r�l�W" ���]��%���f̘�:B%� ����)�N�/ܸq��z�A�y�1��i�9�$3c�ؚd29�)*�l�~ _�P���T��k��E4y���}+�����擕�d�pR{{{���R op��XD����ˮCԐ!�������H$\�(��Ed5��vwwov�R�1�U��\砒��s-&�̪��郣���8�2����ۖ���,��Ӹ�'y&�}����!���A��ٳg/�־^D� ���mD�HUO�<�e�s���׹:=� 6��
 �����\������~7����Mh�ϭ[��@����Ot��i*"�r���;�ܼ�z{{G�0�-��^h�9�
�nGD�qO��I\}������Ƙ%�t�̞��U�t���^�,Y��{��(��DףAp+��T(RYq���@�#r��+�*W7��L&�T�� �2�,p���r���Q��E]]]5[�T��rP��}�G��3g.L��+7nܸ�u�j�(���A�6=�}���։�T,�`�2���Ot:,��TEc�;U��*@�d2�_A�������8�T�����"f��ݻ��u�Z����3Pe�X�������~:�>/�N�Y�n]Cͧ�<�e"�a�9h�N��>�U����9�}rX��a9����L&�Pӿ��t>�Apn,���[׹���r�{	D�#�u�F����-Ƙs���K����[�l��:�"7�\�3ꀪ�������9s��� OT(RYq��ı@�?��i�����wr�ؾ}�� ��`�1��*��T&�w^2�<�u��������U]1<<����璍7�u�5��>�����Aec �0���;4����
f*Nu�8�����D�}���O;1c]�W455%���3թ&c�D?
��קvn�	�Z '��鮞��U����\����O�o�sP�u477��DN�f�w��+��8�}bX��s8�ھ!��}���#n�֭�A��f�gc^
�j �s����\�:@`�^g����ҹݪ�Z H���+����\����@d�;Д����WM�X,�����/9սt,��?ݲ �T~�U&�y4���x��� ��7����}�$�!�LD�$��D`�< p��vQOO�9�tzM:�惠��}%�N�9�b�o�����"��lS��T0Sٸ��[K�P4�����e�ٴ� 5����� n�<�"�v op��dD5�" �|\�^_Z[[�;y+8��ƘU���w����-X��%�X��]砊[�H$���RO��OU/���
U.�|��Ϝ��t�|��3�X�*W7��\�7A�lii�U�BY��M�?�7נ����2�%���7n\����D$��n��:Uŕ�����|����ixx�Z�1"��0���v��U���;��#}}}# � X�L&_d�y�w `wj��$=�;����p�~���"�U�V�"�]U�.�No����y���u��8����+T��J6��{�w���S�lS��(��cDG	��bx�io����ھ�2@�
����Qu���D����z}�J�=� 6��
 ���W�8��d2y* Nmo<�y������ŮP��9qf|��hH�Rg��}�s8�7A��u�FqȨ�e �q��(��jii9alF
���� ���45ӧO�T�> � _K��[+q�F����R(� ^�:9��B���;v�)���W��
f���� ��:D9q�\���yuU��[<�8Q��+�!�*AD0mڴr^�xp{��3g����,�ˣP(|,�ټX,v�DN����L��P��@'W
�ڒ;TRyA0���n
��k� V��:Q�p��a���ո�ӧØ���{��|>����h�֭��鵵 �L���]� �D����g�z�Ν;w�HMl�FG���Pկ�a����a�9�MMMI +T�1י�\S��/^�x���ֻ5�3���C �c����yI:��z˖-����ttt�1�|���BΉ��"RrGGU�_ �
f�
c�N.�K$��:=�֭[� X��Rk�9"� �lR�j��u����r��͜9s����ꊖ���=Z�
�/H��A��r���Z��A���*��*�:��?�V-�TՆa�6��^("/p5�']�"�6�4�?Ţ�F��q��Lh�Dd�����t����g�����V*�J���ͮsP�|��+�	[�� HW0Ut�����ßu�J��f�A�2�{�z)�G\g"���;::�\���A�]%��ۃ߆��ۺ��WlڴiK��ј���E���9(��ZZZJ�nol��*��*�:U��~|Ϟ=|_c����s���A�b���rîsUX�P(��u��a�^�������4�!9 W��������V)���JXk�	��/�H����%��� n�`��TMO�a��!hj2�LO+��B +�F$T�8���X�נ#�y>`���~ѢE����͛7o�n2:h׮]��+\�Hk�	����g�a�NU#"+U�[�ԉm۶�
����?���F ��DT�MdĢ�@�1���H$�~�Qx����{zzn[�z5�:�J�^���sPM�����sJ=8�_�N�P�]�� "������A�N�� VX����i�����Ջ7��8��ͻk���VmPD���������s�-Z��xU��R�Jd�������%�����Uu9��Q�H�:U����=4�����b��@���]g"*��]�V�5���u�1fE>�Ovww�`q-"bFGGo�f�4/�}���(�lv��~�����X�S5ܕ��ֹAճ}��� V�����@�:�� �Ju�,�k���\��ӳj˖-�]�?���GD����D��'�.]:n��C�����l#Q�@���O��@n���=�5��bU��î3M���ֲ@����ܹ��yD������W��A5k����?�z����w �B�P�@�J�i6���ur+�N�s�ܚ N7Ɯ%"k �)�U}���\� �5@D6�a�-�9��:::ex�C    IDATZko��)4]�xq������O�}�P��@�JRc��]��h�d2��� ^�Zp�Ն���\�pMD�]Om���RT]�����8�u�yǎ��|�ԃ������V2�t����d2=�CP4A�� �(
\`��DD��7��A�8U�.g�E��|EUOu��ꃈ���<��㇇���
F�2`�N�bU�k��v�ر'�O���v �x�u&�#�����ѷ�a�mÉDb��tx��_�����Au�UDJ���{��}"rM%�Ա@��P�չ\n��T;����� �Z.�;�Z�z ݮ3=�1�v�:�u�D�z���g������A���W���T�ޚJ��zpss��Z�Hc�N�`c���A�IUm��Ap�XC���3b�� ��@�(U����|����|��� }UF��J=�����|���@����g2�G]��7�P�c�Y n�r��{��{0��1���{�uz�d2y,��8�u�_�zQ2�|q��'�k<U�H4,Щ�D�O�2��� γ�v� v'&W���uW�zd=�M�C�s���j���\g��3Ɣ<��u��A�I�"�:�����N��� �cNp��:�����Y�G���OU��0BD� ��鮳P�x���'�zpSS���Q�Hb�Nee����T�2�̣A\b�y�Q�j��F��lٲ͜9�b�9�O� �˭s�������uj(FD>Z��c��_�`�$�TNw�a��uj�L��A\""/�5��Uǜ������~�g�vuu-���SU��b��D�1
�۪E����/�sP�Q���l�\`_����@�r��� Ԙ��lo6��PDNf�Nՠ�u=ͽ���sٲe׍����ZD^@T��1�A��:�Q*�z �&$WDD�*�� ~/"_�`�����T*u����:�<�+\� �T*�LU?�a�yQ�=={���{{{G])��O>yn"�X."�p����!<��GĞ���%c�T)���ϱ����ujh*"��f�K9��<OD��ե[OA0�u�r�:���@tP6����lk�9 6��Cui����k]��*1��v�k���V755���p�✢EU?��<:�������9�'���R��r9�v%�İ@�r���r?w����0\���:U�B []��R���O?�t����Ý��[��w�@g����p�]d�2ï�Ax��rc�O Lw��h̹���Y���O�w#�:M�����]E��j.�[s��ǿ�
U��:������/Y�����kyWW�m�Ba;��]x�㭵(
������0��|�����PՂ�x��B ?0�u���D��a������a�t\�5�}`�������ے%Kf}\D� �:�6U=7��E�Mͩ��z�1� � p, ��?|Xka�}���� �n��]�  �L��1�H��Bt8"��l���bl���
G���[�w�j޵,Ω����=���_�� ��q$�aƘ� "W�wuu�.��h��'k����<��"
�
�ְg����:mmm���`qN6���~)A<�J�6��++���:M�>c�*�!�&clk��M&��c>`��LT{T��%K�4��������~����������b���p$���g�Y�!]2�<6�H��E���پ�*�{J9�X,^m��q�3�Qp:M��|-��<�:�T�ax��ٳ_�J {]硚3ghh�j�4�L���K=�����[Tu�1fC>������b����������C4:��1Ƭ�R�Y�JT�NK�x��Y�,�i��"�E�!�ʡ��w4�k���I8�쇨dc��+�;�R��o�}���8�g��"�tr�
�35]GG��9�!Ֆ�|�U)�5}�Re��ѰI\D�Z�8U�N.�{��D��y�%"�9 u�t�*f�����rOs
��kT�l9�J��T�ǹ\�|�9���� ���B4Q�zg.���R�M&�ӌ1j�=P�5��:M�1泮3UJ.��9�H���Y�&�>{�Y�p�	�����_
�] �?6B�⼱���\�hd�/���j����y�+J96�gU��
G�q�@��x(��v�ATI۶m��%���]��{�dN���X����T��b���� �K 5��:U��~z��%9�x��٣��,Ω�ȇJ=�Z{-�b��8X��dp�95�0o���K��5At$�HI;��R������-�B���U����*��`Y`P(���M�C���\g!*��S���R� `7wGX��D�iii���D�����t+T�� v��C�t��yg�Ŏ��������f \���ţr���OU߷s���U�)�Cq��8��!���	MŒиX�ӄ��W�E�U.���P(,UU>U��y�4w�T*����P(��� �Gʩ4w�r9>w���}�������BTfoJ�R�K90�{<R�<t,�i"
80͗�a�رcO.�;_U/��-:�ߋ�̟?F*��g��zU�^ o0�u8�) W�ш����Zk9rN�*���,"�V0t*��� ���\� ��\.w���@��,I��olnnΨ���:�&�B�r���,Z��xk�`C8�c��V���%� ��p$z�4_r�(J�0|<�˝�`�S����v���R�]�D��s4�����|>��\g!��fU}_)A0n9[u,ЩT���~�!��FUA\%"��u���jއ�n�:�:D#I&��B�p?����BT"��N8��c��_w��*�TU��:�_��Vd������N��ND4Y�ax������c�1� /p�����b�)��0p_���!X�S)���w\� ���[��r�q��Ө�<DTS,�+�0�z���
��z ��U������cN���It�@��R�����?�:Q-PU��y%�m��Q��R]�h��l��@IͲ����B��Β�=�{ vW8�a�NG��_w����d��tKK�)"��u"�6U�k��O�9E*�Z�. �]g!r�_��䴣���;
����!�:���AT������f�XNy'�#��Ƙ���-w���y��jU�����E�|c�;J9�s,š
c�N���q=��A��s����Qd�HDV��w2�<�u�z�J�^/"?0�u��`WWW�he2�mc���X��xF��<�>$*�L&��ǻ ��:Eګ�1ݾ�߼p��\����_�����:Q���w���R�+����ơ�?ܱc��9��E�ӹ\�� V(��CD�e \\,�|�����\�e���M ⮳E��~XD�h���� `��
c�NG��pD�7���j�[ O��CD�6��<�K{�w��0��������h</K&��9�A���� VW!OC�+:�����ݮCիl6�k�) v���"��"����/.^�x��0�@D$�J}��\g!�"�R�S�+��@��R�o�*;5UP�AKK�_cnv���"/�ݣ���y�W�z�F��Օ�<�fU�W�Y�j��|�?�h�r�<^�<�:��~�u�F���7��d.�>}z���_DD'�ȚT*���c\���d29m׮]��"�Y�j����K9PU9�PA,��p6�a�'cDU4cƌ��͛�X������Tu���&���\g�������X� �:Q-Rշ$�I�hǉ��`�ۊa�N�íՈ�lѢE?�����y�����:Ն6c̏|߿n���3\�q)�J-��ޫ��t����%�1�r��� ��B�����/_(��:Q�Y�zu�7�1�3g�O��:�pyss����3]�q����DU}�Q���Q�(����T�0��:=����{��Q,o �"�3f`����t"*�"k�=��_%"�����Ӭ��8�\"*ɬ|>�OG;�X,���*�i8��J���D�l޼����oii�ܹs�.��J���ݱhѢ�]��4���������U�r�ҥ㮷��Y �U)RCa�N����A��T��C��H$0o�<$	W����������<���E� ���BT��O?���v������hX�ӡ�A0�:Q#+
k <s��1�7oZ[[�"��Yk����A���2��}dl�+�\U��|�h?;�Ν� OU)R�`�N`�Y�:Q�۲e�~ ��^�5kfΜ�u�DT�8�O{���z��."�T*�U�oh�GD�s����w@oo�(�T)O�`�N�.�ͮs�� c�Gzmڴi�;w.��o"*����ttt,t�c���ڦ{��CU]�:Q�P�-�Ns/3��# ��|_U�s�q�� <v���Kg�8"���
�B����:�D-Z���D"q�s]g!j0�koo?q��0\`�Jyt Xk׸�@D$"7��z,üy����\�DDT���T*�V�AJ�J�����t��BԀ�Z{�x���*�i,�	 ��ax��D�G�X�& ��1�`��٘6�M���dͪz������~�睮�X�:Q�8�L�����~�ZaA�0Supz;Q�<��C� ��hǉfΜ�Y�fU!Ցz�������A���7��� �s������b�q{?�a��\���=����D%"Gl�|����7o���D�_(~�dɒH=��}�
�2˽%�"@Uߵt�Ҧq^W ?�b���wr�'��\� �?5cƌ� �Q��lGD���������""���� >�G%������w����Za��58���EӺu�
"�͉���p�1Ǡ�������3�H<���\X�dIs2��6���@DG&"�n�6����*ũk,���r:
Q�YkK��~��`Μ9hm��P"*�" ���R�o�������;E�վ7�FUOM�Rg��zAU\�L��zc���׹ADG����<8��D�f��̙3+���� �$��S�uÅv � ��o��(Tu�QtNs/������îC��&3�~дi�0{�l�H9#Q��g��;�JU|��T*��P(<�ŕ�����Tj�^�6m� �V1O]b���8��6���|��ɞ��҂�s��;�j���Y�"��sUu��_�{Q� �9ҋ}}}#"�*�K|�ָ
(a�e"r���wl94i��ND4GU�hoo�,��=�{������6U���m���3�9����N�@o\�s�;-Ո�Ls?�މh��Zk�������6jW��W �i!Qm����rɑ^����@ M����D�eӦM�x|��9��}ڴieHED�X k���։���M�<� ��<���k�{��m2��S &�ܖ��z���]g ��Q�[�q�̙3�ᝈJu�1��d2���ɩTjA"����ED.��K���k�9��h��zcz4�>�!�hb���M �����DD%��1?�}�DN�}�dU}@Ż�Q��ȿ���O���@o@���D5�G	����lii��y��ᝈJ�R ?I&�%���}���`R#�Di�-\���p/A�+ �*�|Gրb�XY��Q���������x�ܗ&��s�1�["2n�7��� p;�YՉEDUf���?�űfq4	,�ϐ�v��D49CCC��S���b1̝;�މ�x���ý "q�������L�zwY[[ۑ�K�:�I���sOC�C��������7+qmc�Ν����J\�����T���~�㎛�yޏ ��Q&"����D�͇{att�. �U�SX�7No'�qƘ�Os?ԬY�0}�������<�o`�---�Ǳ����8�'w�ܹ��U�RX�7k-׃ո���^U��=f̘��Dt4FDn�}��b��0�]"��{���'�Y[�0��zQ��a>�:M���P�{���`�ܹ��ND��f ǹBDUe�."�A���`-�I໮b���v��q+�g+}���&̙3�E:�G\ �����X,.��l6�>ҁanA��;��j ����N���A ?�ƽ�Q�Vկ���Ap����cG;A����	��aU�>�!��|T�����m؈���~ �xA.�{W����,"wU$Uc�� D�\.���DT>�6mZ`k��g���9s���|�cT�Zq����r��6�� �+� 's�x<~g�s�=��Z{��DT^z�����̞=---���&¥�DDD5�w >a�i�������S��؈{Y�5�c�� DT~�x�z �j�s�H��1��C�DDD�/ p���=��2��Se�6��O ��Plnn��u"*��z(�����{l "oWՂ����mp�X�k�0,�1\�>1l��6mݺu�u"��AU���}����|����� ,������h�Q�υa�-U��L�x<~O>���-�
G���ձ�������j;+��,Ή��j��l�־>�Sr��͕.�`۶m� �U�>��zc��u "�����QU�N����Q,/��}���hB,�����f���jP��վg�b�^�
����� �_���T�<� �m;Q4��R,�Ap^�
b�a?��@����ٳ�u"�����_�\���۷�{�E�~ �ZkAp����a�F�&����z�{�u "���q���Q<�lٛ����p���ApE���@A�`����z��]g ��hjj���J�g�^N�!""��~��|a���rO�t\�,��\�X�:Q�x��~/"?��=���ϩ�DDD����^���*��y�q�{	�z}���"�<k�"��J\�X,b�����4�HD6�ū]tc�
k���p|�h�/T�D��H�̦M����ĵ���U�ĥ���h|��"r���Ҧj```�}�sD�:f���v����M����0FFF�}Y"""�>����y�l��u��R�"��9��z�D�X,^�O���Z��pDDDյ�' ��^��qlt �X�ׯ�ٳg?�:U��͛���\�{��gam��}""":�� ��0��� ���@太5;�Z�$�~m���u���P�D�5S����{�Uރ >���~4�\�.%�n�3>��ׯ�� D�Nss��<=���۷��ለ�*��{�zFgA��z.�������r�#�X��)Ue�����T�Q(0<<\�DDDD4f/�U�zb�s�܃�U��p��8X�שX,������S9���DDDe��'�1�A���r�q�������l6�}�u"r���{cWW� /�蹣���V����<zT��0oUU.�f'�q�@�O[��OD  "7��g'z޾}�*����QX ?��^��Z�a�DU�E�u��������D 0��`BCᣣ����JDDDT��Xe�=1��X���\.�$��u��b�^�D�: ~��'U������s""�	{���0��t|[\�*Nq�C��ND�k�����s""�҉Ȧ�i�\_>��ED�u�#�X�ן�\.���D�-���m� �ю}��g���������Z��0p�Fq�8ŽΈ�c|zGD�Z�zu�7�v\>�g�v""�#pm<A�Y�O��<�:CT�@�?��Q��� ��������������l��Z� �+�����T�r��V lzs,�댪��u"��͛7����Gz�P(p������"��Z{N�A�*C�+U����aqz��:�����ýƵ�DDD������_
Ð[�U��lQ��]��u�Z����P(�I$� �u�筵v����(z �J$7����bu�Q�a�@�/��I���`�!�j0퐿�9�;m����EUg�H�h�U�� ����Q)���! �aj��"2������!��{���"����) ��bO
��bO��Zk�1�P(<�ǋ�l�U-�����b�lٲ���k5������0T�]�NDDT�FD������r�]�i@\�{,��K���.�2 =ы�w驼��Da "G��D����U�Cރ�����<�� {�s�<��"2���Ed�����"�WUEd������bO��}"����S| @�b��-��s    IDAT�Z��}hh�U"""v XU(��cǎ=��4���������5������-M��f��9��/,��y��?���BD`�}΃  <ੱ����O���?�I�m��S(v�a����_R�ڸq�]]]�x	 ����P�ΌDDT�Dd����0�m��۹s�n���p��,Q����:M���)�Rf�}�?������}?`��� {Tu�1f @�X,�Xl{;ǺiR�U�j��ለ����o��3��TG��<���t�#JX��c�c%��Ƒ �`��e��b��(��i����=�E$ �]DU� �M,{b���;\�P��b��
��'�����Q�q����NU�� |-����u:<U} �C�@�#�|�7%���/!",p֡}��������xBD�(��ijjz��Nk�C=���������9Ցa��X,�
�p��0T�'\���cdǎ����)�4Q� t�}@Ua�A�P(����(�U�u,{4��>Zb�BrDDn:�u""�2x����� �t�Jg�}��:F��@��-u�����9�$� ,�8�`�;���}�� ~%"���=a��Y�c׮]!��Q���Uwq`�6cw�!jX�׏R��CD8ŝ*m�?����{���}�@�cLOSSSw__߈ۨ�-�M��lp��ܚ�d�r���&��m�<o@��,Q��~�vǲ@' N���Z����g}�� �a A0��e��{��f�9���J�4������0��:���}��-����,��GI#�"b<��*��i ^1��/ �����t��km�1fC�ZF���%�6�9����aE�AU��Z��0�/h��m��}���W�A,��9E�lU}-�׎5���?�#�Zk7�a��JS���ه����HU��ȍ�b�Ɓ����<Ty���:C��@��X��tct�5�ұ�wc���n T�~c�� 6�]iD$�y�ߺ�ADDt�A ?���̆o�GU�9p�G,����L&�����xS��:�j�| o�7�*<�۟J�Q����---�mݺu�u�(�}���z��DD��Fܡ�kT�{��޸Tu+�?b�^����qtt4���MW�Wx�1���E��� �^U���{v�ر�u�(�֞�_�DD�P�[
�­��L ���9i�X�ׇ������%m�NT�b�/"���q���� �12�̯�FtCD�s������lR�5ƘՙLf��<-�bq�1Fp,�낈dK=�P(p�բ������}?�~��X,�k��s�Tj)�%�sQCx�U�5��z%Qc
��Y��v���D�:`�-�@��b	N!! x ެ�o6���]Ƙ�Tum����: յG�� J�a�8�� �`�^&2�^,9�Nt"r��.�|l�}��\���z���Z�W\NDDe�,�u"�b���0K~OJ�<� ��u�(`�^�1%ƘD%�Ց�X�9k�U���\.�8߄$��iƘ�\� "����NU];::��ݻw�s�j��d9�� �u�P(�\�[k9�N49X�."�����ݹ\�I������T�&�9�����p���-�?m��-T}�:�:CT�@�}������t��Y�r��M�R�Xk׉��###�EmDAU_�:Մ�- �Zk�N�6�����ס�D���j�ԃE���G��Ψ�"r*��777}�conN8�{��t�qF�DDt8E٢�w�+��߿s����CQ�a�>�z��	����&�$���b :tc>�k׮}�Tꡱ�k3�LO5�w�q3[ZZN��=��(���oP��"rW6����P��X��a�^�&�^��mֈ�o����k��!>�ݶ}�����LFss���"�ƴ_DQ���ڵƘA�Et�\.���"r44�5NUwN�xkm�#�D���C|�X�����p��ܝ���ʽ�OD�*����(ҶxPD*��RU��C�GU������u�X��8�5��11��E���KDV?����"r������p��2\�����Y٬�=������m۶M�!Q��`����Mt�"��i ^��� ��w�Ƚ���E�� &�NPD��S*�������1UMc��b�����E�Z����zJ��,Љj�|U]."�X��7c��S�T��v^u�Q� ���Z��X,>���T�Tu�KqY�׼X,6��R��'�]�����= n���<���O(���eGDy��=c���Y����v�!
X��8k턦�����:Qݘ�\ �c���� �BU>gΜ�{{{GE��qF""z��� ��w�3E���D�ڦ�g��3�s8ŝ�~��$����೩T� )ס��X?�GDd�����i�D�'"{�̚z��}oo��DN0�~�5�ic{�Q������y�\e�6��{NU�I:YH�S�T�,]	����:���QFq����������8#��Ό8�˼��Ό��D �����6�t�S�NHwg��|tC�R�9�T�s�+�$9��\Iw��<�y�033�xO�3�De)�OY�Y�[��� �A'"""�ƈ�<>{��&۶ojj����7i:Q#~��F���T������4�y^<�J=>00��t(��bAz����!"""z��<�q ��%�_���fc%Gkk���Ą�Ʊ�7�Jf�-��NDDD	5�w8�YqΊՇ���I�u��k:�I,荭��M∈�(���>+���>n���\�ת�GDG�XЩQ�j%K�9}NDDDqR�S ���� ��ܹ�OU��QyDd��v��az�,�r�QU>�NDDDqbOLL|`xxx�� DTUM��c���V�wp����b���%�3nDq!"c�3�Ƃ��XЉ��(�Dd��DT=Π��7� F+��;�Q��j��DT=Π��74�_�=�(�����Mg ��q��э�{C,�DDD+�e�`:UODX�M�ʉȁ
�aA'""�X�:Q<�*���@��,������:Qp��74�h��7r'"��ض P�g��t�x�`,�]������s���"#"hnnFKKR�,���o���"���0==���	v2BD8�N��Ƃ޸�[�n�*�&)���eYhooG[[�q��m���hmm�ܹs1>>����#�$%z�B�U�D̶�ɤ�`Ao\eϞ\�NDD���ֆ9s�<o��"���6���bll���ڱW�X1��� DT9U�4��4nנT����%�DDt$"���̝;��r~���͛W�XD�R�V���:,�,荬�� t"":���磥�%�1[[[YҩfXЉ:zê�t`f�{�Y����͛7MMM����҂9s�D26ѡT���&Q]���t ���T�`gЉ��P���hm�vⱭ�-� ��t��N�Y�M��T�K):j�ܹ5y.u���*��58Π��7���6���A����m�&�e�6g�)R"�쳙�b����U�M�3�DDtP؛�O�K�)��t "�NKK˴����7(UeA'"���H�g����k�z�,�b�3�D��X�T�E�X,��R�T�^��3�D��X�W��W��;�K��=��ץ�t�gYV����7�*��Wt~:Q=�&qD,���g�Uu<�,DD�xT�LR;E�����qU4����A'""�ڒ�[�PT������:###\�n: UL*��X,r���P(j>�m�5)9����d:Q�X���T����0gЉ� 01Q�}Ck�z�,"�u��qB"jh,�JU�� �95�j��-:EŲ,������W��BD��i,����Y\�NDD(��ͷ������s������DT����j:N,��7(U��//�� `�޽�?^,���H_��M�٭y޵jժf�Y��r���M�3�Ƃ޸8�NDDUSU���Fv욪bϞ=Ǝu�d��g�������fqD*�J���@���Y�A'"�gMMMadd$�}��si;E퐂 \�NԠ,�J�
���t""
����y�LOO�2^�P��O?�xD�b��ټ�-g�q�|SY��r�B�3�P��:��P(`Ϟ=ؿų骊}���g���9��a3�-�T���Q�,�bA7�*������:�����SOa߾}%����i�۷���U|�JV��b9��:,���Y�U��t"":� ��~�߿�m���	�mCD`Y� @(�����l9u�w�깧�~z磏>�7��*P,����[���7(i��vΠQ�jy^:Q%����J�R�_�!�
�7�3�*�&��Y&ΠQlLOO�
��N�`D$�K�Y���8NK%7�:�������122����e�̵kמj:�NU��`z���e�:v""""�T�����ݻ122����+�-[��t6"*�eYsMg0�Ϡ70Um�T��T�:������MNN�����N�up�eY�6�FDG��,�P���tE3�e���"""J@�� >�n?��A�?������6���f��ܤ�.qo`�3��7v"""����eݾk׮�L&�C�q.9餓:L#J:Πs��USйĝ���U�"�hjj���dR�� �q>��L�#JU������� ��&t"""��I��+ �²��������eݔ���פ��%���� T9YX�}MMM{
�B�q������� ^�g��ǹɲ�l۾����t8���g:�i,荭���Ϡ������G��x&��_U7��m:Q�$~���5��ܴcǎ1 A�Y������UU��E۶�p]w��Wuvv^����b:Q�K�:z��
�� �9Q��a˲n,
�d2��]��lgg�M#j@�M0�K�[�K�`�����(Lg�ϳ,닮�n�!�����n���4���-2�4��VMA�Z
"""":�������8��dP՛���OL�#�'����1��4��V�w P��<j�����f�ή۶��u��EUo�?��[�n�2�Ȥ����OX�]�3�"�t""""sVX-"�=8������\n3�]�J��v���UU��u�����.<;��ٝ�d�V�Aܒ��=��j�,�nA6�M���N�{��r�����>-QՋ \dY����UUo�ۧ����o: Q�,�Z�	D�Fg�޽{1��ro�:QC /�� �t:�.���3��o�,�~���g$
g�����D�DTP�+�������J��cY�g<��������ܨA�������e��g۶W(CDDDD����>11��u����=,����� 8�����7<����رc��8 ZB�DDDDD�8���eattt�u��03�~*��o```��D�#"�Mg�,�nv�{�TU]��� �HDDDDT?���;� (���[ �������|>�3�� :M�,�NU�Vq{,�DDDDIbx1��ȇE����� �pGGǣ\Op,�qP�w P��� """J���x/ ���\�}���mo��rO(� �����8N5������*]�>{/�3��R8d�=8�3��� 6�bY֣�\������8�2̬�H<���t ^hA����VD~��"�Ϧ�Q�Y�ͳ?0[���yLD� xTDU��y.{r�Hj�ҥm�^�`���>*!"'�,��KU�
��]�i��^�EdCwX�uG.�<���~ �j�و�(��9 ��قUp�OD~�OD��''''��m2,������������eu X��s��߇��"�q:f������[�K:��op,药�u�e �{�aR��ox:Ql��Uu�eYr���c,;�,�DD��������Ү�H��p]w@�'1S޽ vȧ��;v���ꈈd2���Ba��T*�^(ضݮ��"2?��"�`��,P� ��W��� ,˪4J___�d�s��Y,�1P,W������?�� BEDQ+ ؂�sm7�x�w���N�rc�Z���h�=�| kf@Uqp��B� �q
����W�!˲����U�,���V�۶�l��_,�r��^U��'Ie2���B�N�R� �,��PU)��g�Y0���� f��������"ݮ�� ����q�� �-����������a������� X�ͫg��ǀm� Tx�o �<�8D� �# �W��&''><<�������o]�}�KCMHDDT�f������#�<��S����u] ���� E c���_D�}&ZU�"r���X�*�)��#"����^3�6̜E?�q�g��������C�v+���HwTAz�jW��,�D��p���*"wz��LX��u�ʂNDDqs� /<�o^j�,�u^�kJU�*� X�g���@��7�!�j����%>G^���[�,�#"""
z�X�c@D*.��k>�Ad�v Tu����-�w��W���r�\׽�kk�zDDD���o/�b�u[,�0OCaA��j
�t��zFD6 �5��|��M�o�*:��	U-�zq�X\a�6�,�x�����y�uݝ N1�^���`���͛7�G���� ��BDDD�P��msy�!X��aβe˖��fU�("o;Q�����j��{L:��[�Ne2���'Mg!""��({wn��{,�1���|2��
�eYU���:O XoY�M�\��7wU�X�ʲ,t"""
��>^��At���cA�	U]�
o8�,D	q �� �����<���q]���q�DDD۶-�z���\,���m�~�P((x���l�̳�7�������7i:PH�,�DDDT��;v�,�D��A��Ǆ��\����#����x���p���,����?i:P�.]z�]��@�t"""j\�Z���8N��qĂՖ�{B�(��;� �)�N����?b:P�z{{�3�̿��?��BDDD�KD��s}&�YAkTyz|�@D,U*��. 3QyTUopS>���Gk||�������0�����VY=�F�Q���G���� �Jn�m��b�r$��U�Uu���$�K��1<<��u�o �s�Y����1�H�K�_� ��z���
��;v���[ ����n����t:}����w�To� ��eY�H��BDDDgrɒ%�-�Ue�8z�ض}2���/"w�	��3"rG7MMM�x����L�g�|�s]�Z �5�������<���;]�m\�~�	�`u���%"	+�!� ~�G��߫�|v��e�C�Lg!""��Q��X�Â#"RUA/
�H��<��'"?*���2����e``�	�u���Lg!""��R�q��.�$�,�=^^R��CCC�]������E)৖e]����W�0�+ �!�=����JW��/�,.�;�D�e��8N5����
C�m ��5��uy�w����},���<�w �m:5�,�rn�m��Q�id����e�~C��_��(y ?�LymA�e�@��,DDDT�v�)��#�z�T���� <R�J�pMo�}g�k/��� |�t"""j�ʽAUO�"H�cA��j7�Sբ��V�2���uA����c��y������Z0,�D��0������^Y]D��eih\�?U�Y� �(�q��gZD~�5"rS.�7�~/����{%�/��BDDD�˲��
��+Uu^Tyz̨�EĮ��g۶o)
<n����������o߾�t:�T���
�A����>
�Gʹ^U���Qp�{��d2�V3@��������xTu��|YUO�<�T��d9������DDDT����Se���Ϗ�=���bO�c��ad�ěp���[�l����>��~Ygd�y����/L� ""��T�q��G�%�1$"= ��fU�AD��)UDU��"r��y>�A�    IDAT< T�S"��6�����ꇪ����3�14[Ы2;˹=�8�S����>�ϟ���WX�����GE�Ǯ�s��A\ww�| +#���X�cHU���WG�ȍa���py�Ppr�ܺ|>����S�i�9����~LOOo.�� ր�Q���S[&�9���2��'ÉD13-"?	��|>y2�ȫ 4��ADDDu#�s���rnPյQ������(���������<��pRQ��?A�s>�ϙC�����R(��	�Y������}򓪮�"H\p�{L����E��0�PcS� .O�R��.c9O��˗��P(<�s""":����bA?Π�T}�O �?����<��������E�a��ǹĶ��n:՟rwpw���Q���R��E$���j�inn�����(����Q�S 7A��|��a��N:餎�����w��BD�OU!�����(�N��A�eYYn]tl\�_��^� }}}�"rC�����9��XΓ�uݵSSS�YΉ(,,�D�;�o߾��{Ί*O\��ǘ���8׆1�/� �\.��\.��t�=�u/px6)߃���Ϗ�=�T��a��t������ci���,�˽��M�!3V�\��q�[ |@�t"""j�s��X �e���Pf�{{{��4���n<dY�+g�yY_\)^2�����ӏx��,DDD�PʚA���|	���q���[�q'��,��2�xȩ��}�����}�Ð9�V�jv]���z�e��QC�J�ӏ�s���2�0q�̢�r�;�c,2�̜c~���W+��L4�uWMLL��g��DDDT�G���'ʹAU_U�8����,+���U�("?c,��) _K�R'y�we�_H)~\�};���a:5��7�����k'�ٱ��ƣ�]�J�>��߿�t2oժU�_�	�Y����ᕵ�pww�
 nA�3��wFggg[����0ƢH�VD��y�E,�<���A��Ql��e9�
�s��7,������ ~�X� �wtt�4���j:��u߁�O�O7���b�N���fv�ر������t,��pnXA����O �����S<ϻr�֭S��y���-��~3��7����KUo�}�|���,D=U-��sU��%bAO 	��> ` ��jU���]244�]�	 �8�ɅB�Kډ(r��k۶�PU������|�t&"��C�\��B /�(K찠'��ŋ�c ��e����I��_��~ٟbR|���Ny�i��Q��N�Ro�̼GX�dɇ �b8E����炽�d��J�Tkkkh������� �)
�x����}��n��� p=��y�(�&T�m�?����;��D�~S��(RAkkko97���
G,�	���-s�}#�ma�G%{\D^�y�%;w�6��Ggg�) ~	����Q"������G��9����B O�8E�񾾾�rn�2��'Gh]U�w���k�ZZZzr�ܽ��P}q]���e��Kډ�v>����|�:�7��(�FY矻��	�䈲�zr��jժya�J��������R�ԋ=ϻ���o�t����~�9��Q2��U���c)���y�y ��)QL�jY�E"�����zr����C;ޠ�������KUw��:��.���&zVgg���Fp�v"�!U��󼏕s��y}"� �"�ED5�J��)�z>^>����kB� ��u������Lg����d.�,�A �Mg!�D�������Z,��\.�QU/��`D��?|c����mR��'������Z�<M����r�u�|�)�a���H�u�/��O�]ډ���J�RV���wx��>Ս_�sqWWש :��_,��rʊ+�����oLUok�S _���xa.���t�?'�x�b�qn�Y b:%�����OT;��y?������(ky{��*H���'�쎪����/�����<ϻtxxx��0T2��+S�� �&GD��+ o
��S.�� �xDT;A�U���ݤ`AOU}C������0�L���MOO����]��P}r]�êz�Mg!���2==}��yτ=��y�W�{\"������'K��u�V ��.N|��'�y�V�jk0U-����/!��=ϻlhhh��0T�,Y2'��\�* i�y�(q�,�ܡ��ȎG����_Q�OD��_�j9G,��-�<qƂ�<����g�9�eY��x16�ʎ��5�\n��0T�:;;Oinn~PUי�BD�toKK���D�"����_*"<���1����"I� ,�	$"�.s��r[l	s�z�X,��y��[�n�2��S&�y�eY8�t"J�_LNN�A__�X-^LU����{/�[j�zDT9U���5�Lo
{@��Gv ���jpp�צ�P}�jDTnN�Roڽ{��Z��֭[�� x�{k��DT�g|��ԋ�/_�" 'E�'�XГ����+�0�J}3�����4��TU��JG��d������FDTs"��K��=���*���455] "�M�>�=��zq*�zs�a�=�
��[�o��� ��� �O����y�3��W&�y�����+Lg!�DR _�<�����&�l۶mtzz�� ~c2=_���U5�պI�P"rac�Lt�۶W{���2w��q]�2U� �FDf |��+����Ν;�U�����t"�=۶K.�V������zB��N:�P�u�m� ���� &0��kw���o:կU�V�s�z _�P#"3�x��y_7�p���"�z C�� `,��=Z�����o �a��cAO�����P���>���0�l������9��/���x �;Lg!����U�����鳏����~�OTO�+��-��T�=�� }�;�oD0f�*`�\s��y���o�<B���y@D����GL9��~� ���B�pw�z�U��E��W�=�D�M�W�u	��y���u�	y9�5��}��� n0�t"J��wtt����M)U>�@U/0i:QR�jɛ@����`^�q�=�:�����U��
{�:� ���\.��"�
˖-kw� �~�%"3&|��K�e����w�G���T>��ԋE��Q�I
�aL�(��7773G���쮲��<��|>�����N7�N��]��Qb� ^�y�7M�F.�����	���a&�P�Z���"b� �<���No�P�l۶mTD�s�:p����K=���� T�\�}�eY� zLg!�ĺ�P(��y�C������k |�t�$��^��+ ,�0Nb��Sg&�9;�qc��]Uw�ȅ��]2<<��t���|��7)"2�������;w�6&L��}MU?m:QRAPrAWU��tB��3����7a�[K"r�Ss�܍��P�����OD��6�'�T�t"�� x����c?}��2�+L� J�����e\��Ȓ$:���^�>�[�Yc ޗ��������0T�\�]�8�m >f:K҉��DF��u�T��|>��,Q�<���w�sř��^굙Lf���$
:����2�A���� L�=n�~iY���}�tj��� ��BD��WU/��r����GL����?���b:Q\�s���D$�X�	 ���/s߾}�. 7�=nD
 ����+��C�!�ɼADp��,D�<"�����f7PK�|>�� ��t�ڟJ�~Qʅ"bE�#���  "r�����A�D��eY/�<>�G�s�S�z3����Q�����w���o:�)����\D��t��������gW�vF�'QX��ŝ���
{�|>�|��DE�?� ��d:5�l6�v]�"�/�fpDT{7��j��������)�o��B#%���wG$�X��Y�e��<EU����a��ay[.��h>�?`:5�%K��ٵk� >h:%���R��{�wA�;+���L�G|�t�P���E$����ǂN�R�wf��t�~@=-�MDN��iT�L&�����^ o2����("�)"/�}�j�aꕪ}߿DU�5������r��R.t�< K"Γ8,�t�v��z������>����O����R����/U��n:%�� ���r�<��aꝪ�-[�>U��D�+gy;wo� :=���/�q��b�2lp��y_�3{T�L&s>�{���Qb���}���y��Hz{{�[[[���t�FdY�M�\���ݢ�F�'�X��ptuu-{�|>�3 a�[𵖖���y�x}j`��~pv��y��Q"L�����}߿�(W���o���i:Q��r���R.,
o�q�DbA��5ApQ؃�j "�{��T��<ϻl��5QIDD\��fv��A"�é�թT���.�k:O��<o<� �m:Q�P�����G�%�X��y�Z�n��7LG1�ܖJ�z|���T����Ϙ�BDɡ������0�#N��������x�t�q})�\�r)�7D�%�X��yD��L椰�����>�q3�ٍ�f_��d�V�jv�Z ���,T_��4D�t�1˲�u'}}}c�T�"RҲ]����|If
����'���NG"���H�r��ߨ�˸Ubɒ%s&''o�N�Y����ϟ������t��7g2��C�Q��mۯ��t�z%"ח��YU/�:O����ѼO"�.�<�v }a���������F06��ʕ+�677ߣ���B�����e!�J����-bQ�(��zČfJz*�:3G��a��bI��3�� /�8N����ќ��9a:����8��?�<���!�K	��ݽbzz�^ g��B�����9??X�/^���vX��Rh>Ň�4���Ĳ�7�5�����,�BU}�a���*�X>Š�B�1�x�H�R�y���Ƣ���zq�Px �*�Y�>577#�:�F��eaΜ9X�h�̙۶k��b�$�q^e:D��ijj:�8��P�S��x�^��	�� O����Q��EQ���s��a ?�b�K���;�R��/_�� 6 8�t�_���ǽƲ,���cѢE�?>���j��b���El۶m�MMMo PҌ!Q\S�E###8!�,�ǂN���E4��Ux_^U_�y�e����:��b�q��l۾,�t�m������E���X�`N8�.�J�+���fK���N���_�r��| �0ĂN���(�<�!����T*���]Qd�dp�t� `��,T����mcΜ9X�x1:::8�N�hU�w��۶m���>�ݦ��""�.������#�C`A��{��n���/���/��>�6�jtvv�9[ι<��ɲ����������Yu>�N�PU.s������---op��,DLA��R.�m�R �V,�t\��,zss�� �2ϲ�s=ϻ���+���uݵ�e�`��,T�����fڶm���'�p-Z�����n@G�����ɓ%j���o,�7�����z���>�E"�R�?�A:��=�/���}}}� ��h�/"�U�������~mJ�q^�6 �Mg��������T���.\���vά�sX��'�3$I>�?�N��
�f�Y�jED�Y�u���o�<�84��J1���%�#���(�� _�<�m�|�Gt,�Ϝ���tjMMM5-��ts��98�>����d*�z 7�L��uvvV�����b�ҥop��,D5��y��r�eY�F�~��J��( p�!��S�WqI;��uݗ�>s���da={^�g \'"�3g�����7�������ԴXUש� p����,��C$Moo����.u�,�F��_VU=�u��@U_W�L4��Q�z�y�����`�� ?�,�O�D��0��p+��9���,�����D�� n�����m۶��n����V��sD� ���Z%�.�]�!�FU�"򁮮��b��.�y�"��P(�t�9fNt
wS:&)���L&�JU��t�����y���."�8�Ş��M����3cY�= �Lg����ގ9s�D1���U�aӦM�U;��8���ZD^	`������bFD^��嶚ΑD"b�Z�����q�_Bqs��y��իW7���z �� S��x���t�0q������?�����5,�
�q˲��9�ID�^�^� ���b�Ǐ<�H_�����c�k�w �ͦ���N�,�U=CU��� ���'Վ�~�'L�H"U���Z������7�(,� J:�xtt�"�w9�%t*GS�P�0��5��H�-[�$�J�`��,�xB�� �;Uu}�P��-[v��$������?����8'��� V�� ���h�,[��/����(��̙3�-��޽{M�!����$���J���o�T��d��8��D&uww�O��?�"�Y�1��U�a�S�z�������ٖ-[�H�n��7��9��lz׮]+ �$"˂ X."KUu��,�̬�rp޴�t:� %�D�z�G���즶��˲0::j:Q��T�E���g[��6�0�|,�T�w��� ךBtPggg�eY78�tjL�m����Ƿ��ɲ�����뮻
E����G,����n	��3�!��j��.�<�V>tcD仪�������(��5���r��R.�m�2�=7�����:ՉիW7Y��c g��B�����'D� �oڴiSԙ�E��	 Ϟ����y�eY,�sz&�Y���6��D�� ��nnnƂ022� �i��X,���R�s]� �y4��\�l"r��8���A$"����w ��tjlG9Z� �~ �,
Noo�7n�"I��h,��o5����ΐT���;U���?O��X�`�5�;�+�B��t�y�(8�N�,� ��tJ�����CU/2��[kk�o���KD�S�z{{�����Dx,n�]��������=ǿ�"�] ��I*���g��E���J��W�u���p�q���UDU/���tM��r��|�tj|���{T�U}��������6n�x5��щg�k�5����T�t�� ��5۶�p�B�Ӝh������w�x�{,�2:U*mY��2���uݏ��tj|"���c�-ڴi�%�6mZ�u��)ә�����#|��1 7��ea��G{L��^��R.������q��S5>r�I'u�A���{|�t�U�'�6�e�f�i +M�H"y��8�2�#��w�_ttt�����y�J����[J��q�7 xI�y�8XЩ�&''��tJ�L&s!���$
������p���ܹs%�y�I�,ΐ����x�h�?g�̛7\�@�DU�����w�a�$,�T���l
Q�\�=KU�nnI�z����L�h4�m�b:C½s�ʕKM�H��G`~|�kZ[[�����N��N���(��L&������S��ݻw��t�7�u_ `=���&*��\e:C#RUt�����?`:D�w�Mss3.\�c��8U�\�r��N�+UMU��t��+V����Xl:��ݹ\n���ݼ���m:Dmڴ�n ��K�RX�h���j����T�F��Yʵ]]]+�=�HT"t
C��8\C�[�x��b�x���0���ED��t�F�����8���C$�� ~Pʵ�ea����<�LP �/���s~�W'X�)�e���/�W�njii�	�3Lg���=o޼��ѨD��>p�8CD���%E����j���?Zʅ˖-[���D�JǂN�P��:;;�6���ADdll� ^g:���<�2]]]��M��[�/_�e:Dmܸ� ��sOkk+�K�Z�F��MMM��]*�JPh,���(��?ͥ����6��Q�EΞ�۶mujNI���N��p�B�R<��"�u���J�p���sU�#Q��S������c:5�L&�Q n:�ֽ����6����ח�^����`Y��0�oYl�ƢE����CI({����)�����Xa� :�JU?k:5.�uߡ���t�/U����̲,��r����;M�H��~x;��*��ܹ</�B����}��]�\�l��X�    IDATٲv�dԙ�|,�*U}g&�Ym:5���W�_�(:��z����;��U���	V�fqG����%����~�ԋ�����=E��Sج٣�J��ݽ�X,��g�P��������X����3���!�(� (T3F*�����R*J*U��R��-[����"�DbA�(\��*�!�1�Z�j^�P�QD���B������D�p��tD3 �6o�<,"�GD�����ب����kJ�8�N���PX�)
6��M�����f�����x��,{��|��!Y&�Y��|uHU߽r�J~�iFU��u�(6۶��BD>��A)��Ξ�Yđ�
,���wvvr)$��ݻ�&"�7��⏛�U/~M�_ͅBღC$���ԏ�k��G�577�5$���r��m�^����p�����STl˲>g:�/�q��goR��omm�������7U��l6�6�#i�lٲ_Dn
sL˲0�|̛7�����LA��R/���nQՒ�'3X�)Jwuu�j:��q.����$���\���7f:G��kuo�����L�H�Ж����w��N��|>��R/.��<�<t���L�����dֈȷ��?T#A|�t�8�z��f�����(�>��{[[[�SS�]MMM_��K�,�Ó�� S����_�+Vt��M �N�je ���m:DL�l: �+�9�t�����V��_D0w�\tttp�;�o۶m�ԋ���?>{�X�)j���7��s]wa�X���@���Rw��������"�eY<�� U�d���ZZZp�	' ��V�_�s�Zgg�	 >a
:��y��dƺu��5kּ&�Jm�%�TK*"%����K��+p���{\��4�#iy�{��u,��w
D�����`��_�a&
:Մ��_��v�>��֞��֬Ys����GGG�*
]�sQ�ܝ�嶙"r��T�4OȨ=���Z��ܹs�`�X��'��r��R/���tU��Q�p�_5��k3��L���d��֬YsI6�����԰�ܨ�޷oߒ��q��(�D��Åg�� T:������j���PMMM�����uɨ�T*�7��`Y���D��"��N5��_������:�;��^���s;����m h���	�߿�hFJ�����?2".T���,L�R�5"i6o޼��Z���`�' ��}�|m2�o����J��u�U �a� V�Zzigg�� pV���]��TU�HU���w������hɛ��JU8<<��t�aAo0"�i�7I�-U����]�_v�ҥKG�z꩗��� 8�ƯO���ҥK���D���j��=˲`�6���MG�+�ͤ��������&dݺuv6�='��~5���Al�ݙ��h��E����0%�sqy{�X��Ɏ��t��Q��(y�]�cǎ~��_� �2P�D�ӽ��%7Y�u�RՋ��TAKK�<t��N˲>n:�i������sAOO��۷o�� >�;A�={� 8iC������q1�h�
�9�|"�#�jl�����K/�g�u�"U-x�w���VUw�A��q.����T��Pǧo455��m�1�:�p��8�L���:��3�n�>�N?#"7��� t�3���(�E~pO��w�9~��m����f�9�|�z��8��Α@5�,nVS�Px����r�{&''_
��03�O��m��˹�q�u"rNT��e�6���LǨ[,�d�|˲>g:k׮]��f/�f��Y��kv��� ���޽{155nH�2ٶ���Ĳ,.ool���4�ǭ���Z��П��<�Ry�|��Ph��cǎ�w�_�zu��}����M叅��P�?u]��s$��X====k֬�"���:�m ���rԁp���PrUa�����Cĉ���70�8��,7�#I6o�<�v/�����e�Ῐ��nU��T�Z��:A|�����>�n�c777ò~_A����X�ɔ��t/.�=�ܖ�kמ��f�����H��&o/�5����oOw!�f7h�A���ؚU���5V�3�gY�B��G�����}�ݪ���5�E����|ɳ��,Rտ�2S5R�������Q�u���t�8:��f�ًzzz�޻w�� n��&o'��Z�B###���A "?4"n8����o:D�
���̹��7}߿.�N���7�*U�g�\�rn�+ ����fngR
��z<��+"�-Cp�gv���|8�ͮ������M��F������Q�s�<��s��cAo|�
�¥�C$ɖ-[�Xo��X�v�Ǻ`���|߿PU�`o�rQy�R���sCgg�) ���yKK�s�����O)AT�7e8����C4��kמ��f?;��[��\��M��Q���bdd�B!�"*	��G�$��z������{g���#�#.s?���W�ŗ �+�HT&�������cY�?���*�J��N�e��Ă� "R��@D��y�Zi֭[gg��s������Al�E���[��c;ՙ���沖��-^�x.�L����B��^�9�DDn𔁗�XJ\29888����03�?�XT�_-Y��k�ܐ�d���M��cNr��'�� u��d���������n���`͚5Wm߾=�^ ���T���q����zy��Q��m�6j:G�477s�<^>#"u� �z{{�\g�W�q�/+�bUU��^,� �a.:�@U/���S�իW7��F�����|Ķ�5�_��7i���/1�^�u�Y�֬YsI6������n�QU?`��lSSS3��9L-%�;n;';��6�!���&˲�S�=�����}�l ��9T�*��Y�=###��"U�����A>��cR �l:�Ig�uVw6�������b�8���p�9��T,1:�IJ�;#,��t���z�\n:@�lڴ�~ ;����=��T�7�j��+d<~,:U�e�vYG�9���_D���[�NGǂ�`�������u�L�B�!ji�ڵ��Y��l6�[,�cfW��0�E]	� ###��t��P՟nݺ��=P�n�(tk\�}��I�3Ӄ?0�ҋ���Ϋ�f��~�J�^�J ��b��X������=e��O����C���r�z�ꪝQ��������e˖����C6y�j6��� ت���c:۱�*��Ƹc;�%1�g"�g��.g��*�k��1�D?����	��.�,�5 ~J":"U�=��}��{�����uQe�FSSl��S�����X�β�z[�I�ӟ3"L�l����炞����o��4f6y� �p���۷����c�HGG��!bl�� �7��{��I�y��' ��֯+"�8�Ӫ����K����L���˹AD� �5>���e���gٟ�=a��)U9�r�ȟuuu�j:D5�<��ų�������(���w�arTe���oU�e&7n�vUO&q%��L����
(
Y]����\o����sUXQ�uUv�"  w��P � Xu$�骆I�:������c�1��L�tu�S]��y��'�>��L��[�=�� ��֬b���{���!Ĥ���}&�irT�m�Q�#@�fq�,�
��-�uG]�=����D�)��
�?4�۶?��&Z�ɺs�A))�cf��TD�ۮ�j���F���őG������������2���I ���6�\.˦pBk���>��� �J�l6ۯ:D�\@�&.-�����y.\��p�N�A�c*��r3/�f�K |�MyZ�H$t��$)�c��S*�4�*҉�X�qޣ:�T��X�jժ�Mޞ�}�I 8�5�Z�bǎ�c1ioo�J��U�A�3Zu����ry �=.�i͚5���\�<���j"��{�3���ZC���;2u�%�L
�����D�Vwf�(���:Ǿ�?����GyB�%�V��(7���+Tg3ˎ�B{Dt����3K�����8�vm�LE�{������Ʈ��v��GAf�g����<�gͼ�q�S��M�Z"G�G
����k\�#4㋪Cv�a������jժ�w�޽����`|��Ū�����.���}ioo#)�c����s���%�������}_��t"Z`]���@ϔJ�O6�����pi��$�N�vts��W2f�ۈA������d�{Е+W��Z�����;��� 7Nl�67�,aA�XTC����o��~�:D'3C6��f>-�ͮP�#~��_?��a��̯9�#��s�|>���1>�.ǾL��>4<<���פ�����' ���D"�:FG�=f�O$�,+�41ø�����}3Gy�����Nl�6HD�a|���|�J%�����!D#����bf)���`��T��"R��N�e���lf�L�M_���/�����74�?Ц<36�]�_Lvq))�c�ы �J�ԪrH�\|#��kך�������_������7� ��[�*�
v��!�"��N�b@
��xG&�y��q�̷أ`ܶ������<�x g���/����j�Dd��>EMЬ^���2C�Vw":/��l�>��U�V��z���6m�T �+ �8��V�N�s"���1У:��IDZ��ir��^"�M�ЯZ�zuhK��w]�r�0p_X�ꎙ�-
n3�q�#̼�]�fʲ,imo)�E]�e��� pUӟk֬9p���g����X*����|���ǌ��;w�Z���!D�~944�]u�N�bŊ$��s���Z۶W�#&�W4�;�phhh��y�����;4�B�py3/�m�`f��
4SA������KI�3�^���x��-[>��_\�fMo�9�V��I�Zf� �`v{#FϞ={06&����`fioo��{n1�!n���Cu�8�={��l	{\f~)8����u��M�<@SǊu�������_KD}@Ws�H*�
��'�N�҆��S�pW��/Y�d�3Ǐ<��CW�^}~�Z�np1� @�6 ��E�ND�@u�Ng���ov�8�!:�}��W!��������85�7o�<�f~�gU�P�s�B�ͼ���xm���X"���]f�_J
1���r��:
 �L��&���6mz5�g�����Y�\Ʈ]�T��Y���;�:D�#�Ū35��? �Fu�NGD�1s�rOl�@���3>�zٲe?*��_p��,!zl�_i�K�.��]GK;&�H���t��vi<�C�ͦM����&o��M�};w�DE��)�㋈��f�oP��ӭ[��7 �v&��mӦM[\�=��O�ԦiS1�s�\ó\DD��_�e����[��^������ނ�"###k���<�9�J6�Q����!�}_
�c�/�X�'��D�b�����D�N����� .�����hhhh}3/p���|B��T"�h���R����a�i"�L��`�b޵k�\�3�k�.�J%�1����O=��C�CĄ�A��U�m�Mu�N����*��L�F�r]���_�	�y4 ��ؗ,Y����)ό���ey�RR��L��N��R	����cD���|�D������"Z�:�P�:�Bw���������+Vh�>](~�p���� ���03��u݆o���,˺��6暑v����d�K�Qi��qquu�s���ݻQ�TTǈ�ND�Tu��t���������:�����:Y�����re�u/$�~ ��3SDt��yM�βm�C:��'�I���:F�H�3A<�jg��LH�9=���}�vy�!"�Z����\�@ ��d2�������w�`�nm�/���7z�w4���V��IC����h�Gk��n��V��q!�������e�ٳGuU<@D���3Ϭgf9VQD�S�B���C�Y T�Cha?"jj�hΣ�>Z`�_)���zի(�a�̮�^ND� �Mu�1��m۶�*�e��U �iQ����q"�����.m6vػw�.紫6
�.f>۲�L.�;vxxx)3�RL�V�OTg�����!�b��8�_����T��[�D��
�mZ>��u�S�y-����L���|�Gͼ�q��Xݦ<3�ӾSq#_��	r#"�]���,3_`m�X\���N^�~��>��۶��>��h�����<$�Je��B+&��U��d�r�&��M�6��<�&��p��,u���tS��L�hf>�]�fJ����H
��	z�;�L��Lę�T*qjup�a'Ι3g�������r7mܸ��/��8k��r���}��3˚c�b��f���ѩ~���ng�f]r�G�T��3V(�q]�L ��Ӳ'p���@�#-Z�h�a���C0mQh��1�X����M;.�t:���-.��{�"�Lv�O�M��߹~���S��e˖-p3���B�����y��q���|I胙������������� ���L�|4ܜl:��������J�rƏeS}�s��?l��D�R }m�3ca�������hY�O��k�.�~���C� >bY����]�n����Dd�����CI)D�ݯ:@�����򱱱��ѩ�Ν{;��
�>C���,��{>�� �򔏂eY�l��l�� ��Myf�4M$����arOGR��@X��M����عsgT/�� �"��T�Ճr�ܱ�\�|���C۶�
��E"t�'�aH�.&�̟�8J���+�]�Я����&���x�w3���
"�opppG�ٶm���hg��P1��{���]&�NkӪR*��w�^�1����a�Sv��y@.�;yݺuW?��#��8��. jCF!T�=D�]L!e��7I�_���U��Dl���03{�wu"�{�+]׽�ѿLD]��L�ӡ��.%��c�St"BWW�6������d��:M��. 7�_�����rO�mۯ�M�D�<��T��)��T��m� \�:H�Y�|���6m�`a�C�-�k�"�M|�δm���[ n�pO�����8�=qfNU'�̠ONf�c���N�20�N��>��D�9f~e.�[������r���q��� ݭGB+똹�:D�h7�#������E�Ct�o��
�FCgW�\y��q����|�?����wx�����F_�8�qD��6di�ʽ�d}rR���%���[d�V�ص��/�Vd�{|��}'���Ol��l  �`Y��+�&��=|�T�ۿ\.���m��͝�"���b�Ba�뺟�
������im_�x�|��ԯՑj��%��L�iG�*Jt�vu/�k���":�\.�~��s��%6lx�]ڶ}�7����PL
���V@菈�&�ɜ�:G�ٰa�C �T0��+V�У2`�����c0�GO;��ņO4 "2M�
 K;P�DB�M�şI�.�B�Vw ؽ{7��r��>OD�3�)�bq�����\�n��{챑vXc��i ��ѱ�y��14Wu �a\�hѢ�st�RT1�~`*��+ㆂ�}�u�nY�!hm9��o۶mw�/p�D���""�R�����G&�mR�*��g�33v�څ8 �6�' �	����?�
ztl�>��� xD�z�󼆏���:����D�[ ަ:H���g�t����������0�3��f�5ul 3_�y�/����	����CWW��ה̠��ҩսR����
� 癦��\.wh.�;ob��Ћ��&�[!3]���Vu���wьS'����r��A��oY�bE,��u�hѢW8@���������1�9 � �i)��L&a������I�3a_�����f��p3�mYV&�����.|衇��ƈI��Wx��B���T�����4�����L&�U�èhs�N�RoU0��\���D������ �q]��M������Ř�3CZ�5'-�1���%�J�Z��Z��>�dv��˲�=8x���&�;���=7n�v��d�ُ1�Z�9���!�--�b���?Dt����N�����a\��w��[ ׆<�R�|�I o�d2'�� �$���>��{f2��A�|u�n����Q�{S�u.�v��wm�f ��q�9s�_���\.w���y&�9��D���    IDAT��:�a`f)�C�H$d������m��Ct���_~��Dt�QG�0�quP(�L&�+ \��5�̛7��u�m�Y��΁�I3Z���d=fT赝"��F���W�ZŎ;�͛��Gy$�D���.2�& 	�Y�wuu=�:D���߭:���3��O
��T��8>�1�r�|��y\-<��;���d�c�7�=7n,5���K�����pT�e��>�~xD{������r����3Ϝ�:G#�ȪT*7B�34�h��3��Q̌���|H�(�6M󺉽D����� ���
��J�Px��c�8�u݆��z{{��j�& �9^ӈH��vY39)�cF���N��ju�۶OWb:�m_�5�sioWC
t�*f^966&K���#�� pO��ѫ׬Y���fac������F�~�R�:�Um�4c�T
��_٧YM���S���Z�5BDteOO��;�g��w 8Gu!�DD�ޮ�a��F���?��fOQ��C��͝*��;�Y���U瘌i�H$��hW=q�+)�E���ns|߿���w?�A^,�ɼ��/S�C������Hf�E@����f��,�Es�̹�ΰ�%�w�=fTe2������ѵ�]LM
t�D*�ҭ���R�|�����r���s��V sUg"l�jU
tÐ]e>3_����(���� nU0�+V�\�*�FJ&���q+ -w_K��Z�����wL(AD���R���j��J-�R���`�9�P�Z���G�,��q�L�\�!���T����b�Y�T��2�f Tg��eYZm�<iq���B��ѧm�^�: x�w���d-�f����V�!�Hf�EЈ�s�L��9�,����Sa�KD�""�&A�m�WX�:�d��mϧIi�M���bF�'U�*IDt��8�� �|�G ��W�E��ʊ�t��a�uG������} 7):�z�j9Af�m���ix=)��]������I���W�pǲe�� �����^��>��8Y�3�}�h� W�n7!��͝����E��� |Au�z�����bj�8ft|R�c�;��r�|[oo�O���Sccc�#�;Ug"��\�0��3��uR&�9Ou��Z�n��P��O���ӿW:$�L�f� -7?��8c1R�-h���Q�j�j]��oݺu�뺧Bӣ<����I�.چ��#�ɜ�:GT��
�����{��q�c����a�`��,�tuui�-+��]E$�K�Vw0��m���5�\u]����/ �FZt�?�W�jU>WD;Dt���>3��_�h�ط������� }��ԓL&a�ZN�&I�3:��ט��k[�g�y����<�b 'Avx���A���0��������e�l�֯_�'"ʅ=.3����_�Y�v#"�T*W 8Zu�z��k���\��$z�����H$t|�G ��m�ժ���u���<���,Bh��yϪW��.Br�m۟W"�Tl�&��(W�L�� ���ٗ�.�H�3�?��}�h� !��%K�����B���4�� ֩�"D@6�g��.Btn6�}��Q��7@������f����Uu��Hk{�]h�0$�I�1^���q�ng�n޼�i˲^໪��*"ڬ:C�I��1��d��媃DI.�{��~�`��:�(-��K6�}-3Ku���z�,Z#�В�O�� �9~�fpp��y� ���#�L1�f�⌈��C�if����o�� ���ݬT*k����qj��va7���Ku�R�ǌ�-�������L���������� {U�b&�hHu�8�}_f�E�)�W�r�i��y3�QCǢͽ��w�a? ���,SI�R:Q, �՘���?"�vGJf>=��|]u��x�w����pUg�Y2���i�e�D,�5��|Ju��x��w1��
�>�#����� ̟?N�Z��e��LŲ,$	�1Z���0I�3Q����@D��l6�1�9&S(!�� �~��0c��q�����"����m��:G��hs�i��P1n����t�ff^�:�tt��jV�&�$��^*���f�/۶}������O�����Uu!U�V7��s*�f�  ���[�d�+T��]�v� �Cwd�;�֭[� �W��L'�NwLk{�&���]��4?ߑ��L&s�� ��<�4"� ���+g����E�D��1M���˗�SDwc�|�������~��Y�L�"f>Su��tJk{�蓓]D�eY�,Ku�z��a�d��᪃L���|>�i"z'd�8���� qW�T�@���T*]��F�:bf%m��Y�l6�q"�����|�jFt�UM>�b&�O����tn�ُ�~��dQ��|>�=f>Z6�{Ju��۲e����Ŷ�SBw�<��}P�`�k׮��,��f��d�U�hD:�6�uI;i[�1͟�7ㇶm۪���y�c̼�}��1	)�cf@Iu! ��8��U������=C/ٴi�k�(�q���W!�P"�й�TL�H!�e�&�ɤ�S�!��-[�l�� �
�g<��+ ��:��bf)�� m�B�{zzUDg��_�h�H��g2���@��:;,�C
t9�TJ�Vw �+��?����Ou�z�����@�=Z0�i� )Ѕ>����lW߆r �P0�i}}}��m�>�0� ��:K#���:��]LM�*G�z4ou�WU*�d2�n�A����a������"��]�]���r�|�lW3ߨ`���͛�&�$�ͮ �{h;���d2	�����	�a3��CZ��h�4o���׺}jhh�~ � ֫�"�MZܵ!��
3�l��gU��]5G�F��=��.g�8Pu�F�!��1%��*�
J������\.���i߻�Zd��T��O޲e����A=��,�:������bfiq� �q�BG��m�t�!t����N��'���Gb�A&�q��� ��҈N<Rm2�2q4�P{��ɖJ%���6ThדL&��ݍY�fMZ�w҅P��Qe:�r�BD�0�㪖�Dt�m�|� O��T*���y��BL���ʞ��Ǉ��T����u �y�43�
�;!�۔ŋ�7M�G zTgiT&���I�A�pň�"��n߾�������s (�Jرc���1666�x-��n������m�[��7���u���T r�.´{�֭{T�  �>]��}��E�-PD7�r�z ���%"���m�>в�{����4*"�8�I�A�]!"J��� �1Y�Z�3�<��{_ة؉B��2�϶��u/� ������ 6��"b��:�'3�Bs��e}?�;���c�=��}
��˕+W.Q0�z{{�#�8Lu�fġ�]LM
tE&��+�خ1�۷o�t&�Ӥ��t�׶�U�h��y{5��Vď��k��d]h����Lu�0�u
�5��no�����*�ʏ1�	ndD�(a�	P�ma��Z�މ3���J���g�ٯ�ш�[�����9/]��� "�A�c��8�s��:I$�@�)Z��/_�|^�R��ժ�4#N��5�^�̔�
L̞>��*��6R�ԋ!�H�����!3��m����(�u/'� ��":���}_f�ET|1�;Uu]<���� ܥ`�#׬Ys��q_b����J�ҏ��y-�ck{D�_C'�G u���E�Tju}�q�ϩ�Ѩ|>�K���=�:��<rĚ>d]D����e��H͔���6wT*�w�w_Q.λ��b��ީ�����O�
Di�_�� ���#�J�X\<7����O�!�n!�N�������#3蚐5�"b���6۶m�AtP,��\��ѻ�s_}}}sK����ܲ��t��pD㧁�4L��Z��:����R �C��� �l�/�R� �H(9\�e!�H�\�̒�Oضm
��s���8�q�u .C�?�BL�4M)�5!���Zb��-z�������smܸ�������<��V�\ٿaÆ\���f��pT�c�*�K"�(�ǟ���:DP�U4n�g�GI:�F�Z�̿��>�8�,"�gf�Dh�u��m{#��WuyR�k���D�Y�/��+��UD�6*�G��:�_���D�@�������{ �	sܠ�R��,��J�{G}��mO8"��; ��϶m�2"��u	��e�� ~�:��6��e�&�y��B���3����C��~��_ ����ޱv�Z3��-[�����#��y"��Eg�h^T
��� �$.3#�V��y�m��QT�[�y޳��	�y谇i"4�\�Uq4��3oW�A��"�sG�zh�&:nP0��?��O�c��K�..��?pX���"7��q�I��]n��V�T*�]1��8�w���#�t���u���T ;U���j变��"������:�JD�d7��6��Z�dIO�Z��C�=V�D��!��T.R�(NO��]]]�c4���nٲ冾��H=^���wT��W���,"R�� ��T*I�.�.	��l6�\uU֭[������N;���v��d^n��� "��M&��k����1� �@2�Tc&�V,���뛫:H3�z�!��^�BȖ�1Ϩ �l۶m�D�!�8���X�|�<�AR��>�\.�u;޸��畆a�@d�ԋ�=�QT
tY��8��$�I�fh����b��۶T��\q]�<"z+��*����@׏l':�+K��uD��V�q<(�}��A���8G���+ K�~�0%��Xއ��I�FE�@�� ��b��fG�U&�qTiV>�����É��Y��|ߗ]?��.:�_۶�M�!Tx��7x(�q���Gq�~A��mۯp/��zOU��"*���ڐ���J�.3����`�fd�t"z�a��m�`�Y�U(\�u_�s��mbr�I�~�@��}�l�c�C(�b���eYo��y�`N遼��Q)�'�qҰQ)�;�^Ղ��n�q�"�� =D��L&s�� ͚hy?���70��y�^��]K�4Etf���8m�a\7��� @E5���:��~ �M �9�2���Q�˲�G\'�C�(ֈNp���U ��7g�ge {������ g�y]�,Y��a���;�Ej˘###Q~P����S�½��̄m����/�Q�Eh���ޢ:��3�q�� n���L����,
�V$L�W������~�R�>�装���q�s\p&��i$�9U7p{��	�~|�뺑_���h���|��T�� �|�\�[����ۢ��X,��2S�ø�q�wG���<�#��m���� :�<�Md]K��.:Q�0�;l�>��?��� �]��Db-��5�""2m�����K/�{Ѹ��,k+�1V�>��Cn�o�D"�3(� ��8�'U�	f���{>3��i�y�ZR�뇙�@��@"�gѢET	K*���^C7Յ��חr�zĤ8�)��mw���I�� 3��rX�fϞ�p��J���U@ .�m�""��?�󼟕����Xu���ؘ�1C
t�ɖ%�;3�L�� a����wѝa�����W�~y#�q���⏙��v��Q\�t�A�\$o�;�� c�y��`͹\�È���"��ٶ}��8�l���y�_c|�w9�!~x˖-�!�~�@��H�4���3�b7w ��L��K��x �k�G_q,�e}rq�P�3�p
���g֬Y2{>�0:���m ~��dRd&j-� ��'�qD��3��7�)�E�c��m����a`�{��HKf~�T�8Κj�� �CB���b��R��:Fhd�prR�+�̛ ��X;��ܹ��������}�ݻ��>^m�o�y�� 3��C�bq%��Ug���v=IW���O:��A�!�-�˕���
�~�ʕ+�'��qN�3 ���ccc�*��KI��3opd*��$�����4,X��sU����,�k^���Lf�� 3�m۶ݮ��4(x�/B'��d�83g�ٷ��nG���0����g�ُ�@,�h������T��D���f��a�_�J%�J%T�U����k��a��,�R�i�8����\��k���ު:H+z{{U*���&�YD{0���u��q�ضm��:�!��x�uV�]��V�Z�	�Ґ�~jٲe�o��:q��� :�k!�T
�dRu��ٽ{wo�q���f��$fϞ�y��a���o����s��Eww���9���j�s ��f۶?�:H+�=�;��> �׋)I+��*��̠���pے%KzTiw����lڴ���ϟc����a����{��=��zAT�U������o�m۾>�;� 3��|���a�б3qED�Tg/5<<<�3�
��o�i�?�����|�YI�{�\~oWW���Y��Q&���#�����#�w ��e���Ҋ���'<�;��?@~Su�Aה�C1u��������Ui�6<`c�c�J%�ر����qT+�JR�ǈ������|�.�˹L&s�� �`��y_��M_�:�h���""�ވ�zM�\��{�f�膰�������~|�WD����=��T��dC�Fنa�2�͞�:H�����<�h �Af�#�0��3���@�ED�ض�5�9ځ����#fƞ={�k׮v;�R	Ţl���@���lW�V122"���f�[�9�"�����u/p$d6=��y��brD$G������8���~x�����̌;v`dd�]C�Z�\t�?�O
���Q[s.&e� ������7Wu�V���[��p6 yT=2K�)fު:��R6��;�!���v�i�Zų�>۱;����#>O�VR��P�_q��DtJ�X|8���:K���w]�r�4!��T���}_f�5EDR�3_��fߠ:H���� *A�����}�YT�� �V��vw�O�O
t�03*�
J�R��U*��~�;����i/7�l6��A��y�����Z��O�W�GL/�L�tM��/G�	1.��7e2��م������?��FFF�c���
Y�\�t�.&g�  "�/�J���>����'�L����g���Y��T�U�ݻWu�(��̷:���}��}ՁZU(�����E�X�<��|�i�R�����z!^`�a?t��uT�	�a�3�	�����عs���+T.������REDf�#�3�ill콭��x��Ν;1<<��וJE����sm۾}����T�	����.�u��}��U��s]7^V"-�B��| �,Z�h�� A0M�f 3�~-��x��8�@�R�\i���M
t��� �p`��[۠c���A���jJ"'�������番��P(��u�7��"��U����ޮ1���@⥖'��3�L�� �z��w�g&���o.���Q�TP,#S�Ʊ۷QR�+BD�v��s��Ig��r�6B����+|��9�󏪳�P(ܻp��# |�� "�>hLZ܅��(�0n���O���vs��|�N����J%2����O}R�+@D� .
c�N~�)�y[u��q��z{{Ӫ�%�˕]׽�R�LD���>Y���n wPBL��[�l�_"�����9s�D�G�����۷���+��rq��P���H�13wd��|���J���q^�:H��~��m�|�_��r���r��r�\�E���˶�KT�h�}��Wd�ۧ�{�#�Z�/I�C&��M
��Q7�S���m�Qo))�ˑi����`��Z�A�6<<��u���` �Bf�CEDR��O֡1�:��I�!ZaF�6�ZK��;���?�%V�H�.)��w�P7�}�;lFyS��ښ�?d��9D�=�q.[�bE(�a�<ϛ���� �@��B��R�kN֡ѐ��o��ٳ�I�U�Uii�8��t�������!�E/j��y�s�!��<��1՟���/Tx���#&	���[V��L�<d��mR�]�/_>�T*��OX�8N'�O�u�UB��8�-��K���X��-���D�7 ����cccعs�Q�4Mtw�u�@����]�= �7�E�bW7�8Eu�(�w��(Π��e��}��5��?j��<ϻFu�vx��'w�����[���CD�p��\�Ff��GD[�]��� ��?q�    IDAT�f�o���R�Y�|=� ���#���Z�b�޽���d7Qiq�E/��͖�Z�CDW;�s������.c��]�yޡ ���#u�0�@ל����.D㺘�N۶W�Y6l��R��{�9)�;T�Z���h��8�J�ޙ�)��T*Iq��w����e2�cTi'f�]׽�u���/��2�:�����d�M�GD?X�ti�� ��d2g<��sd���&Ez4D�@�� E���T*�n���c���9������1����|>�O�tz	��<�:STQ��a�Hvq�yK�����ŋϷm�v"���������C���R��z��pA�Qj�c��m�?�m�V&�\׽�� �7�@Eu�(�}��bj��K�.Ds�8�I��WOOω�e=JD��S�T�U���(�	"��J���2� �/ik����w�m��:HX������\�=ղ,�7fO��2��?iq�a% �W*����{���(����M;�s���?��T[��+mw����RQ)�e=@:_����#��m۾�q��:�b:����7f/3��� ��IS�0�A�\"��t!���M�i���O?�����9�R�� ����-!"$�I�1��rM���*E���⼳�;���L&s��,*�w]�l�����Q ��Τ�J�"�����bRDt/3����k7o�<�:�T��r�\ 8Tu��$	̚5�T
�TJu-�*�u�0T-*�̠w���1)�;-4��q�^�`�l�yT(
�x��5�u7�P �c�ͪs���,iq�3W<�:��Y�̯���'z����0�Y�d�+l��5� ĢJ5]]]H�����&�I)�먝�f�,z}Q)���}�C�o���J������H&��s�8�ATz�u����r�0^�����"ϟ??�����6w!�=����<�>�a�CD��8g����Zu��$	twwò���Y2��v�:|��H���^�����̠�Q�ƷVB�s�����x}���6����WR��-�S�q�jYֿ�v'@f���~�q>��'љ ވ�|.��������hx�+U�B�<�/x�w�DW����m�; �V�%,D�t:=ia���,���T�H���n{-3��Q�8Dԍ�[r*��I"Z��wx&",^���Yt�4���f�IIqkO2���0�l6���O'�3�y��<m����U��s� �V�C���eY�D�2�m���U �T�	K"�@*�j�������h{���S�]��M�#Q�w"z�aa��J�0���u(��CQ`|��7��⧶m��ma���9���3 ��"�y�`�u�e�C��9�� >�:�!���b���(�~r����f9�aH�R�Κ�#������k�����0��})���Ν�p�*��a(��ϟ����g�ٷ�������]�=��<����; v(�$YD4�:�!p�a�]�=?*����� x1*ΧZkިT*�D"`����t�gR���= ���vwwk�ce�XD�,�N�,a�۲�썙L� �at��U�u�y��{�w�>���T��E��� �נ��� \�H$���{����vՁe���m��ňIK{m���;����u�q��R�+ �<�S�m^��H$����O6~;��K�������JM���h��骳芙�CCC���{v:�^���) ��Ku���`f)�E�*��4�W��{ΦM����(�q�ǹ��r �U�	�eY�5kV��]]]R��Q�I�}9T+,R�+��� 8
������t��ϟ�ɢ�c�8�ϲ,��i$	̚5K���@D��F�q�\�dI��<:+
w��{�eY���o@t
ߨ�=���@���"z��gn޼yPu�fLY�(�s��!�N����m��R����>FGG-�eV�>)��(�O�OD�-���,p :蠺�:�}AHq^�i����z��k�f�,A��L�|<��~����4�����y�;-˚��̺�E�^�Dc����@��'�� ���|>�SuZ��d�f�Wa|r�`�qBc�f[f�'#Ez}2���]��W*�~>66�j��j��c6��a�4M�R)$��i_cf�
g����Y��������2�~�����¯U��E��J&�'1�i ���'~�uݳT��qg����>}�Z�~�P(�Au�fe2�3��" �:���a��{�6|/7D����wwp����]i���d2�P�����T*�ch�4�iל�f���rP�PD�a�a��8ε���P(<�:PT�`|S������K�ұ�a���=0��FD#*�M�\u!�� ~�����c�����&p� �j�Y�T�Oj�_��������`f����|�L�'-�1�!�y}���F�P��d�צ  g���q�")D���`�P(���9�����_�O�"�*Ẁl'"�����*�uO�</r������9�s��&p�)Ή�T*��Vstww��ޫ� ���V�>)�c�����5S��K֦?�  �ٶ�3�q�Bu���g7��\��3c��Xb)�#D�B� nc敮�\(Q�YDD�㼻T*����M�L�Dww�Vݤ��w��l3-�e�>����v^R��gF˻�&�Iy�;�u 68��u�q:jݑ
CCC���{����i.�"z �7��"��E�̠���1�w]�T��Uh&zzz^i���0�ɧ�eHa�a�|2A���T�"}&Kd�>�i��⼾�xF:>aV�� r�"��S� l޼y�u�K���� f�' w(<�̠G���M�Dt����N̘oPh&zzz�w������ب�Ю�=u�L:��`�&,˂i����jkқ-�e�>�$N�l�f\Y��+�J��,�Ÿ���?��m���l6{N>����@��u��� \�8N����Ll2w�%-��̠G�aO�͔�H	�`~>���3SDdٶ� >`��<ak��!���v�X�D"1e�e��J�2����L�tyC
t�fF�X�⼎ �ڧR{��QQv83��q������z�!Ձ:�뺣 ����C}�?�I Vb|#�f�z�����������y�ô¶��۶�5 �������Q+�j3�{���~��0$�Ɇ��3M�i"�L�Z��T*ͨ+���{Ծ���]�X�8���ɵk�|22��'��y��8_.��M5&644�8�����ۻ�R���d �0�� �ժ̠G���ò^P(���х�|�)�aZ�8N}��NV�E�d2�ok�v�����o��5�mh\*�P*��z��l��?�P)ڋ)ČqA�.@)�'W{����M�Y �O$��W֧�����f�u��� ����?���^CDR�GH�R�t��n 2�R�uωrq��ۻ�m���̱+�;�4�vwG�T��3��qmc�f��R#�������k�9���s��i��3ݱ1t��Z��l�>��� |��Tg�����e����� ���c
�¯��#"ö�"���%�h�6"�$�H|��'�ܩ:L+���[�l�{�t�9!�HtDa�b���u�����`Y�7G���IDH��u3X�ow]��N��]Q*Х8����R��7�b�rYu����?�#x�n���s��� ����E�B���Џ�8. [u����+Dt�ľ�ED��dN#�/X�:�
����~>�j����Q�Ez�7�k�aD���@�O
tMD�@��ڧ7k�,�~���C#>}�R�|B6��q��<`���#�g�K��w�9�7�m��a���+UgQ%�k͛��>��ı�Zِx��})��ӫ��i�CD���nk��4M̞=��<c�`��M�|�q�K-Z��C!f��:��(>��|�?�u�~��zq�����l6{#��⼓֚7�����5�a}�S�Ԍ���&�9�U"�\`���8�\m͹.m����i-75Q��������g�ϟ���Bt>)�E� \S�VW��{r�Px@u�V-]���q��}��3��:�*�D"�C�H�,+ԯw+m�/.ҥ��>)�c�ы���D6�O�5�ӱ,�f͒������/�N:�s��8]�	�))�E+�p!-s]�̧�z��Tj�m۶�8�T���pbz_]��H�ӱ�0M�������µs�}��8��LG�A��F.
��;籶�'�0���C��Q�VQ�V#�  J�yMmWM�4166&O0��@  ���8͛7�7n��b+!:��:���M .�}�ۅB�#�W\�x�|˲>FD� �"�Lm�v)��Y����n��Ώz�z�������Q��i�����1��S~��֜�Z0'��i�oL�|~F��Q*�f�	E��u�EX���E��z��;w����8��<��" 2�.�� _�<�Vf����:2��A�a�kY�?c|�Tl��T*���v������� "R�`���pN��V1�ښ�V.�D"�Y�f!�J55�LDH�R�3g��m�Q/�kjG�Ľ-��> �ڶ�G�q�"��Åh��b:cDt���Ǹ�{�����|���s�9�0�?�8b^��֚w�}P�X���{+U�mA���2�>�����T�N�aY�ŢVq-W'I$��e6�%��̶�Od��/��{-3�IĎ��O�Zx��J忟~��m��%��DD�����:�j�%r�v�.���b�ؖ�����%�k"�s�';���✈ڲ&[����J��Z���\.�����Z:�������h�Xq�9 ���!�@D��I�P���\.Z�hA"��g �� d�y+��r[�t"��ٳ��hxdZǝ�.��b������[)�j�mߵ<*��8瀬Mo@�����G���eY�����)@
����F _���S&H�L&k����� ȉ�Y� �s&}�=��A&p�O��������9o�k�F!�i"�J��Mh:�T*�yMmm�̦O)��r��)�q�eY�Ń��;T���
 V�!�X�r ׸���ݯB�t���j���0�B�weߗ̚'�H�������~��	�N^�%z�1sn��d��&�H$P.�C�`H�R���tT[�>::*�u�B ��T*�m��J����᭪s	�&r�Z�0�"�
�����4۶_ED� � �:3��dּ=��$�(�ɦR�����=�^0��K�Q��lX��6^\��"Bww���>����_�D�q��3���U�d'��Wp3�]�h��V�����8ΝD��wA���Y��Y�fIq�&�D"���J�j�c�\m�8��/���j`��a~��������C4�d6�a) g��.�q��y�uVJ��H�ޙ|"�3_�N�oإ:P�������o��1_�:�nj���i9�*�ɦR������!�n��]�q%zL�^��	�eY�}�ՓL&C�����l��Mo��$ 'e��{'v:���������! ���C�PpUj�����cccg1�9Dd�Σ�0��/d�^.����]|�o����3)�EKT�����)������X,���0�	Dt�m���\:66���[��Q�K���h� ���̷��۱����ޥ�J� �0Wqm���R)0s m㣣����~��A`f��P�W�8)�EKT<mmǇOM"��M��x�wѐ> ��J���8��Z������ͪC	ф��e�d����LDw�����L����s,3��O����e�&��t[���j����̌�����<���LƄ��EU�l�5��K�9�������x����H��+�����/��3��{���^�a�h��8��V�C�52���^�0������o�z{{��ry-}�a��茈�L&e����@f҃�K�Z�btt4
����{��A�'�B`�U_��gNf�g� p�a'9���o���]'��Bs�CT����7 d�<��1s,��N�_�� ����W�Gw2k��t:fF�Ri�}j��J�TjF���y�c�:R�k��#����JfЃdYV�gHv��Sy˲d6}f� pY*����8�ѷ���Fա��DR��R�[ 0�z˲~�y��Aա�DD�m��� �92�!rl�����0::�r���V�T`�&��$LӜvYj�ZE�RA�\�¬��ZCME
tM��'��/��䘦iJq0�0��ݍR�$��33����������:� ��g�|���`;����.`�%Lł ,RB�D�&4�6U��Ҩ�J���6Q�V�ꗪ$U�B)A�P�*bPp>ʚ$�ر��s��m`����3s��?f�@�ػ;���;�O�����#dݹ�}�=���� �
�� f�"Z���W�qyQUwx��7��=766֓����V�uW�T�,��]�I
N͓��%xs�:��Q���{H�*����&�������:C����D��z=��f���K�;u��伻��r��e�
�W �������W���Aס�籠w�������3k�O�$��u0��2-�,��r޷.�����ׇ�'Ov|%bEi]�ȂN��y��I,1�ˬ�qk�ڎ\\�(Swe2�Z�
sss<?sy6���~qa��l6�����n�Dg "դNZk xi~*�WU_�d2�\.��W���i��pj�|����NcA��ظq�G�qcI����N,�^X��∸^���O����Q1s��d��{���7T�� ~�:��(�����4���TT��b��x�W�V�㽲y�R����fff~MD�V�[�{�%��r��6D���]���P�
:�Y���g�~�4q
�BG�tx/�V��{4K�r���]�WD�����T*�|�G�Q*����~�9:m	���4�ry����7��:ORc:~6�É'8�x"��j�z���ħ��2��t,q���޶�D�-���G�����izW\���l6�������B���\6Kݠ���(�4^L# G�ީ>��Z;n����Ac��C�-�È0444h����b>�:O����,��)�0I�=�i���i��ǈ�� ���K��{w���.��ԭl�<�z��lv�q ����Z�U�';u���G��!i�L�����[U'Uu���ƍ���Q^���X,�g2���� >��ma��WN��Z���Y��w�����a�9:��x9�:�rXkq��Ɏ~Xt��r_�Fp���|FD>S*�j��?j�yx||�Y��(�D$P�8�WО|0!"GUur���Ƙp��յ={����$"�͛7�h���1�㪺�u�4�Լ�,��r��Ni|��)��w�ꃮstB'��h6����[ֹ�|�������"�_"� ߗ���}�1 ��9`JD�T�m��Z{�sDU'֯_��;>D$S,?$"w ���\gJ�k���a�o�Xk�Z�v�u�NbA���/�S�9:��\.��5�n6�h4�~B��y�Z-��u~�� �H/�C����?��E��:�%{RU��^n>`b~����y� ��1�C��pl��b�x�|)��י�haj�������oS	���!:�=FDĔJ�# 6���I"�L&��`����������Z�V��V�ձ������y�*���8M_y{<E�C�\��x+��wϿK�֢��B�V�W=ϛ�WEd�e;}D$S.�����ړ��Li%"����ԜN�$�MU���w\��4���}�Q�?�h���=:�-�� <b�yd|||��0D[�l�����оO�R6P�#N��tX�U�t�����i,�1���� ���I��y�Xk177ױ��$c��-�v�Ϫj�:�����U���""���Zיz���P(��3�^��tU��0]��4��9��.���q�#�V�Z�r�B���ƫ"���|>�̓θDD�7<<<�j�n�Q ; �&�-���bDQ����^�G:�E�Ctz̈��J� @�u�������Y)����뜦�GCU��oy����C��DDK#"^�T��	�� .u�'qjNKգ%�_� ������C�����9�����N�ck?�� �����yB�6����ͪz��|�9�3�2N�i�z��[k���j�w��X�c��������iz�D�G��mc̓�j�y��S��ÅF�����e���9Ʃ9�Wt�  	IDATuR������+�0���ނ=�|��1�+\爻��>~��0N����t��L&����Ó������0����,"����Eo�Ԝ�!�"�<��El��\����*�J_��s�#�X�	�N�	�sU�	��V������Qׁ�ҠX,^l����z����u&z'c��<�a�kR>IW�R�V��-,�1588���� �]g�#�s�E��'��`'����L��8�D{""��_� �[ko`!�?N�i��Z-�������a��:G7��ǘ��� ��s��9���bvvQģ�L��}�E�j��~ס�\�\.�Z��� l��m*:["�|>�l6�:
��f��z��:F���ӮCtz��J����s�%.
�?��8MO��D��Tu���Yc̮ R�v� ������Ƙ�D�:U�pU]"y��B���99����� �u��X�c�����]�9���Z�z��iz:�x����Zk����ܯ��u0������\� ר�"2�6u�](RT�?����m,�1����h/���5��|����i:��� �W�Qc̨��A��PD����> ��ȕ�z�+� `�KN��l,����Y�{z���h4�l6������0�N��joł� �R�oE�]�p�圖�Z���YX�k��𼈼 ��(�^���qll�OlhElٲem�Ѹ�Z{�|!��%���i�yr��Y��n݋/��v��[.������-�U]�Ƙ���ǟud%��'�ƍ�
�} ����4�s�N�i^@��w�ꋙLfo�Z��O�;�mۖ=v���(�.��D�RU��� ��|DDI�����o�αRX��\.RU��:�J��r���cP���t:�� ���>�`��v���`ett4�k�s6mڴ:��n�d2[U�"Q�_p!8'"��f�y����Q�AV
z����'Tu��+�场��hp�Ng�	���^ �E䀪V�������ӥ϶m۲�����:_ķ�`+zp%�K"�{�j�_]�XI,�	2<<<�j��p��,ݔ�fQ(\ǠE��:�M��j 8���cLEU+�Z���<8�8����LfHU�DdHD�Uu��%��p""�T��Z�����0�=a����T�1 ����\���C��p���U �Ƙ	UW�	 ���Z���!�dxx�`��`sE�Ed��=�P�����(�&������}z���W�?p���X��%N�ɑ9 � pTD�Yk�c����D�1�H��|����x�M�E��`�=�Z���`���;��&ٌv	���DD�	�A<�:�,�	422���������)�l�|�煒s��SL����¯U=n�9��3 fE�uUm��y#��"r"��4T������9��j��j��K	�iӦ�}}}�(�L&�Y7��� @E�UU�1kU5#"kUu�1f����NU׉�U]+"k �A�l�_��!""J�?��ˮC��P���p��,�%"K�n�eޘŝt�͇|oQavv����=�H��'DD��P�V�T��w�V,�	����������u�n�^yȱ�_�h4�䝈��he�,
������1;,�	W.��V��X�:���y��:�:�k��Q�T���D�v�7""""""J��l�f��6N�S��� |��3}-Q�6��[{�8���=%� xFD����BDDDDDt�-
7���z�T��=��mp�u"""""��x�P(|dll�5�A�K�S�.X�h4����k��0���G����)�J�p/���<DDDDD��Bk��Zm�� qƂ�r�ry��>�|�Y������'=��w�a��� qǂ�Ve��{ �	8M'""""��1��\���Wϳ�C���E�L�Uu��,DDDDD�Z���N���ǈ���;|ID��!""""�ty�Z{O�V��� IĂޣD���_G��_�:%��<i���0�:K�������~�����]�!""""��h��c �:ß��,�t��͛/�d2�p'��;��� �o6�NMMu&MX������ ��Rי�����ș9 ?�'U�� �\J+t:����(�nT�|�V }�cQw�`��|/���Ƙ]A̺�X�i�DD��lv��nU�� �Sյ"��* k�$""""�w�"2���8��o x�S���\DA�됽��������(�� DDDDDDDĂNDDDDDD�n|��1l�    IEND�B`�PK
     E"BY��C�I  I  /   images/d1a57a69-e5a0-4805-bdaf-8d975fdf5bdb.png�PNG

   IHDR   d   S   i��A   	pHYs  A  Ak!T�   tEXtSoftware www.inkscape.org��<  �IDATx���U�u��0<��y#�W|E�b�M�5V��6�������Sc�hMl�1I�G���51jbk5IU���F06A"UE�	�0�83�c�a�������s�=�{��~]߷�{�9���^{=����7`��ɦ��ǿT+8Qp���
{w򅱬��1���z�B��O?$8=����8��}����8<�}�1A��'�s�ۥ��r����C���O��ÇM�~��._�
��54���u~www�D�
t����wK 8�Np�`�`���"�>����0�mۛ�~�3v�	�_���r�u��R��3\�g&�@]]������_9��Ѓf!=j|I�E�u��	6K��%��� 8Dp��$�Y��
��#86���F�7hР�8y'΁�	絋��'�U������uMxQ�Cͤ���ꊈ4��^&���1v���C[��@�[p��s�fm �s��y���f������Q;!�rK`\ ���͡C���&�ǂ�'k�ȭi���y���}������g"
� b����|Bp�I�?f�l-8��C�S���b��竂���/c�}�������L�7��O�3����\�`~����N�jC��+��rD��$��f�w�Q�gq��H�~k7v�R���XL�so0V� �]�q��e�o��]"ߗ
�zX	��~0�&}� �q��'�5�S�52+AJ
�`���r`~'E	hY�d��'�%����K��p!�"���D�(��?%�Y�q>#���%�	����-HDc��S�uttDc�Qv���� ���@2�<��Cs0$
���*��4n�\�P����N�/����
n�5c�!S� !�pH}���6?%���|�Up�_X��0�>1�eT�;�H��~�=dȐh��L@�3�>�`���zfWða�v�{�ƍ�˭Ok�1��36g� T;�T�4�*�E�{�7+��J���I?�I�����	��P�R��*���ݣG��b^-?뛛�omii�$�8/�3�˂�͏$.��#��0�,�	�A�@����1��O��q 1mY�bOVE<��t�҆�����,!�b�U���ۯ*c��D�@�Ϗ)S��-[��k��Mu���Qx��#��F��!��\Ey�T%��BL��|�c`�|�-�lr��?'��`S�=q�����8S���/�D�rW
�,�wq�)�,P�X��3���X/�{3�A��1.4�X}B�,Vtm۶M�Yp��%t�.�r"R-(��_�Q~�+x\X^��<P��`��:{`mt�n�{���}F� -��3�}�TF�Ǔn̛7���է�P7jԨ�{������v�?q0|�y�*�!��|�`��=\�x�9�����C)f0��0I��X ?�/,X������4�]xekk��q^����	FO�
A�4�� �#� �ϭ��"�������3g�M�6�nz�f��Y�S����2nܸ!��A�뽂��b�e�p���-�8DT���4�'YEWE�E�#0��&oV����� ��9�FP��E�������f":��y��k@Q��B,B|��	��o֊�F9��]$U�*���lM����O�� ��ޒRn{���Ks>|�� %Q���o�䎎�C2����P����a�cC�K�^�UAQE,�G�����8P-��a��w��%�MNb<.3|�����4����|�'�\&�xF��V�>*�*�����ͥ�^�+
��x������5/��r���2p�0�	�qG�2{�V*��	&���/��M4�ս�bM	w|9�
��]�W��`�/�ҠAtQ�a�k{<�%�@TUCo��"��]�n�{�tV�E,(O�M����E�"!J�z�!,(�����2T���@���I�,�K
����MG�	��̾��ZU�����<y���s�obz�9��2]@��Sf��?��}�m߾�O�/���Z"��j���Cc�"�M��IVWn�0�@l0VnF�=��E���Y�_"��&a�4'\&��W���{�d o�s�|��Y��_��kiiQ�L?N��FV �&V3�׋IAH�J����������H/"�;Y�F13��<���2�mӦMC���"�f�PF����i��7���755�?Q��h'�z�޿���5�d��l�^}����I�&�k�@8B^�7�����X�a!s��':�h���뎝;w*q�ٻf�?� z�5� [��o7v�J�J���_�=����4��x�c�E�Z*�#�r����666�'��Ῐ�7����`�}2�|3�:�g��S� �6���g)a12+a�?2v-39O蜥^�~UpP����o׆�5 �I�f���} �����}���YwY@	��TWI}ɵ32V5��D�"��s�<?!$@�Θ`�L:�b�]�
!��P��X�gJH�~)&�_�㵒L�
�hӀ4 ,�>�4�n^������[u�@�_�%��,j��9�L�:��͛7�Q6����e��@���u���* i�������U��"!� �K�ڵ�T 
��M�6��-�2��.�p	6:��mG�9GO0vB�O*�� *C��]xX�p�8l���w�c�-�e���r�D��1�|f��*��f�	
W]ƿ���������zIN�GB�y��+���lv�X��&�yR������$3�*��s?ق�Gj���M��a,�l;׸��N��!T6�X+���ٕ�^�QD
��B.�����^��!$����;�i!��g���A������L�X�%+����E�(�=�P�̒�r�X�&�B�u�$�����Դ_���ls샆�p�Dd|b�D1��������OV���9��e���ث�Ʀp��
ΪnY`�M`b�56-	O���'��� A����J�"	�Q-B��!q)DY#ˍe���fo�����I��!��W8C��VWlJT�t��y������-��
��Xfv'$B�c������u�<"qr�=���[$�r�b2�rc��z���"�M���2y�VT�9��6lX���w�G��39 JL3f�Y�zu���YZ]Ie�z��s��5���2�{SA;����BC�i����on�ԩSu	7�ayCB���Ŧ �HWID�rVqf}�A�ys�M^����S���	10]��1�F���PF��ɚ	Y���M-G�V$�j��B�e�Tͼ�{V%�� B�g8d;��4����J"�qH8(Z�цH�5G�� W������<�C��è�<;$�#H��ˍ=���IKͱ�]�:��fAG�śBd������@D���At��'v�9��~���o���Y��_0v� �.�"��W�c��Gc��Z�`�w��!��,��+�� ';˅,B8�M1�).)����f_ɇ����g�!i���K��'	 �r�o�W���dEh�D� Ib�ƾ�c	�{*�8��������z\�����i7��3?cB�`��=����I@�P̕����$e�j�%��"Z�LG�,.S���+zJ�b�F�Sɣ�Fp@1�m.F��9J�am1��r��$9`a@�����⸩���z^��֮]۫`@�\���lm^@��s���M�ِE�[ӀX�g�+T� g��������c�ql�z�?��=�q�6`�)�ω�`��z�^�\�5�ё��Ϧ�%����EB62�l�o�z�8����n�EI������VnWR/���*�������ȭwĈ��N��UQ�ó����*�JJ��Y͌�L����E9bx��:2��,"�p�}��� ±y�L��o��� �X��E��PS9�TM��ⴂE	5ֻٰ�.�R�ܪ�r�#����p.����~z����:t�۷o%��XeX1i&9��F�'nӏ;��	�ۄ�?[I��ِlV:.�`Q���XXQ��q�)�DIN<�%-71<?dȐ�tvv;R����V��B!���0駶8�a��O����y\�	v
<��p%�C{4_�L�Ę;wn�\FQ#F�@��r[Ȇ|�7�#577�ٳgG�ۺu���A�e�g�X������\�2~�x�6�Z)�9�\c�_�(��L��L�� ����u�dV���;�q�t�4���K����E��q�~�)�&�Q���!�3�Mr�����w�!)w�1��fp��?	@R::r����>��� b���e����(Z�9g�+���,�P�F��q��utJ��8�m���vD�s!�ľ�^*�C�Y�'Z�.ܒ9�FS�@�Q	!7A�%Rcu�礡rއ� f>J�"��H��y XE*ǲ����y�G�<�_�7�\c<x��H��F�]?hР�ك��I�
�V��0�Yed�K�"��t�*�@t�e��G��'��=R��]r�V���+����l�C�� v��p�"�\l��U������Q�w7:nY���K(�3^X��&8�w��{R��)XR�]"�Q>Sk���o ��Y�����d=�"~�w�H���/w655�����Fyk�u���!�*�`�$(���<sD��$Q�,i"xL��+��2T���J	�?K/-�1��	��lժU*�XGG�ÊA�����-_4V���`�RVO�. �"�a�g<)��G���{!
l}���M/R�3�B@�UI��u���� K�;` ����9;�0�~L��K� �〔����}��n����5����!r�r������Y͌#
�������ߩ����J��(�/1BQU�KJI*rgk��yԨ�!]]}䎞���<Y��5v��PI��`;3��2���pPduA���2����E8�pv�=GV�e��ұ�*͓�r#J�����ڶ��/��/j��o +F'N�Â��ޒ���t�ia�� 9�!�� )����刣=@y�Z��=��v3�>�_*3�N�eVF�hA5|�BHƜ1N�a�EoE8��g�k83Ɣ�7���[]��_�>X���o{^`v�t���]I�>�Cp`��Nu�ݙ��4���	�Ń߰{�nD��~%pF�7�a̱�鐾Lk����+����~B�|Ѓ�P�QP����]�CX3��y�$��ve���YQ�:�Y&P�~A��1>���K�3@��Uro�|_V�����!�Dx��%����d����55�B�ڤwM%3��B��*��]��v:��ń���th��)� 'e9�&��{D�%��,�*�G� 7�����zC�I_�]*�Dw�9|��Ƭ�x���Ms��Ɖ��W/����4
1Ȓ��݄(�<ĩB��;d9����b���d�x�4�����m۶�<s�̗:::NOz=�B���LT"�h2�<�?��pa���p���`89�>wn�K�"�-q�!�sF������b�8��C�Nj;v�g�3N�ed���a�{GD�bq�a�{��:��}R���#}J<�(y:����Mc�B���:b��$	;�#C�Pw����j��A�gI�G��&�,�mH�ަ�B
E7���I�
�����I(%X��g$��i��i@p�/�!�p�W�=���1���u�&�����m�__`9A��)�:�����jڪ���C�ꦯ~J{�E&O]de����=�S���eM�3{�}M����Ʀ���nu�(#�&����� ! i?��ܻ�y$���#t���ߥ��qqi'(�e���{�[�|��;�3G_&pyJ�ǩk�����U�Y����u ����+4
]�Hð��`q
{F9�]��}�ɞ�"�(L\�
����?g%�9�¯�K�T�Ǝ��w�� l}�t�H)���l��kG�v,i"��G؃��w8��>���$LF�~��#Jc7���r�.A�ϥ/݌���PPV���KAB=�_�%�+T����Z�n�,�rѓ���1�6�Db��2��GXRE$�e��Z��:�5��:Y�_�K�����}�Gd�b�"�������,�P٪��M Xn�C�9~A�<J���z^:���ۢ	��~�_ �p�,4eN��3�}��}ǔer��C�<A��GD��x!z�Nk��HE`��3o�8�4�M ���A��_��k�=d�8"%sB�[pT��?O�@g ��o�3���.8�b�W    IEND�B`�PK 
     B"BY.u��� �                  cirkitFile.jsonPK 
     B"BY                        � jsons/PK 
     B"BY�h���`  �`               � jsons/user_defined.jsonPK 
     B"BY                        �u images/PK 
     B"BYP��/ǽ  ǽ  /             v images/0b351edc-7875-4477-b820-546ce15be531.pngPK 
     B"BY$7h�!  �!  /             #4 images/e0155ecf-753f-4e63-a512-9d8bb2c3e0aa.pngPK 
     B"BY,��2�� �� /             aV images/e28c3bbb-5472-4456-9ec9-e60c5bfdece2.pngPK 
     B"BY�ʩ��*  �*  /             � images/9a88a734-d46c-4092-86bc-e9f7b966a1ec.pngPK 
     B"BY�U���? �? /             �7 images/05596fff-4f8f-4556-8b1d-73ff55b6eaa8.pngPK 
     B"BY<��G�4  �4  /             �w images/e4b09d94-725a-4fc8-8861-adc4f6b1a3b4.pngPK 
     C"BY���+� +� /             �� images/c49304c6-1828-42f7-9c78-6513b79a7c1a.pngPK 
     C"BY���    /             %? images/86ae6a4b-562d-4e93-9595-3c4b0d09f42e.pngPK 
     C"BY"-�' ' /             �Z images/43e4be74-284e-4582-91bd-e4a77387caa5.pngPK 
     C"BYW�����  ��  /             �a images/a3b4885c-2487-4906-a080-ee9b44acb175.pngPK 
     D"BYq���W W /              images/7c9bed20-c7d7-43dc-b689-820375f46db8.pngPK 
     D"BY$�3  3  /             de" images/7ade412b-fa94-47ea-987a-d6c9baa14438.pngPK 
     C"BYg�Ѧ�h  �h  /             �|" images/4d53c106-8e41-4afb-b8f1-56dd58def1e6.pngPK 
     C"BYw��V�e  �e  /             ��" images/d004afae-d6a3-4a65-a5d4-4f8d37106046.pngPK 
     D"BYW���  /             �K# images/19f08d4b-a68c-4e36-96dd-32682874608f.pngPK 
     D"BY��Ed  d  /             W$ images/5779bcfa-264f-4061-b24b-5c8b50561781.pngPK 
     E"BY	��} } /             �i$ images/bbfae99c-8036-4c5e-89fd-a87441410720.pngPK 
     E"BYd��   �   /             �% images/a262aa33-74c4-460b-b0ad-c746896f6744.pngPK 
     E"BY?S�2� 2� /             �& images/da48ab5c-24bb-4ba8-ab59-39208c7b2ba2.pngPK 
     E"BY$�8��  �  /             k�) images/b96c8ad8-7845-422d-b49f-326b2968fdb8.pngPK 
     D"BYWC�� � /             ��) images/f1393e3f-31c1-44d6-9d33-bf195c230c11.pngPK 
     D"BY��_3
  3
  /             R�* images/1ff35573-e276-4514-8c59-6294c96ecf57.pngPK 
     E"BY
�8b  8b  /             �+ images/a7e3301e-fb46-458d-916f-a05c0bde95f4.pngPK 
     E"BY'�Y��  �  /             Wi+ images/4bf63cb1-3675-4452-8ab6-1403298522d5.pngPK 
     E"BY�}���) �) /             jm+ images/146a6d58-0553-42c9-b8c7-03425202d69a.pngPK 
     E"BY��C�I  I  /             ��, images/d1a57a69-e5a0-4805-bdaf-8d975fdf5bdb.pngPK      ]
  :�,   